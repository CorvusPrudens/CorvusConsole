// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 27 2020 03:05:37

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    BUFFER_DATA_OUT,
    BUFFER_DATA_IN,
    BUFFER_ADDRESS,
    A13,
    D6_in,
    A9,
    D3,
    CLK,
    A6,
    RX,
    D8_in,
    D7,
    D12,
    CE,
    D9_in,
    D5_in,
    D0_in,
    B_OE,
    A10,
    D10_in,
    A8,
    D11_in,
    D0,
    A1,
    GPIO11,
    D4_in,
    GPIO9,
    A14,
    LB,
    D4,
    D13_in,
    D11,
    B_CE,
    A5,
    D14_in,
    B_WR,
    A2,
    A11,
    D6,
    D13,
    B_LB,
    D1,
    A0,
    OE,
    D8,
    D15,
    D15_in,
    A15,
    UB,
    D5,
    D10,
    A4,
    GPIO3,
    D1_in,
    TX,
    D7_in,
    A3,
    D9,
    D14,
    WR,
    D3_in,
    A12,
    D2_in,
    D12_in,
    D2,
    B_UB,
    A7);

    output [15:0] BUFFER_DATA_OUT;
    input [15:0] BUFFER_DATA_IN;
    output [15:0] BUFFER_ADDRESS;
    output A13;
    input D6_in;
    output A9;
    output D3;
    input CLK;
    output A6;
    input RX;
    input D8_in;
    output D7;
    output D12;
    output CE;
    input D9_in;
    input D5_in;
    input D0_in;
    output B_OE;
    output A10;
    input D10_in;
    output A8;
    input D11_in;
    output D0;
    output A1;
    output GPIO11;
    input D4_in;
    output GPIO9;
    output A14;
    output LB;
    output D4;
    input D13_in;
    output D11;
    output B_CE;
    output A5;
    input D14_in;
    output B_WR;
    output A2;
    output A11;
    output D6;
    output D13;
    output B_LB;
    output D1;
    output A0;
    output OE;
    output D8;
    output D15;
    input D15_in;
    output A15;
    output UB;
    output D5;
    output D10;
    output A4;
    output GPIO3;
    input D1_in;
    output TX;
    input D7_in;
    output A3;
    output D9;
    output D14;
    output WR;
    input D3_in;
    output A12;
    input D2_in;
    input D12_in;
    output D2;
    output B_UB;
    output A7;

    wire N__80918;
    wire N__80917;
    wire N__80916;
    wire N__80907;
    wire N__80906;
    wire N__80905;
    wire N__80898;
    wire N__80897;
    wire N__80896;
    wire N__80889;
    wire N__80888;
    wire N__80887;
    wire N__80880;
    wire N__80879;
    wire N__80878;
    wire N__80871;
    wire N__80870;
    wire N__80869;
    wire N__80862;
    wire N__80861;
    wire N__80860;
    wire N__80853;
    wire N__80852;
    wire N__80851;
    wire N__80844;
    wire N__80843;
    wire N__80842;
    wire N__80835;
    wire N__80834;
    wire N__80833;
    wire N__80826;
    wire N__80825;
    wire N__80824;
    wire N__80817;
    wire N__80816;
    wire N__80815;
    wire N__80808;
    wire N__80807;
    wire N__80806;
    wire N__80799;
    wire N__80798;
    wire N__80797;
    wire N__80790;
    wire N__80789;
    wire N__80788;
    wire N__80781;
    wire N__80780;
    wire N__80779;
    wire N__80772;
    wire N__80771;
    wire N__80770;
    wire N__80763;
    wire N__80762;
    wire N__80761;
    wire N__80754;
    wire N__80753;
    wire N__80752;
    wire N__80745;
    wire N__80744;
    wire N__80743;
    wire N__80736;
    wire N__80735;
    wire N__80734;
    wire N__80727;
    wire N__80726;
    wire N__80725;
    wire N__80718;
    wire N__80717;
    wire N__80716;
    wire N__80709;
    wire N__80708;
    wire N__80707;
    wire N__80700;
    wire N__80699;
    wire N__80698;
    wire N__80691;
    wire N__80690;
    wire N__80689;
    wire N__80682;
    wire N__80681;
    wire N__80680;
    wire N__80673;
    wire N__80672;
    wire N__80671;
    wire N__80664;
    wire N__80663;
    wire N__80662;
    wire N__80655;
    wire N__80654;
    wire N__80653;
    wire N__80646;
    wire N__80645;
    wire N__80644;
    wire N__80637;
    wire N__80636;
    wire N__80635;
    wire N__80628;
    wire N__80627;
    wire N__80626;
    wire N__80619;
    wire N__80618;
    wire N__80617;
    wire N__80610;
    wire N__80609;
    wire N__80608;
    wire N__80601;
    wire N__80600;
    wire N__80599;
    wire N__80592;
    wire N__80591;
    wire N__80590;
    wire N__80583;
    wire N__80582;
    wire N__80581;
    wire N__80574;
    wire N__80573;
    wire N__80572;
    wire N__80565;
    wire N__80564;
    wire N__80563;
    wire N__80556;
    wire N__80555;
    wire N__80554;
    wire N__80547;
    wire N__80546;
    wire N__80545;
    wire N__80538;
    wire N__80537;
    wire N__80536;
    wire N__80529;
    wire N__80528;
    wire N__80527;
    wire N__80520;
    wire N__80519;
    wire N__80518;
    wire N__80511;
    wire N__80510;
    wire N__80509;
    wire N__80502;
    wire N__80501;
    wire N__80500;
    wire N__80493;
    wire N__80492;
    wire N__80491;
    wire N__80484;
    wire N__80483;
    wire N__80482;
    wire N__80475;
    wire N__80474;
    wire N__80473;
    wire N__80466;
    wire N__80465;
    wire N__80464;
    wire N__80457;
    wire N__80456;
    wire N__80455;
    wire N__80448;
    wire N__80447;
    wire N__80446;
    wire N__80439;
    wire N__80438;
    wire N__80437;
    wire N__80430;
    wire N__80429;
    wire N__80428;
    wire N__80421;
    wire N__80420;
    wire N__80419;
    wire N__80412;
    wire N__80411;
    wire N__80410;
    wire N__80403;
    wire N__80402;
    wire N__80401;
    wire N__80394;
    wire N__80393;
    wire N__80392;
    wire N__80385;
    wire N__80384;
    wire N__80383;
    wire N__80376;
    wire N__80375;
    wire N__80374;
    wire N__80367;
    wire N__80366;
    wire N__80365;
    wire N__80358;
    wire N__80357;
    wire N__80356;
    wire N__80349;
    wire N__80348;
    wire N__80347;
    wire N__80340;
    wire N__80339;
    wire N__80338;
    wire N__80331;
    wire N__80330;
    wire N__80329;
    wire N__80322;
    wire N__80321;
    wire N__80320;
    wire N__80313;
    wire N__80312;
    wire N__80311;
    wire N__80304;
    wire N__80303;
    wire N__80302;
    wire N__80295;
    wire N__80294;
    wire N__80293;
    wire N__80286;
    wire N__80285;
    wire N__80284;
    wire N__80277;
    wire N__80276;
    wire N__80275;
    wire N__80268;
    wire N__80267;
    wire N__80266;
    wire N__80259;
    wire N__80258;
    wire N__80257;
    wire N__80250;
    wire N__80249;
    wire N__80248;
    wire N__80241;
    wire N__80240;
    wire N__80239;
    wire N__80232;
    wire N__80231;
    wire N__80230;
    wire N__80223;
    wire N__80222;
    wire N__80221;
    wire N__80214;
    wire N__80213;
    wire N__80212;
    wire N__80205;
    wire N__80204;
    wire N__80203;
    wire N__80196;
    wire N__80195;
    wire N__80194;
    wire N__80187;
    wire N__80186;
    wire N__80185;
    wire N__80178;
    wire N__80177;
    wire N__80176;
    wire N__80169;
    wire N__80168;
    wire N__80167;
    wire N__80160;
    wire N__80159;
    wire N__80158;
    wire N__80151;
    wire N__80150;
    wire N__80149;
    wire N__80142;
    wire N__80141;
    wire N__80140;
    wire N__80133;
    wire N__80132;
    wire N__80131;
    wire N__80124;
    wire N__80123;
    wire N__80122;
    wire N__80115;
    wire N__80114;
    wire N__80113;
    wire N__80106;
    wire N__80105;
    wire N__80104;
    wire N__80097;
    wire N__80096;
    wire N__80095;
    wire N__80088;
    wire N__80087;
    wire N__80086;
    wire N__80079;
    wire N__80078;
    wire N__80077;
    wire N__80070;
    wire N__80069;
    wire N__80068;
    wire N__80061;
    wire N__80060;
    wire N__80059;
    wire N__80052;
    wire N__80051;
    wire N__80050;
    wire N__80043;
    wire N__80042;
    wire N__80041;
    wire N__80034;
    wire N__80033;
    wire N__80032;
    wire N__80025;
    wire N__80024;
    wire N__80023;
    wire N__80016;
    wire N__80015;
    wire N__80014;
    wire N__80007;
    wire N__80006;
    wire N__80005;
    wire N__79998;
    wire N__79997;
    wire N__79996;
    wire N__79989;
    wire N__79988;
    wire N__79987;
    wire N__79980;
    wire N__79979;
    wire N__79978;
    wire N__79971;
    wire N__79970;
    wire N__79969;
    wire N__79962;
    wire N__79961;
    wire N__79960;
    wire N__79953;
    wire N__79952;
    wire N__79951;
    wire N__79944;
    wire N__79943;
    wire N__79942;
    wire N__79935;
    wire N__79934;
    wire N__79933;
    wire N__79926;
    wire N__79925;
    wire N__79924;
    wire N__79907;
    wire N__79904;
    wire N__79901;
    wire N__79898;
    wire N__79897;
    wire N__79896;
    wire N__79895;
    wire N__79892;
    wire N__79891;
    wire N__79890;
    wire N__79887;
    wire N__79884;
    wire N__79883;
    wire N__79882;
    wire N__79881;
    wire N__79880;
    wire N__79879;
    wire N__79878;
    wire N__79875;
    wire N__79874;
    wire N__79873;
    wire N__79872;
    wire N__79871;
    wire N__79870;
    wire N__79867;
    wire N__79866;
    wire N__79863;
    wire N__79862;
    wire N__79861;
    wire N__79860;
    wire N__79859;
    wire N__79858;
    wire N__79857;
    wire N__79854;
    wire N__79851;
    wire N__79850;
    wire N__79847;
    wire N__79846;
    wire N__79845;
    wire N__79844;
    wire N__79843;
    wire N__79842;
    wire N__79841;
    wire N__79840;
    wire N__79839;
    wire N__79838;
    wire N__79835;
    wire N__79834;
    wire N__79833;
    wire N__79832;
    wire N__79831;
    wire N__79830;
    wire N__79819;
    wire N__79818;
    wire N__79815;
    wire N__79812;
    wire N__79809;
    wire N__79808;
    wire N__79801;
    wire N__79798;
    wire N__79795;
    wire N__79792;
    wire N__79789;
    wire N__79788;
    wire N__79787;
    wire N__79784;
    wire N__79783;
    wire N__79778;
    wire N__79775;
    wire N__79772;
    wire N__79769;
    wire N__79766;
    wire N__79763;
    wire N__79762;
    wire N__79761;
    wire N__79758;
    wire N__79755;
    wire N__79752;
    wire N__79751;
    wire N__79748;
    wire N__79747;
    wire N__79744;
    wire N__79741;
    wire N__79738;
    wire N__79735;
    wire N__79732;
    wire N__79729;
    wire N__79726;
    wire N__79723;
    wire N__79716;
    wire N__79715;
    wire N__79714;
    wire N__79711;
    wire N__79708;
    wire N__79705;
    wire N__79698;
    wire N__79695;
    wire N__79692;
    wire N__79683;
    wire N__79678;
    wire N__79675;
    wire N__79672;
    wire N__79667;
    wire N__79662;
    wire N__79657;
    wire N__79652;
    wire N__79649;
    wire N__79644;
    wire N__79641;
    wire N__79638;
    wire N__79635;
    wire N__79628;
    wire N__79621;
    wire N__79614;
    wire N__79613;
    wire N__79610;
    wire N__79605;
    wire N__79598;
    wire N__79591;
    wire N__79584;
    wire N__79581;
    wire N__79578;
    wire N__79573;
    wire N__79556;
    wire N__79553;
    wire N__79532;
    wire N__79531;
    wire N__79530;
    wire N__79529;
    wire N__79528;
    wire N__79527;
    wire N__79524;
    wire N__79523;
    wire N__79522;
    wire N__79519;
    wire N__79516;
    wire N__79515;
    wire N__79514;
    wire N__79511;
    wire N__79508;
    wire N__79507;
    wire N__79504;
    wire N__79503;
    wire N__79502;
    wire N__79501;
    wire N__79500;
    wire N__79499;
    wire N__79498;
    wire N__79497;
    wire N__79496;
    wire N__79495;
    wire N__79490;
    wire N__79489;
    wire N__79488;
    wire N__79487;
    wire N__79486;
    wire N__79483;
    wire N__79474;
    wire N__79469;
    wire N__79464;
    wire N__79461;
    wire N__79458;
    wire N__79457;
    wire N__79456;
    wire N__79455;
    wire N__79454;
    wire N__79453;
    wire N__79452;
    wire N__79447;
    wire N__79440;
    wire N__79437;
    wire N__79434;
    wire N__79433;
    wire N__79432;
    wire N__79431;
    wire N__79428;
    wire N__79425;
    wire N__79422;
    wire N__79421;
    wire N__79420;
    wire N__79419;
    wire N__79418;
    wire N__79417;
    wire N__79416;
    wire N__79415;
    wire N__79414;
    wire N__79413;
    wire N__79412;
    wire N__79411;
    wire N__79408;
    wire N__79405;
    wire N__79398;
    wire N__79395;
    wire N__79392;
    wire N__79391;
    wire N__79388;
    wire N__79381;
    wire N__79378;
    wire N__79373;
    wire N__79370;
    wire N__79367;
    wire N__79358;
    wire N__79355;
    wire N__79352;
    wire N__79343;
    wire N__79342;
    wire N__79341;
    wire N__79336;
    wire N__79333;
    wire N__79328;
    wire N__79327;
    wire N__79324;
    wire N__79323;
    wire N__79322;
    wire N__79321;
    wire N__79320;
    wire N__79319;
    wire N__79318;
    wire N__79315;
    wire N__79314;
    wire N__79309;
    wire N__79306;
    wire N__79301;
    wire N__79300;
    wire N__79299;
    wire N__79298;
    wire N__79297;
    wire N__79294;
    wire N__79293;
    wire N__79290;
    wire N__79287;
    wire N__79286;
    wire N__79277;
    wire N__79274;
    wire N__79269;
    wire N__79262;
    wire N__79259;
    wire N__79256;
    wire N__79253;
    wire N__79250;
    wire N__79249;
    wire N__79248;
    wire N__79245;
    wire N__79238;
    wire N__79233;
    wire N__79228;
    wire N__79223;
    wire N__79220;
    wire N__79217;
    wire N__79214;
    wire N__79211;
    wire N__79210;
    wire N__79209;
    wire N__79208;
    wire N__79207;
    wire N__79204;
    wire N__79201;
    wire N__79196;
    wire N__79193;
    wire N__79190;
    wire N__79185;
    wire N__79182;
    wire N__79179;
    wire N__79176;
    wire N__79171;
    wire N__79162;
    wire N__79157;
    wire N__79150;
    wire N__79143;
    wire N__79142;
    wire N__79139;
    wire N__79134;
    wire N__79131;
    wire N__79126;
    wire N__79123;
    wire N__79116;
    wire N__79111;
    wire N__79104;
    wire N__79091;
    wire N__79088;
    wire N__79067;
    wire N__79064;
    wire N__79061;
    wire N__79058;
    wire N__79055;
    wire N__79052;
    wire N__79049;
    wire N__79048;
    wire N__79045;
    wire N__79044;
    wire N__79043;
    wire N__79040;
    wire N__79037;
    wire N__79034;
    wire N__79033;
    wire N__79030;
    wire N__79027;
    wire N__79024;
    wire N__79021;
    wire N__79016;
    wire N__79011;
    wire N__79006;
    wire N__79001;
    wire N__78998;
    wire N__78997;
    wire N__78996;
    wire N__78995;
    wire N__78994;
    wire N__78993;
    wire N__78990;
    wire N__78989;
    wire N__78988;
    wire N__78985;
    wire N__78984;
    wire N__78981;
    wire N__78980;
    wire N__78977;
    wire N__78972;
    wire N__78969;
    wire N__78966;
    wire N__78963;
    wire N__78960;
    wire N__78957;
    wire N__78956;
    wire N__78955;
    wire N__78952;
    wire N__78949;
    wire N__78944;
    wire N__78943;
    wire N__78940;
    wire N__78937;
    wire N__78934;
    wire N__78929;
    wire N__78924;
    wire N__78921;
    wire N__78918;
    wire N__78915;
    wire N__78912;
    wire N__78905;
    wire N__78900;
    wire N__78887;
    wire N__78884;
    wire N__78881;
    wire N__78878;
    wire N__78875;
    wire N__78872;
    wire N__78869;
    wire N__78866;
    wire N__78863;
    wire N__78862;
    wire N__78861;
    wire N__78860;
    wire N__78859;
    wire N__78858;
    wire N__78857;
    wire N__78856;
    wire N__78855;
    wire N__78854;
    wire N__78853;
    wire N__78852;
    wire N__78851;
    wire N__78850;
    wire N__78849;
    wire N__78846;
    wire N__78845;
    wire N__78844;
    wire N__78843;
    wire N__78842;
    wire N__78841;
    wire N__78840;
    wire N__78839;
    wire N__78838;
    wire N__78837;
    wire N__78836;
    wire N__78835;
    wire N__78834;
    wire N__78833;
    wire N__78832;
    wire N__78831;
    wire N__78830;
    wire N__78829;
    wire N__78828;
    wire N__78827;
    wire N__78824;
    wire N__78823;
    wire N__78820;
    wire N__78819;
    wire N__78818;
    wire N__78815;
    wire N__78814;
    wire N__78813;
    wire N__78812;
    wire N__78811;
    wire N__78810;
    wire N__78809;
    wire N__78808;
    wire N__78807;
    wire N__78806;
    wire N__78799;
    wire N__78798;
    wire N__78797;
    wire N__78796;
    wire N__78795;
    wire N__78794;
    wire N__78793;
    wire N__78792;
    wire N__78791;
    wire N__78790;
    wire N__78789;
    wire N__78788;
    wire N__78787;
    wire N__78780;
    wire N__78779;
    wire N__78778;
    wire N__78777;
    wire N__78776;
    wire N__78775;
    wire N__78774;
    wire N__78773;
    wire N__78770;
    wire N__78769;
    wire N__78768;
    wire N__78767;
    wire N__78766;
    wire N__78761;
    wire N__78754;
    wire N__78753;
    wire N__78750;
    wire N__78747;
    wire N__78746;
    wire N__78745;
    wire N__78744;
    wire N__78741;
    wire N__78738;
    wire N__78737;
    wire N__78736;
    wire N__78735;
    wire N__78734;
    wire N__78733;
    wire N__78732;
    wire N__78731;
    wire N__78730;
    wire N__78729;
    wire N__78728;
    wire N__78727;
    wire N__78724;
    wire N__78721;
    wire N__78720;
    wire N__78719;
    wire N__78718;
    wire N__78715;
    wire N__78714;
    wire N__78713;
    wire N__78712;
    wire N__78705;
    wire N__78704;
    wire N__78701;
    wire N__78700;
    wire N__78697;
    wire N__78696;
    wire N__78695;
    wire N__78694;
    wire N__78693;
    wire N__78692;
    wire N__78689;
    wire N__78688;
    wire N__78687;
    wire N__78686;
    wire N__78685;
    wire N__78680;
    wire N__78679;
    wire N__78678;
    wire N__78677;
    wire N__78672;
    wire N__78663;
    wire N__78652;
    wire N__78641;
    wire N__78640;
    wire N__78639;
    wire N__78638;
    wire N__78637;
    wire N__78636;
    wire N__78635;
    wire N__78634;
    wire N__78631;
    wire N__78626;
    wire N__78625;
    wire N__78622;
    wire N__78613;
    wire N__78606;
    wire N__78597;
    wire N__78594;
    wire N__78591;
    wire N__78588;
    wire N__78583;
    wire N__78574;
    wire N__78573;
    wire N__78570;
    wire N__78569;
    wire N__78560;
    wire N__78555;
    wire N__78552;
    wire N__78547;
    wire N__78544;
    wire N__78543;
    wire N__78542;
    wire N__78537;
    wire N__78532;
    wire N__78523;
    wire N__78516;
    wire N__78507;
    wire N__78506;
    wire N__78505;
    wire N__78502;
    wire N__78499;
    wire N__78496;
    wire N__78489;
    wire N__78484;
    wire N__78483;
    wire N__78482;
    wire N__78479;
    wire N__78476;
    wire N__78475;
    wire N__78474;
    wire N__78473;
    wire N__78472;
    wire N__78469;
    wire N__78468;
    wire N__78457;
    wire N__78454;
    wire N__78447;
    wire N__78442;
    wire N__78437;
    wire N__78434;
    wire N__78431;
    wire N__78426;
    wire N__78417;
    wire N__78410;
    wire N__78407;
    wire N__78406;
    wire N__78405;
    wire N__78404;
    wire N__78399;
    wire N__78396;
    wire N__78391;
    wire N__78388;
    wire N__78379;
    wire N__78372;
    wire N__78369;
    wire N__78366;
    wire N__78363;
    wire N__78362;
    wire N__78361;
    wire N__78360;
    wire N__78359;
    wire N__78358;
    wire N__78355;
    wire N__78352;
    wire N__78345;
    wire N__78340;
    wire N__78339;
    wire N__78338;
    wire N__78337;
    wire N__78336;
    wire N__78335;
    wire N__78334;
    wire N__78333;
    wire N__78332;
    wire N__78331;
    wire N__78330;
    wire N__78329;
    wire N__78328;
    wire N__78327;
    wire N__78326;
    wire N__78325;
    wire N__78324;
    wire N__78323;
    wire N__78322;
    wire N__78321;
    wire N__78320;
    wire N__78319;
    wire N__78316;
    wire N__78315;
    wire N__78312;
    wire N__78305;
    wire N__78300;
    wire N__78295;
    wire N__78290;
    wire N__78287;
    wire N__78282;
    wire N__78277;
    wire N__78272;
    wire N__78265;
    wire N__78258;
    wire N__78237;
    wire N__78234;
    wire N__78227;
    wire N__78214;
    wire N__78209;
    wire N__78206;
    wire N__78203;
    wire N__78194;
    wire N__78185;
    wire N__78178;
    wire N__78169;
    wire N__78160;
    wire N__78151;
    wire N__78142;
    wire N__78133;
    wire N__78124;
    wire N__78107;
    wire N__78100;
    wire N__78071;
    wire N__78070;
    wire N__78069;
    wire N__78068;
    wire N__78067;
    wire N__78066;
    wire N__78065;
    wire N__78064;
    wire N__78063;
    wire N__78062;
    wire N__78061;
    wire N__78060;
    wire N__78059;
    wire N__78056;
    wire N__78055;
    wire N__78054;
    wire N__78051;
    wire N__78050;
    wire N__78049;
    wire N__78044;
    wire N__78043;
    wire N__78042;
    wire N__78041;
    wire N__78040;
    wire N__78039;
    wire N__78038;
    wire N__78037;
    wire N__78036;
    wire N__78035;
    wire N__78032;
    wire N__78029;
    wire N__78028;
    wire N__78027;
    wire N__78026;
    wire N__78025;
    wire N__78024;
    wire N__78023;
    wire N__78022;
    wire N__78021;
    wire N__78020;
    wire N__78017;
    wire N__78012;
    wire N__78011;
    wire N__78006;
    wire N__78003;
    wire N__77996;
    wire N__77995;
    wire N__77994;
    wire N__77993;
    wire N__77990;
    wire N__77989;
    wire N__77988;
    wire N__77983;
    wire N__77982;
    wire N__77981;
    wire N__77978;
    wire N__77977;
    wire N__77976;
    wire N__77975;
    wire N__77974;
    wire N__77973;
    wire N__77970;
    wire N__77967;
    wire N__77966;
    wire N__77965;
    wire N__77962;
    wire N__77961;
    wire N__77958;
    wire N__77957;
    wire N__77956;
    wire N__77955;
    wire N__77954;
    wire N__77953;
    wire N__77950;
    wire N__77947;
    wire N__77944;
    wire N__77941;
    wire N__77940;
    wire N__77937;
    wire N__77934;
    wire N__77933;
    wire N__77932;
    wire N__77929;
    wire N__77926;
    wire N__77921;
    wire N__77912;
    wire N__77911;
    wire N__77910;
    wire N__77909;
    wire N__77908;
    wire N__77907;
    wire N__77906;
    wire N__77903;
    wire N__77900;
    wire N__77899;
    wire N__77898;
    wire N__77897;
    wire N__77896;
    wire N__77895;
    wire N__77894;
    wire N__77893;
    wire N__77892;
    wire N__77889;
    wire N__77888;
    wire N__77887;
    wire N__77886;
    wire N__77885;
    wire N__77884;
    wire N__77883;
    wire N__77882;
    wire N__77881;
    wire N__77880;
    wire N__77879;
    wire N__77878;
    wire N__77877;
    wire N__77876;
    wire N__77875;
    wire N__77874;
    wire N__77873;
    wire N__77870;
    wire N__77867;
    wire N__77866;
    wire N__77865;
    wire N__77864;
    wire N__77863;
    wire N__77862;
    wire N__77859;
    wire N__77856;
    wire N__77853;
    wire N__77850;
    wire N__77847;
    wire N__77844;
    wire N__77843;
    wire N__77842;
    wire N__77841;
    wire N__77840;
    wire N__77839;
    wire N__77838;
    wire N__77829;
    wire N__77826;
    wire N__77817;
    wire N__77816;
    wire N__77813;
    wire N__77812;
    wire N__77809;
    wire N__77808;
    wire N__77807;
    wire N__77806;
    wire N__77805;
    wire N__77804;
    wire N__77803;
    wire N__77800;
    wire N__77797;
    wire N__77796;
    wire N__77795;
    wire N__77794;
    wire N__77793;
    wire N__77790;
    wire N__77785;
    wire N__77778;
    wire N__77775;
    wire N__77766;
    wire N__77755;
    wire N__77752;
    wire N__77745;
    wire N__77744;
    wire N__77743;
    wire N__77740;
    wire N__77733;
    wire N__77730;
    wire N__77723;
    wire N__77720;
    wire N__77715;
    wire N__77708;
    wire N__77701;
    wire N__77700;
    wire N__77697;
    wire N__77694;
    wire N__77693;
    wire N__77692;
    wire N__77691;
    wire N__77690;
    wire N__77689;
    wire N__77688;
    wire N__77685;
    wire N__77682;
    wire N__77675;
    wire N__77668;
    wire N__77659;
    wire N__77654;
    wire N__77647;
    wire N__77642;
    wire N__77639;
    wire N__77636;
    wire N__77627;
    wire N__77624;
    wire N__77621;
    wire N__77620;
    wire N__77619;
    wire N__77618;
    wire N__77617;
    wire N__77616;
    wire N__77615;
    wire N__77614;
    wire N__77613;
    wire N__77612;
    wire N__77611;
    wire N__77610;
    wire N__77609;
    wire N__77608;
    wire N__77605;
    wire N__77598;
    wire N__77591;
    wire N__77590;
    wire N__77587;
    wire N__77584;
    wire N__77583;
    wire N__77580;
    wire N__77577;
    wire N__77576;
    wire N__77575;
    wire N__77568;
    wire N__77559;
    wire N__77548;
    wire N__77539;
    wire N__77532;
    wire N__77525;
    wire N__77518;
    wire N__77515;
    wire N__77512;
    wire N__77507;
    wire N__77498;
    wire N__77489;
    wire N__77480;
    wire N__77473;
    wire N__77466;
    wire N__77459;
    wire N__77450;
    wire N__77441;
    wire N__77438;
    wire N__77427;
    wire N__77420;
    wire N__77415;
    wire N__77408;
    wire N__77401;
    wire N__77392;
    wire N__77383;
    wire N__77378;
    wire N__77373;
    wire N__77366;
    wire N__77343;
    wire N__77318;
    wire N__77317;
    wire N__77316;
    wire N__77315;
    wire N__77314;
    wire N__77313;
    wire N__77312;
    wire N__77311;
    wire N__77310;
    wire N__77309;
    wire N__77308;
    wire N__77305;
    wire N__77304;
    wire N__77303;
    wire N__77302;
    wire N__77301;
    wire N__77298;
    wire N__77297;
    wire N__77296;
    wire N__77295;
    wire N__77294;
    wire N__77293;
    wire N__77292;
    wire N__77287;
    wire N__77284;
    wire N__77283;
    wire N__77282;
    wire N__77281;
    wire N__77280;
    wire N__77275;
    wire N__77274;
    wire N__77273;
    wire N__77272;
    wire N__77271;
    wire N__77268;
    wire N__77265;
    wire N__77262;
    wire N__77259;
    wire N__77258;
    wire N__77257;
    wire N__77256;
    wire N__77255;
    wire N__77254;
    wire N__77253;
    wire N__77252;
    wire N__77251;
    wire N__77250;
    wire N__77249;
    wire N__77248;
    wire N__77247;
    wire N__77246;
    wire N__77245;
    wire N__77244;
    wire N__77243;
    wire N__77242;
    wire N__77241;
    wire N__77240;
    wire N__77239;
    wire N__77238;
    wire N__77237;
    wire N__77236;
    wire N__77235;
    wire N__77234;
    wire N__77231;
    wire N__77222;
    wire N__77219;
    wire N__77214;
    wire N__77205;
    wire N__77202;
    wire N__77201;
    wire N__77200;
    wire N__77199;
    wire N__77198;
    wire N__77197;
    wire N__77196;
    wire N__77193;
    wire N__77192;
    wire N__77191;
    wire N__77190;
    wire N__77189;
    wire N__77188;
    wire N__77187;
    wire N__77186;
    wire N__77185;
    wire N__77184;
    wire N__77183;
    wire N__77182;
    wire N__77181;
    wire N__77176;
    wire N__77175;
    wire N__77174;
    wire N__77173;
    wire N__77172;
    wire N__77171;
    wire N__77166;
    wire N__77165;
    wire N__77164;
    wire N__77161;
    wire N__77152;
    wire N__77151;
    wire N__77150;
    wire N__77149;
    wire N__77148;
    wire N__77147;
    wire N__77146;
    wire N__77145;
    wire N__77144;
    wire N__77143;
    wire N__77142;
    wire N__77141;
    wire N__77140;
    wire N__77137;
    wire N__77132;
    wire N__77129;
    wire N__77126;
    wire N__77125;
    wire N__77124;
    wire N__77123;
    wire N__77122;
    wire N__77121;
    wire N__77120;
    wire N__77119;
    wire N__77118;
    wire N__77117;
    wire N__77116;
    wire N__77115;
    wire N__77114;
    wire N__77109;
    wire N__77100;
    wire N__77093;
    wire N__77088;
    wire N__77081;
    wire N__77074;
    wire N__77073;
    wire N__77072;
    wire N__77071;
    wire N__77070;
    wire N__77069;
    wire N__77068;
    wire N__77067;
    wire N__77066;
    wire N__77065;
    wire N__77062;
    wire N__77055;
    wire N__77048;
    wire N__77039;
    wire N__77034;
    wire N__77027;
    wire N__77020;
    wire N__77017;
    wire N__77010;
    wire N__77003;
    wire N__76998;
    wire N__76995;
    wire N__76988;
    wire N__76985;
    wire N__76982;
    wire N__76979;
    wire N__76978;
    wire N__76977;
    wire N__76970;
    wire N__76967;
    wire N__76966;
    wire N__76965;
    wire N__76960;
    wire N__76957;
    wire N__76954;
    wire N__76947;
    wire N__76938;
    wire N__76937;
    wire N__76936;
    wire N__76935;
    wire N__76934;
    wire N__76933;
    wire N__76932;
    wire N__76931;
    wire N__76930;
    wire N__76929;
    wire N__76928;
    wire N__76927;
    wire N__76926;
    wire N__76925;
    wire N__76914;
    wire N__76913;
    wire N__76912;
    wire N__76911;
    wire N__76910;
    wire N__76909;
    wire N__76904;
    wire N__76899;
    wire N__76890;
    wire N__76879;
    wire N__76872;
    wire N__76865;
    wire N__76858;
    wire N__76851;
    wire N__76838;
    wire N__76831;
    wire N__76822;
    wire N__76811;
    wire N__76802;
    wire N__76797;
    wire N__76792;
    wire N__76787;
    wire N__76784;
    wire N__76775;
    wire N__76762;
    wire N__76753;
    wire N__76746;
    wire N__76743;
    wire N__76732;
    wire N__76723;
    wire N__76704;
    wire N__76679;
    wire N__76676;
    wire N__76673;
    wire N__76670;
    wire N__76667;
    wire N__76664;
    wire N__76661;
    wire N__76658;
    wire N__76655;
    wire N__76652;
    wire N__76649;
    wire N__76648;
    wire N__76645;
    wire N__76642;
    wire N__76637;
    wire N__76636;
    wire N__76635;
    wire N__76634;
    wire N__76633;
    wire N__76626;
    wire N__76625;
    wire N__76624;
    wire N__76623;
    wire N__76620;
    wire N__76619;
    wire N__76618;
    wire N__76617;
    wire N__76616;
    wire N__76613;
    wire N__76610;
    wire N__76609;
    wire N__76608;
    wire N__76607;
    wire N__76606;
    wire N__76605;
    wire N__76604;
    wire N__76603;
    wire N__76602;
    wire N__76601;
    wire N__76600;
    wire N__76597;
    wire N__76594;
    wire N__76593;
    wire N__76592;
    wire N__76591;
    wire N__76588;
    wire N__76587;
    wire N__76586;
    wire N__76585;
    wire N__76584;
    wire N__76583;
    wire N__76580;
    wire N__76579;
    wire N__76576;
    wire N__76575;
    wire N__76574;
    wire N__76573;
    wire N__76572;
    wire N__76571;
    wire N__76570;
    wire N__76569;
    wire N__76566;
    wire N__76563;
    wire N__76560;
    wire N__76559;
    wire N__76554;
    wire N__76551;
    wire N__76546;
    wire N__76541;
    wire N__76536;
    wire N__76535;
    wire N__76534;
    wire N__76533;
    wire N__76532;
    wire N__76531;
    wire N__76530;
    wire N__76529;
    wire N__76528;
    wire N__76527;
    wire N__76526;
    wire N__76523;
    wire N__76522;
    wire N__76519;
    wire N__76516;
    wire N__76513;
    wire N__76510;
    wire N__76507;
    wire N__76504;
    wire N__76501;
    wire N__76500;
    wire N__76499;
    wire N__76498;
    wire N__76493;
    wire N__76486;
    wire N__76485;
    wire N__76484;
    wire N__76483;
    wire N__76482;
    wire N__76481;
    wire N__76480;
    wire N__76479;
    wire N__76476;
    wire N__76475;
    wire N__76474;
    wire N__76473;
    wire N__76472;
    wire N__76471;
    wire N__76470;
    wire N__76467;
    wire N__76464;
    wire N__76463;
    wire N__76462;
    wire N__76461;
    wire N__76460;
    wire N__76459;
    wire N__76458;
    wire N__76455;
    wire N__76454;
    wire N__76449;
    wire N__76448;
    wire N__76447;
    wire N__76446;
    wire N__76441;
    wire N__76434;
    wire N__76429;
    wire N__76424;
    wire N__76421;
    wire N__76414;
    wire N__76411;
    wire N__76406;
    wire N__76405;
    wire N__76404;
    wire N__76403;
    wire N__76396;
    wire N__76391;
    wire N__76388;
    wire N__76381;
    wire N__76378;
    wire N__76375;
    wire N__76374;
    wire N__76373;
    wire N__76372;
    wire N__76369;
    wire N__76362;
    wire N__76357;
    wire N__76354;
    wire N__76351;
    wire N__76350;
    wire N__76349;
    wire N__76346;
    wire N__76341;
    wire N__76336;
    wire N__76331;
    wire N__76326;
    wire N__76323;
    wire N__76322;
    wire N__76321;
    wire N__76318;
    wire N__76313;
    wire N__76310;
    wire N__76305;
    wire N__76302;
    wire N__76299;
    wire N__76294;
    wire N__76293;
    wire N__76292;
    wire N__76291;
    wire N__76288;
    wire N__76287;
    wire N__76286;
    wire N__76277;
    wire N__76274;
    wire N__76273;
    wire N__76272;
    wire N__76271;
    wire N__76270;
    wire N__76269;
    wire N__76268;
    wire N__76265;
    wire N__76264;
    wire N__76263;
    wire N__76262;
    wire N__76261;
    wire N__76258;
    wire N__76251;
    wire N__76248;
    wire N__76241;
    wire N__76232;
    wire N__76225;
    wire N__76222;
    wire N__76215;
    wire N__76210;
    wire N__76203;
    wire N__76192;
    wire N__76185;
    wire N__76174;
    wire N__76173;
    wire N__76168;
    wire N__76159;
    wire N__76152;
    wire N__76145;
    wire N__76142;
    wire N__76139;
    wire N__76136;
    wire N__76131;
    wire N__76128;
    wire N__76123;
    wire N__76118;
    wire N__76113;
    wire N__76110;
    wire N__76103;
    wire N__76098;
    wire N__76089;
    wire N__76074;
    wire N__76071;
    wire N__76062;
    wire N__76059;
    wire N__76028;
    wire N__76025;
    wire N__76022;
    wire N__76019;
    wire N__76016;
    wire N__76015;
    wire N__76012;
    wire N__76011;
    wire N__76010;
    wire N__76009;
    wire N__76008;
    wire N__76005;
    wire N__76004;
    wire N__76003;
    wire N__76002;
    wire N__75997;
    wire N__75996;
    wire N__75995;
    wire N__75994;
    wire N__75993;
    wire N__75992;
    wire N__75991;
    wire N__75990;
    wire N__75987;
    wire N__75986;
    wire N__75985;
    wire N__75984;
    wire N__75983;
    wire N__75980;
    wire N__75977;
    wire N__75974;
    wire N__75973;
    wire N__75970;
    wire N__75969;
    wire N__75968;
    wire N__75967;
    wire N__75966;
    wire N__75965;
    wire N__75964;
    wire N__75963;
    wire N__75962;
    wire N__75961;
    wire N__75960;
    wire N__75959;
    wire N__75956;
    wire N__75955;
    wire N__75954;
    wire N__75951;
    wire N__75950;
    wire N__75947;
    wire N__75942;
    wire N__75941;
    wire N__75940;
    wire N__75939;
    wire N__75938;
    wire N__75935;
    wire N__75934;
    wire N__75933;
    wire N__75932;
    wire N__75929;
    wire N__75926;
    wire N__75923;
    wire N__75920;
    wire N__75919;
    wire N__75918;
    wire N__75917;
    wire N__75916;
    wire N__75915;
    wire N__75914;
    wire N__75913;
    wire N__75912;
    wire N__75911;
    wire N__75910;
    wire N__75909;
    wire N__75908;
    wire N__75907;
    wire N__75906;
    wire N__75905;
    wire N__75904;
    wire N__75903;
    wire N__75902;
    wire N__75901;
    wire N__75900;
    wire N__75899;
    wire N__75896;
    wire N__75893;
    wire N__75892;
    wire N__75891;
    wire N__75890;
    wire N__75889;
    wire N__75888;
    wire N__75887;
    wire N__75886;
    wire N__75885;
    wire N__75882;
    wire N__75881;
    wire N__75880;
    wire N__75879;
    wire N__75876;
    wire N__75871;
    wire N__75868;
    wire N__75865;
    wire N__75860;
    wire N__75857;
    wire N__75856;
    wire N__75853;
    wire N__75852;
    wire N__75851;
    wire N__75848;
    wire N__75847;
    wire N__75846;
    wire N__75843;
    wire N__75840;
    wire N__75839;
    wire N__75836;
    wire N__75833;
    wire N__75832;
    wire N__75831;
    wire N__75830;
    wire N__75829;
    wire N__75828;
    wire N__75825;
    wire N__75822;
    wire N__75821;
    wire N__75818;
    wire N__75817;
    wire N__75816;
    wire N__75815;
    wire N__75814;
    wire N__75811;
    wire N__75810;
    wire N__75809;
    wire N__75808;
    wire N__75805;
    wire N__75804;
    wire N__75801;
    wire N__75800;
    wire N__75799;
    wire N__75796;
    wire N__75795;
    wire N__75792;
    wire N__75791;
    wire N__75790;
    wire N__75789;
    wire N__75786;
    wire N__75781;
    wire N__75770;
    wire N__75763;
    wire N__75754;
    wire N__75751;
    wire N__75750;
    wire N__75747;
    wire N__75746;
    wire N__75743;
    wire N__75740;
    wire N__75737;
    wire N__75736;
    wire N__75733;
    wire N__75730;
    wire N__75727;
    wire N__75726;
    wire N__75725;
    wire N__75722;
    wire N__75721;
    wire N__75720;
    wire N__75719;
    wire N__75718;
    wire N__75715;
    wire N__75712;
    wire N__75711;
    wire N__75710;
    wire N__75709;
    wire N__75708;
    wire N__75705;
    wire N__75702;
    wire N__75695;
    wire N__75692;
    wire N__75689;
    wire N__75688;
    wire N__75685;
    wire N__75684;
    wire N__75681;
    wire N__75680;
    wire N__75677;
    wire N__75676;
    wire N__75673;
    wire N__75672;
    wire N__75671;
    wire N__75670;
    wire N__75669;
    wire N__75668;
    wire N__75665;
    wire N__75660;
    wire N__75659;
    wire N__75656;
    wire N__75655;
    wire N__75654;
    wire N__75653;
    wire N__75650;
    wire N__75647;
    wire N__75646;
    wire N__75645;
    wire N__75642;
    wire N__75639;
    wire N__75638;
    wire N__75637;
    wire N__75636;
    wire N__75635;
    wire N__75632;
    wire N__75631;
    wire N__75630;
    wire N__75627;
    wire N__75620;
    wire N__75619;
    wire N__75616;
    wire N__75615;
    wire N__75614;
    wire N__75613;
    wire N__75612;
    wire N__75611;
    wire N__75606;
    wire N__75599;
    wire N__75598;
    wire N__75597;
    wire N__75594;
    wire N__75587;
    wire N__75580;
    wire N__75577;
    wire N__75570;
    wire N__75561;
    wire N__75556;
    wire N__75551;
    wire N__75546;
    wire N__75541;
    wire N__75540;
    wire N__75539;
    wire N__75538;
    wire N__75535;
    wire N__75534;
    wire N__75533;
    wire N__75530;
    wire N__75529;
    wire N__75528;
    wire N__75527;
    wire N__75526;
    wire N__75521;
    wire N__75516;
    wire N__75513;
    wire N__75502;
    wire N__75501;
    wire N__75500;
    wire N__75499;
    wire N__75496;
    wire N__75493;
    wire N__75490;
    wire N__75483;
    wire N__75474;
    wire N__75467;
    wire N__75460;
    wire N__75453;
    wire N__75446;
    wire N__75439;
    wire N__75430;
    wire N__75425;
    wire N__75424;
    wire N__75423;
    wire N__75422;
    wire N__75419;
    wire N__75416;
    wire N__75413;
    wire N__75410;
    wire N__75407;
    wire N__75404;
    wire N__75401;
    wire N__75394;
    wire N__75385;
    wire N__75384;
    wire N__75383;
    wire N__75380;
    wire N__75377;
    wire N__75366;
    wire N__75361;
    wire N__75348;
    wire N__75339;
    wire N__75336;
    wire N__75329;
    wire N__75320;
    wire N__75317;
    wire N__75314;
    wire N__75311;
    wire N__75308;
    wire N__75307;
    wire N__75306;
    wire N__75305;
    wire N__75304;
    wire N__75303;
    wire N__75300;
    wire N__75299;
    wire N__75296;
    wire N__75293;
    wire N__75292;
    wire N__75291;
    wire N__75288;
    wire N__75287;
    wire N__75284;
    wire N__75283;
    wire N__75280;
    wire N__75277;
    wire N__75272;
    wire N__75263;
    wire N__75258;
    wire N__75249;
    wire N__75248;
    wire N__75247;
    wire N__75244;
    wire N__75243;
    wire N__75240;
    wire N__75237;
    wire N__75236;
    wire N__75235;
    wire N__75234;
    wire N__75231;
    wire N__75224;
    wire N__75215;
    wire N__75212;
    wire N__75205;
    wire N__75196;
    wire N__75179;
    wire N__75172;
    wire N__75161;
    wire N__75158;
    wire N__75151;
    wire N__75144;
    wire N__75137;
    wire N__75126;
    wire N__75123;
    wire N__75118;
    wire N__75109;
    wire N__75106;
    wire N__75101;
    wire N__75090;
    wire N__75083;
    wire N__75074;
    wire N__75061;
    wire N__75050;
    wire N__75041;
    wire N__75034;
    wire N__75021;
    wire N__75010;
    wire N__75003;
    wire N__74978;
    wire N__74975;
    wire N__74972;
    wire N__74969;
    wire N__74966;
    wire N__74963;
    wire N__74962;
    wire N__74959;
    wire N__74956;
    wire N__74953;
    wire N__74950;
    wire N__74945;
    wire N__74942;
    wire N__74939;
    wire N__74936;
    wire N__74933;
    wire N__74930;
    wire N__74927;
    wire N__74924;
    wire N__74921;
    wire N__74918;
    wire N__74915;
    wire N__74912;
    wire N__74909;
    wire N__74906;
    wire N__74903;
    wire N__74902;
    wire N__74899;
    wire N__74896;
    wire N__74895;
    wire N__74894;
    wire N__74891;
    wire N__74890;
    wire N__74889;
    wire N__74888;
    wire N__74887;
    wire N__74886;
    wire N__74883;
    wire N__74882;
    wire N__74879;
    wire N__74876;
    wire N__74873;
    wire N__74870;
    wire N__74867;
    wire N__74864;
    wire N__74861;
    wire N__74860;
    wire N__74857;
    wire N__74856;
    wire N__74855;
    wire N__74854;
    wire N__74853;
    wire N__74850;
    wire N__74847;
    wire N__74844;
    wire N__74841;
    wire N__74838;
    wire N__74835;
    wire N__74834;
    wire N__74833;
    wire N__74832;
    wire N__74827;
    wire N__74826;
    wire N__74825;
    wire N__74824;
    wire N__74817;
    wire N__74816;
    wire N__74815;
    wire N__74812;
    wire N__74809;
    wire N__74804;
    wire N__74801;
    wire N__74798;
    wire N__74793;
    wire N__74788;
    wire N__74785;
    wire N__74782;
    wire N__74779;
    wire N__74778;
    wire N__74775;
    wire N__74772;
    wire N__74771;
    wire N__74768;
    wire N__74765;
    wire N__74762;
    wire N__74759;
    wire N__74756;
    wire N__74753;
    wire N__74750;
    wire N__74739;
    wire N__74736;
    wire N__74733;
    wire N__74730;
    wire N__74727;
    wire N__74724;
    wire N__74715;
    wire N__74712;
    wire N__74709;
    wire N__74706;
    wire N__74703;
    wire N__74700;
    wire N__74697;
    wire N__74694;
    wire N__74691;
    wire N__74686;
    wire N__74683;
    wire N__74682;
    wire N__74681;
    wire N__74674;
    wire N__74671;
    wire N__74666;
    wire N__74663;
    wire N__74658;
    wire N__74655;
    wire N__74652;
    wire N__74649;
    wire N__74646;
    wire N__74643;
    wire N__74636;
    wire N__74629;
    wire N__74618;
    wire N__74615;
    wire N__74612;
    wire N__74609;
    wire N__74608;
    wire N__74607;
    wire N__74604;
    wire N__74603;
    wire N__74600;
    wire N__74597;
    wire N__74596;
    wire N__74593;
    wire N__74590;
    wire N__74587;
    wire N__74584;
    wire N__74581;
    wire N__74578;
    wire N__74575;
    wire N__74572;
    wire N__74571;
    wire N__74570;
    wire N__74569;
    wire N__74566;
    wire N__74563;
    wire N__74560;
    wire N__74555;
    wire N__74548;
    wire N__74545;
    wire N__74542;
    wire N__74539;
    wire N__74528;
    wire N__74525;
    wire N__74524;
    wire N__74521;
    wire N__74518;
    wire N__74515;
    wire N__74512;
    wire N__74507;
    wire N__74504;
    wire N__74501;
    wire N__74498;
    wire N__74495;
    wire N__74492;
    wire N__74491;
    wire N__74490;
    wire N__74489;
    wire N__74488;
    wire N__74487;
    wire N__74484;
    wire N__74481;
    wire N__74480;
    wire N__74477;
    wire N__74474;
    wire N__74471;
    wire N__74468;
    wire N__74465;
    wire N__74462;
    wire N__74459;
    wire N__74454;
    wire N__74451;
    wire N__74448;
    wire N__74447;
    wire N__74444;
    wire N__74439;
    wire N__74434;
    wire N__74431;
    wire N__74428;
    wire N__74423;
    wire N__74416;
    wire N__74411;
    wire N__74410;
    wire N__74407;
    wire N__74406;
    wire N__74403;
    wire N__74400;
    wire N__74397;
    wire N__74394;
    wire N__74391;
    wire N__74386;
    wire N__74383;
    wire N__74378;
    wire N__74375;
    wire N__74372;
    wire N__74369;
    wire N__74366;
    wire N__74363;
    wire N__74360;
    wire N__74357;
    wire N__74354;
    wire N__74351;
    wire N__74348;
    wire N__74345;
    wire N__74342;
    wire N__74339;
    wire N__74336;
    wire N__74333;
    wire N__74330;
    wire N__74329;
    wire N__74324;
    wire N__74321;
    wire N__74318;
    wire N__74315;
    wire N__74312;
    wire N__74309;
    wire N__74306;
    wire N__74303;
    wire N__74300;
    wire N__74297;
    wire N__74294;
    wire N__74291;
    wire N__74288;
    wire N__74285;
    wire N__74282;
    wire N__74279;
    wire N__74276;
    wire N__74273;
    wire N__74270;
    wire N__74267;
    wire N__74264;
    wire N__74261;
    wire N__74258;
    wire N__74255;
    wire N__74252;
    wire N__74249;
    wire N__74246;
    wire N__74243;
    wire N__74240;
    wire N__74239;
    wire N__74236;
    wire N__74233;
    wire N__74230;
    wire N__74225;
    wire N__74222;
    wire N__74219;
    wire N__74216;
    wire N__74213;
    wire N__74212;
    wire N__74207;
    wire N__74204;
    wire N__74201;
    wire N__74198;
    wire N__74195;
    wire N__74192;
    wire N__74189;
    wire N__74186;
    wire N__74185;
    wire N__74182;
    wire N__74179;
    wire N__74176;
    wire N__74171;
    wire N__74168;
    wire N__74165;
    wire N__74162;
    wire N__74159;
    wire N__74156;
    wire N__74153;
    wire N__74150;
    wire N__74147;
    wire N__74144;
    wire N__74141;
    wire N__74138;
    wire N__74135;
    wire N__74132;
    wire N__74129;
    wire N__74126;
    wire N__74125;
    wire N__74122;
    wire N__74119;
    wire N__74116;
    wire N__74111;
    wire N__74108;
    wire N__74105;
    wire N__74102;
    wire N__74099;
    wire N__74096;
    wire N__74093;
    wire N__74090;
    wire N__74087;
    wire N__74084;
    wire N__74081;
    wire N__74078;
    wire N__74075;
    wire N__74072;
    wire N__74071;
    wire N__74070;
    wire N__74069;
    wire N__74068;
    wire N__74067;
    wire N__74066;
    wire N__74065;
    wire N__74062;
    wire N__74061;
    wire N__74058;
    wire N__74053;
    wire N__74050;
    wire N__74045;
    wire N__74042;
    wire N__74039;
    wire N__74038;
    wire N__74037;
    wire N__74034;
    wire N__74031;
    wire N__74024;
    wire N__74023;
    wire N__74020;
    wire N__74017;
    wire N__74012;
    wire N__74011;
    wire N__74008;
    wire N__74007;
    wire N__74004;
    wire N__74001;
    wire N__73998;
    wire N__73997;
    wire N__73994;
    wire N__73989;
    wire N__73986;
    wire N__73983;
    wire N__73980;
    wire N__73977;
    wire N__73972;
    wire N__73969;
    wire N__73964;
    wire N__73959;
    wire N__73946;
    wire N__73945;
    wire N__73942;
    wire N__73937;
    wire N__73934;
    wire N__73931;
    wire N__73928;
    wire N__73925;
    wire N__73922;
    wire N__73919;
    wire N__73918;
    wire N__73915;
    wire N__73912;
    wire N__73911;
    wire N__73906;
    wire N__73905;
    wire N__73902;
    wire N__73899;
    wire N__73896;
    wire N__73893;
    wire N__73892;
    wire N__73891;
    wire N__73886;
    wire N__73883;
    wire N__73880;
    wire N__73877;
    wire N__73874;
    wire N__73873;
    wire N__73870;
    wire N__73867;
    wire N__73864;
    wire N__73861;
    wire N__73858;
    wire N__73857;
    wire N__73852;
    wire N__73849;
    wire N__73846;
    wire N__73841;
    wire N__73838;
    wire N__73829;
    wire N__73826;
    wire N__73823;
    wire N__73820;
    wire N__73817;
    wire N__73814;
    wire N__73813;
    wire N__73812;
    wire N__73811;
    wire N__73810;
    wire N__73809;
    wire N__73808;
    wire N__73805;
    wire N__73800;
    wire N__73797;
    wire N__73794;
    wire N__73791;
    wire N__73788;
    wire N__73787;
    wire N__73784;
    wire N__73781;
    wire N__73778;
    wire N__73773;
    wire N__73770;
    wire N__73767;
    wire N__73766;
    wire N__73761;
    wire N__73752;
    wire N__73749;
    wire N__73742;
    wire N__73741;
    wire N__73740;
    wire N__73737;
    wire N__73734;
    wire N__73731;
    wire N__73730;
    wire N__73729;
    wire N__73728;
    wire N__73725;
    wire N__73722;
    wire N__73721;
    wire N__73720;
    wire N__73719;
    wire N__73716;
    wire N__73713;
    wire N__73712;
    wire N__73707;
    wire N__73702;
    wire N__73697;
    wire N__73694;
    wire N__73691;
    wire N__73688;
    wire N__73687;
    wire N__73686;
    wire N__73683;
    wire N__73680;
    wire N__73679;
    wire N__73678;
    wire N__73677;
    wire N__73672;
    wire N__73669;
    wire N__73668;
    wire N__73665;
    wire N__73662;
    wire N__73661;
    wire N__73658;
    wire N__73655;
    wire N__73652;
    wire N__73649;
    wire N__73642;
    wire N__73637;
    wire N__73636;
    wire N__73633;
    wire N__73628;
    wire N__73627;
    wire N__73624;
    wire N__73619;
    wire N__73614;
    wire N__73611;
    wire N__73608;
    wire N__73605;
    wire N__73600;
    wire N__73595;
    wire N__73588;
    wire N__73585;
    wire N__73574;
    wire N__73573;
    wire N__73572;
    wire N__73569;
    wire N__73566;
    wire N__73565;
    wire N__73562;
    wire N__73559;
    wire N__73554;
    wire N__73553;
    wire N__73552;
    wire N__73549;
    wire N__73546;
    wire N__73543;
    wire N__73542;
    wire N__73539;
    wire N__73536;
    wire N__73533;
    wire N__73530;
    wire N__73527;
    wire N__73524;
    wire N__73519;
    wire N__73516;
    wire N__73505;
    wire N__73504;
    wire N__73503;
    wire N__73498;
    wire N__73495;
    wire N__73492;
    wire N__73491;
    wire N__73488;
    wire N__73485;
    wire N__73482;
    wire N__73475;
    wire N__73472;
    wire N__73469;
    wire N__73466;
    wire N__73463;
    wire N__73460;
    wire N__73457;
    wire N__73454;
    wire N__73451;
    wire N__73448;
    wire N__73445;
    wire N__73442;
    wire N__73439;
    wire N__73436;
    wire N__73433;
    wire N__73430;
    wire N__73427;
    wire N__73424;
    wire N__73421;
    wire N__73418;
    wire N__73415;
    wire N__73412;
    wire N__73409;
    wire N__73406;
    wire N__73403;
    wire N__73400;
    wire N__73397;
    wire N__73394;
    wire N__73391;
    wire N__73388;
    wire N__73385;
    wire N__73382;
    wire N__73379;
    wire N__73376;
    wire N__73373;
    wire N__73370;
    wire N__73367;
    wire N__73364;
    wire N__73361;
    wire N__73358;
    wire N__73355;
    wire N__73352;
    wire N__73349;
    wire N__73348;
    wire N__73345;
    wire N__73342;
    wire N__73339;
    wire N__73336;
    wire N__73333;
    wire N__73330;
    wire N__73327;
    wire N__73324;
    wire N__73319;
    wire N__73316;
    wire N__73313;
    wire N__73310;
    wire N__73307;
    wire N__73304;
    wire N__73303;
    wire N__73302;
    wire N__73299;
    wire N__73294;
    wire N__73293;
    wire N__73292;
    wire N__73291;
    wire N__73290;
    wire N__73287;
    wire N__73286;
    wire N__73283;
    wire N__73282;
    wire N__73281;
    wire N__73280;
    wire N__73279;
    wire N__73278;
    wire N__73277;
    wire N__73276;
    wire N__73275;
    wire N__73274;
    wire N__73273;
    wire N__73272;
    wire N__73271;
    wire N__73270;
    wire N__73269;
    wire N__73268;
    wire N__73267;
    wire N__73266;
    wire N__73265;
    wire N__73264;
    wire N__73263;
    wire N__73262;
    wire N__73261;
    wire N__73260;
    wire N__73259;
    wire N__73258;
    wire N__73257;
    wire N__73256;
    wire N__73255;
    wire N__73254;
    wire N__73253;
    wire N__73252;
    wire N__73251;
    wire N__73250;
    wire N__73249;
    wire N__73248;
    wire N__73247;
    wire N__73246;
    wire N__73245;
    wire N__73244;
    wire N__73243;
    wire N__73242;
    wire N__73241;
    wire N__73240;
    wire N__73239;
    wire N__73238;
    wire N__73237;
    wire N__73236;
    wire N__73235;
    wire N__73234;
    wire N__73233;
    wire N__73232;
    wire N__73231;
    wire N__73230;
    wire N__73229;
    wire N__73228;
    wire N__73227;
    wire N__73226;
    wire N__73225;
    wire N__73224;
    wire N__73223;
    wire N__73222;
    wire N__73221;
    wire N__73220;
    wire N__73219;
    wire N__73218;
    wire N__73217;
    wire N__73216;
    wire N__73215;
    wire N__73214;
    wire N__73213;
    wire N__73212;
    wire N__73211;
    wire N__73210;
    wire N__73209;
    wire N__73208;
    wire N__73207;
    wire N__73206;
    wire N__73205;
    wire N__73204;
    wire N__73203;
    wire N__73202;
    wire N__73201;
    wire N__73200;
    wire N__73199;
    wire N__73198;
    wire N__73197;
    wire N__73196;
    wire N__73195;
    wire N__73194;
    wire N__73193;
    wire N__73192;
    wire N__73191;
    wire N__73190;
    wire N__73189;
    wire N__73188;
    wire N__73187;
    wire N__73186;
    wire N__73185;
    wire N__73184;
    wire N__73183;
    wire N__73182;
    wire N__73181;
    wire N__73180;
    wire N__73179;
    wire N__73178;
    wire N__73177;
    wire N__73176;
    wire N__73175;
    wire N__73174;
    wire N__73173;
    wire N__73172;
    wire N__73171;
    wire N__73170;
    wire N__73169;
    wire N__73168;
    wire N__73167;
    wire N__73166;
    wire N__73165;
    wire N__73164;
    wire N__73163;
    wire N__73162;
    wire N__73161;
    wire N__73160;
    wire N__73159;
    wire N__73158;
    wire N__73157;
    wire N__73156;
    wire N__73155;
    wire N__73154;
    wire N__73153;
    wire N__73152;
    wire N__73151;
    wire N__73150;
    wire N__73149;
    wire N__73148;
    wire N__73147;
    wire N__73146;
    wire N__73145;
    wire N__73144;
    wire N__73143;
    wire N__73142;
    wire N__73141;
    wire N__73140;
    wire N__73139;
    wire N__73138;
    wire N__72833;
    wire N__72830;
    wire N__72827;
    wire N__72824;
    wire N__72821;
    wire N__72818;
    wire N__72815;
    wire N__72812;
    wire N__72809;
    wire N__72806;
    wire N__72803;
    wire N__72800;
    wire N__72797;
    wire N__72794;
    wire N__72791;
    wire N__72790;
    wire N__72789;
    wire N__72786;
    wire N__72785;
    wire N__72784;
    wire N__72781;
    wire N__72778;
    wire N__72777;
    wire N__72776;
    wire N__72775;
    wire N__72774;
    wire N__72773;
    wire N__72772;
    wire N__72771;
    wire N__72770;
    wire N__72769;
    wire N__72768;
    wire N__72761;
    wire N__72752;
    wire N__72749;
    wire N__72746;
    wire N__72743;
    wire N__72742;
    wire N__72741;
    wire N__72738;
    wire N__72737;
    wire N__72732;
    wire N__72731;
    wire N__72730;
    wire N__72729;
    wire N__72728;
    wire N__72727;
    wire N__72726;
    wire N__72725;
    wire N__72724;
    wire N__72723;
    wire N__72722;
    wire N__72721;
    wire N__72720;
    wire N__72717;
    wire N__72714;
    wire N__72713;
    wire N__72712;
    wire N__72707;
    wire N__72704;
    wire N__72699;
    wire N__72698;
    wire N__72697;
    wire N__72696;
    wire N__72695;
    wire N__72694;
    wire N__72693;
    wire N__72692;
    wire N__72691;
    wire N__72690;
    wire N__72689;
    wire N__72688;
    wire N__72685;
    wire N__72684;
    wire N__72683;
    wire N__72682;
    wire N__72681;
    wire N__72676;
    wire N__72673;
    wire N__72672;
    wire N__72669;
    wire N__72666;
    wire N__72657;
    wire N__72656;
    wire N__72655;
    wire N__72652;
    wire N__72649;
    wire N__72648;
    wire N__72637;
    wire N__72630;
    wire N__72627;
    wire N__72626;
    wire N__72619;
    wire N__72618;
    wire N__72615;
    wire N__72612;
    wire N__72609;
    wire N__72608;
    wire N__72607;
    wire N__72606;
    wire N__72603;
    wire N__72600;
    wire N__72597;
    wire N__72588;
    wire N__72583;
    wire N__72580;
    wire N__72577;
    wire N__72572;
    wire N__72567;
    wire N__72564;
    wire N__72563;
    wire N__72560;
    wire N__72557;
    wire N__72554;
    wire N__72549;
    wire N__72546;
    wire N__72541;
    wire N__72538;
    wire N__72535;
    wire N__72532;
    wire N__72529;
    wire N__72526;
    wire N__72523;
    wire N__72520;
    wire N__72515;
    wire N__72512;
    wire N__72511;
    wire N__72508;
    wire N__72505;
    wire N__72504;
    wire N__72503;
    wire N__72500;
    wire N__72495;
    wire N__72490;
    wire N__72485;
    wire N__72480;
    wire N__72475;
    wire N__72470;
    wire N__72461;
    wire N__72454;
    wire N__72451;
    wire N__72446;
    wire N__72439;
    wire N__72436;
    wire N__72433;
    wire N__72430;
    wire N__72427;
    wire N__72424;
    wire N__72415;
    wire N__72404;
    wire N__72383;
    wire N__72380;
    wire N__72377;
    wire N__72376;
    wire N__72373;
    wire N__72370;
    wire N__72367;
    wire N__72364;
    wire N__72361;
    wire N__72358;
    wire N__72353;
    wire N__72352;
    wire N__72349;
    wire N__72348;
    wire N__72345;
    wire N__72342;
    wire N__72339;
    wire N__72336;
    wire N__72331;
    wire N__72328;
    wire N__72325;
    wire N__72320;
    wire N__72319;
    wire N__72318;
    wire N__72317;
    wire N__72316;
    wire N__72315;
    wire N__72312;
    wire N__72311;
    wire N__72308;
    wire N__72307;
    wire N__72306;
    wire N__72305;
    wire N__72304;
    wire N__72301;
    wire N__72300;
    wire N__72299;
    wire N__72298;
    wire N__72297;
    wire N__72294;
    wire N__72293;
    wire N__72290;
    wire N__72289;
    wire N__72288;
    wire N__72285;
    wire N__72284;
    wire N__72281;
    wire N__72274;
    wire N__72273;
    wire N__72272;
    wire N__72271;
    wire N__72268;
    wire N__72265;
    wire N__72264;
    wire N__72263;
    wire N__72262;
    wire N__72261;
    wire N__72260;
    wire N__72257;
    wire N__72256;
    wire N__72253;
    wire N__72252;
    wire N__72251;
    wire N__72250;
    wire N__72249;
    wire N__72248;
    wire N__72247;
    wire N__72244;
    wire N__72239;
    wire N__72236;
    wire N__72231;
    wire N__72228;
    wire N__72227;
    wire N__72226;
    wire N__72225;
    wire N__72224;
    wire N__72223;
    wire N__72222;
    wire N__72221;
    wire N__72220;
    wire N__72217;
    wire N__72214;
    wire N__72213;
    wire N__72212;
    wire N__72209;
    wire N__72206;
    wire N__72201;
    wire N__72198;
    wire N__72195;
    wire N__72194;
    wire N__72193;
    wire N__72192;
    wire N__72191;
    wire N__72190;
    wire N__72189;
    wire N__72188;
    wire N__72185;
    wire N__72182;
    wire N__72181;
    wire N__72180;
    wire N__72179;
    wire N__72178;
    wire N__72177;
    wire N__72176;
    wire N__72171;
    wire N__72166;
    wire N__72161;
    wire N__72158;
    wire N__72155;
    wire N__72152;
    wire N__72149;
    wire N__72146;
    wire N__72141;
    wire N__72140;
    wire N__72137;
    wire N__72134;
    wire N__72133;
    wire N__72132;
    wire N__72131;
    wire N__72130;
    wire N__72129;
    wire N__72128;
    wire N__72123;
    wire N__72118;
    wire N__72115;
    wire N__72110;
    wire N__72105;
    wire N__72104;
    wire N__72103;
    wire N__72102;
    wire N__72101;
    wire N__72100;
    wire N__72097;
    wire N__72092;
    wire N__72081;
    wire N__72078;
    wire N__72075;
    wire N__72068;
    wire N__72061;
    wire N__72052;
    wire N__72047;
    wire N__72044;
    wire N__72033;
    wire N__72026;
    wire N__72013;
    wire N__72010;
    wire N__72009;
    wire N__72008;
    wire N__72005;
    wire N__72002;
    wire N__71997;
    wire N__71994;
    wire N__71987;
    wire N__71976;
    wire N__71973;
    wire N__71968;
    wire N__71963;
    wire N__71960;
    wire N__71951;
    wire N__71948;
    wire N__71935;
    wire N__71932;
    wire N__71925;
    wire N__71922;
    wire N__71915;
    wire N__71910;
    wire N__71895;
    wire N__71892;
    wire N__71879;
    wire N__71876;
    wire N__71875;
    wire N__71874;
    wire N__71873;
    wire N__71872;
    wire N__71871;
    wire N__71870;
    wire N__71869;
    wire N__71868;
    wire N__71867;
    wire N__71866;
    wire N__71863;
    wire N__71860;
    wire N__71855;
    wire N__71854;
    wire N__71853;
    wire N__71852;
    wire N__71849;
    wire N__71842;
    wire N__71835;
    wire N__71832;
    wire N__71831;
    wire N__71830;
    wire N__71829;
    wire N__71828;
    wire N__71827;
    wire N__71826;
    wire N__71825;
    wire N__71824;
    wire N__71823;
    wire N__71822;
    wire N__71821;
    wire N__71820;
    wire N__71819;
    wire N__71816;
    wire N__71813;
    wire N__71810;
    wire N__71807;
    wire N__71806;
    wire N__71805;
    wire N__71804;
    wire N__71803;
    wire N__71802;
    wire N__71799;
    wire N__71792;
    wire N__71789;
    wire N__71786;
    wire N__71783;
    wire N__71776;
    wire N__71765;
    wire N__71762;
    wire N__71759;
    wire N__71758;
    wire N__71755;
    wire N__71752;
    wire N__71749;
    wire N__71746;
    wire N__71745;
    wire N__71742;
    wire N__71739;
    wire N__71730;
    wire N__71727;
    wire N__71722;
    wire N__71715;
    wire N__71712;
    wire N__71709;
    wire N__71706;
    wire N__71701;
    wire N__71698;
    wire N__71693;
    wire N__71690;
    wire N__71683;
    wire N__71676;
    wire N__71657;
    wire N__71654;
    wire N__71651;
    wire N__71648;
    wire N__71645;
    wire N__71642;
    wire N__71639;
    wire N__71636;
    wire N__71633;
    wire N__71630;
    wire N__71627;
    wire N__71624;
    wire N__71621;
    wire N__71618;
    wire N__71615;
    wire N__71612;
    wire N__71609;
    wire N__71606;
    wire N__71603;
    wire N__71600;
    wire N__71597;
    wire N__71594;
    wire N__71591;
    wire N__71588;
    wire N__71585;
    wire N__71582;
    wire N__71579;
    wire N__71578;
    wire N__71573;
    wire N__71570;
    wire N__71567;
    wire N__71564;
    wire N__71561;
    wire N__71558;
    wire N__71555;
    wire N__71554;
    wire N__71553;
    wire N__71550;
    wire N__71547;
    wire N__71544;
    wire N__71539;
    wire N__71536;
    wire N__71533;
    wire N__71530;
    wire N__71527;
    wire N__71522;
    wire N__71519;
    wire N__71516;
    wire N__71515;
    wire N__71512;
    wire N__71509;
    wire N__71504;
    wire N__71501;
    wire N__71500;
    wire N__71495;
    wire N__71492;
    wire N__71491;
    wire N__71490;
    wire N__71487;
    wire N__71484;
    wire N__71481;
    wire N__71478;
    wire N__71471;
    wire N__71470;
    wire N__71469;
    wire N__71468;
    wire N__71467;
    wire N__71464;
    wire N__71463;
    wire N__71460;
    wire N__71455;
    wire N__71454;
    wire N__71453;
    wire N__71452;
    wire N__71451;
    wire N__71450;
    wire N__71449;
    wire N__71448;
    wire N__71445;
    wire N__71442;
    wire N__71441;
    wire N__71440;
    wire N__71437;
    wire N__71436;
    wire N__71435;
    wire N__71432;
    wire N__71429;
    wire N__71426;
    wire N__71425;
    wire N__71424;
    wire N__71423;
    wire N__71418;
    wire N__71411;
    wire N__71410;
    wire N__71407;
    wire N__71402;
    wire N__71401;
    wire N__71400;
    wire N__71399;
    wire N__71396;
    wire N__71395;
    wire N__71394;
    wire N__71391;
    wire N__71388;
    wire N__71385;
    wire N__71384;
    wire N__71381;
    wire N__71380;
    wire N__71377;
    wire N__71372;
    wire N__71367;
    wire N__71364;
    wire N__71361;
    wire N__71358;
    wire N__71353;
    wire N__71350;
    wire N__71347;
    wire N__71344;
    wire N__71341;
    wire N__71338;
    wire N__71333;
    wire N__71330;
    wire N__71327;
    wire N__71324;
    wire N__71321;
    wire N__71320;
    wire N__71315;
    wire N__71314;
    wire N__71309;
    wire N__71304;
    wire N__71297;
    wire N__71292;
    wire N__71289;
    wire N__71282;
    wire N__71279;
    wire N__71274;
    wire N__71269;
    wire N__71266;
    wire N__71263;
    wire N__71260;
    wire N__71257;
    wire N__71254;
    wire N__71251;
    wire N__71248;
    wire N__71245;
    wire N__71236;
    wire N__71219;
    wire N__71216;
    wire N__71215;
    wire N__71214;
    wire N__71213;
    wire N__71212;
    wire N__71211;
    wire N__71208;
    wire N__71207;
    wire N__71204;
    wire N__71201;
    wire N__71200;
    wire N__71199;
    wire N__71198;
    wire N__71197;
    wire N__71194;
    wire N__71193;
    wire N__71190;
    wire N__71189;
    wire N__71186;
    wire N__71183;
    wire N__71180;
    wire N__71177;
    wire N__71176;
    wire N__71173;
    wire N__71170;
    wire N__71167;
    wire N__71164;
    wire N__71163;
    wire N__71160;
    wire N__71157;
    wire N__71154;
    wire N__71151;
    wire N__71148;
    wire N__71145;
    wire N__71140;
    wire N__71137;
    wire N__71134;
    wire N__71131;
    wire N__71128;
    wire N__71125;
    wire N__71122;
    wire N__71119;
    wire N__71116;
    wire N__71113;
    wire N__71110;
    wire N__71105;
    wire N__71102;
    wire N__71097;
    wire N__71094;
    wire N__71089;
    wire N__71084;
    wire N__71081;
    wire N__71076;
    wire N__71071;
    wire N__71066;
    wire N__71063;
    wire N__71060;
    wire N__71057;
    wire N__71052;
    wire N__71049;
    wire N__71046;
    wire N__71043;
    wire N__71038;
    wire N__71035;
    wire N__71030;
    wire N__71021;
    wire N__71020;
    wire N__71019;
    wire N__71012;
    wire N__71009;
    wire N__71008;
    wire N__71007;
    wire N__71006;
    wire N__70997;
    wire N__70994;
    wire N__70993;
    wire N__70990;
    wire N__70987;
    wire N__70986;
    wire N__70983;
    wire N__70980;
    wire N__70977;
    wire N__70974;
    wire N__70971;
    wire N__70968;
    wire N__70965;
    wire N__70962;
    wire N__70959;
    wire N__70956;
    wire N__70953;
    wire N__70948;
    wire N__70943;
    wire N__70942;
    wire N__70941;
    wire N__70940;
    wire N__70937;
    wire N__70936;
    wire N__70935;
    wire N__70932;
    wire N__70931;
    wire N__70922;
    wire N__70915;
    wire N__70914;
    wire N__70913;
    wire N__70908;
    wire N__70905;
    wire N__70902;
    wire N__70897;
    wire N__70892;
    wire N__70891;
    wire N__70890;
    wire N__70889;
    wire N__70888;
    wire N__70887;
    wire N__70884;
    wire N__70883;
    wire N__70882;
    wire N__70875;
    wire N__70866;
    wire N__70865;
    wire N__70862;
    wire N__70859;
    wire N__70856;
    wire N__70853;
    wire N__70844;
    wire N__70841;
    wire N__70838;
    wire N__70835;
    wire N__70832;
    wire N__70829;
    wire N__70828;
    wire N__70825;
    wire N__70822;
    wire N__70819;
    wire N__70816;
    wire N__70815;
    wire N__70812;
    wire N__70809;
    wire N__70806;
    wire N__70799;
    wire N__70798;
    wire N__70797;
    wire N__70796;
    wire N__70795;
    wire N__70794;
    wire N__70791;
    wire N__70790;
    wire N__70789;
    wire N__70788;
    wire N__70787;
    wire N__70786;
    wire N__70785;
    wire N__70782;
    wire N__70779;
    wire N__70776;
    wire N__70773;
    wire N__70770;
    wire N__70767;
    wire N__70766;
    wire N__70765;
    wire N__70764;
    wire N__70763;
    wire N__70762;
    wire N__70761;
    wire N__70760;
    wire N__70759;
    wire N__70758;
    wire N__70757;
    wire N__70756;
    wire N__70755;
    wire N__70754;
    wire N__70751;
    wire N__70746;
    wire N__70733;
    wire N__70730;
    wire N__70727;
    wire N__70724;
    wire N__70723;
    wire N__70722;
    wire N__70721;
    wire N__70718;
    wire N__70715;
    wire N__70712;
    wire N__70711;
    wire N__70710;
    wire N__70709;
    wire N__70708;
    wire N__70703;
    wire N__70700;
    wire N__70693;
    wire N__70690;
    wire N__70683;
    wire N__70678;
    wire N__70671;
    wire N__70668;
    wire N__70661;
    wire N__70646;
    wire N__70643;
    wire N__70640;
    wire N__70631;
    wire N__70626;
    wire N__70613;
    wire N__70610;
    wire N__70607;
    wire N__70604;
    wire N__70603;
    wire N__70600;
    wire N__70597;
    wire N__70594;
    wire N__70591;
    wire N__70586;
    wire N__70585;
    wire N__70582;
    wire N__70579;
    wire N__70576;
    wire N__70573;
    wire N__70570;
    wire N__70567;
    wire N__70564;
    wire N__70561;
    wire N__70556;
    wire N__70553;
    wire N__70552;
    wire N__70551;
    wire N__70550;
    wire N__70549;
    wire N__70548;
    wire N__70545;
    wire N__70544;
    wire N__70543;
    wire N__70542;
    wire N__70541;
    wire N__70540;
    wire N__70539;
    wire N__70536;
    wire N__70535;
    wire N__70528;
    wire N__70527;
    wire N__70526;
    wire N__70525;
    wire N__70524;
    wire N__70523;
    wire N__70522;
    wire N__70521;
    wire N__70518;
    wire N__70515;
    wire N__70514;
    wire N__70511;
    wire N__70500;
    wire N__70497;
    wire N__70494;
    wire N__70491;
    wire N__70478;
    wire N__70475;
    wire N__70472;
    wire N__70469;
    wire N__70468;
    wire N__70467;
    wire N__70466;
    wire N__70463;
    wire N__70462;
    wire N__70461;
    wire N__70460;
    wire N__70459;
    wire N__70458;
    wire N__70457;
    wire N__70456;
    wire N__70455;
    wire N__70452;
    wire N__70445;
    wire N__70442;
    wire N__70437;
    wire N__70432;
    wire N__70425;
    wire N__70422;
    wire N__70417;
    wire N__70404;
    wire N__70401;
    wire N__70398;
    wire N__70395;
    wire N__70390;
    wire N__70373;
    wire N__70370;
    wire N__70369;
    wire N__70366;
    wire N__70363;
    wire N__70360;
    wire N__70357;
    wire N__70354;
    wire N__70351;
    wire N__70348;
    wire N__70345;
    wire N__70340;
    wire N__70337;
    wire N__70334;
    wire N__70331;
    wire N__70330;
    wire N__70329;
    wire N__70328;
    wire N__70325;
    wire N__70322;
    wire N__70319;
    wire N__70318;
    wire N__70317;
    wire N__70314;
    wire N__70309;
    wire N__70306;
    wire N__70303;
    wire N__70300;
    wire N__70297;
    wire N__70292;
    wire N__70285;
    wire N__70282;
    wire N__70279;
    wire N__70276;
    wire N__70271;
    wire N__70268;
    wire N__70265;
    wire N__70262;
    wire N__70259;
    wire N__70256;
    wire N__70253;
    wire N__70250;
    wire N__70249;
    wire N__70246;
    wire N__70243;
    wire N__70240;
    wire N__70239;
    wire N__70236;
    wire N__70233;
    wire N__70230;
    wire N__70227;
    wire N__70224;
    wire N__70221;
    wire N__70218;
    wire N__70215;
    wire N__70212;
    wire N__70209;
    wire N__70206;
    wire N__70199;
    wire N__70198;
    wire N__70197;
    wire N__70192;
    wire N__70191;
    wire N__70188;
    wire N__70187;
    wire N__70186;
    wire N__70185;
    wire N__70184;
    wire N__70181;
    wire N__70178;
    wire N__70175;
    wire N__70172;
    wire N__70171;
    wire N__70170;
    wire N__70169;
    wire N__70168;
    wire N__70167;
    wire N__70160;
    wire N__70159;
    wire N__70158;
    wire N__70157;
    wire N__70154;
    wire N__70147;
    wire N__70140;
    wire N__70139;
    wire N__70134;
    wire N__70131;
    wire N__70128;
    wire N__70123;
    wire N__70118;
    wire N__70117;
    wire N__70114;
    wire N__70111;
    wire N__70106;
    wire N__70103;
    wire N__70100;
    wire N__70097;
    wire N__70096;
    wire N__70095;
    wire N__70094;
    wire N__70091;
    wire N__70090;
    wire N__70089;
    wire N__70088;
    wire N__70085;
    wire N__70080;
    wire N__70075;
    wire N__70072;
    wire N__70065;
    wire N__70062;
    wire N__70055;
    wire N__70054;
    wire N__70047;
    wire N__70042;
    wire N__70037;
    wire N__70034;
    wire N__70031;
    wire N__70028;
    wire N__70025;
    wire N__70016;
    wire N__70013;
    wire N__70012;
    wire N__70011;
    wire N__70008;
    wire N__70007;
    wire N__70004;
    wire N__70001;
    wire N__70000;
    wire N__69999;
    wire N__69998;
    wire N__69995;
    wire N__69992;
    wire N__69989;
    wire N__69988;
    wire N__69983;
    wire N__69978;
    wire N__69977;
    wire N__69974;
    wire N__69973;
    wire N__69972;
    wire N__69969;
    wire N__69968;
    wire N__69967;
    wire N__69966;
    wire N__69965;
    wire N__69962;
    wire N__69959;
    wire N__69954;
    wire N__69951;
    wire N__69948;
    wire N__69945;
    wire N__69944;
    wire N__69943;
    wire N__69940;
    wire N__69937;
    wire N__69932;
    wire N__69929;
    wire N__69928;
    wire N__69925;
    wire N__69922;
    wire N__69919;
    wire N__69914;
    wire N__69909;
    wire N__69908;
    wire N__69907;
    wire N__69904;
    wire N__69901;
    wire N__69898;
    wire N__69891;
    wire N__69886;
    wire N__69885;
    wire N__69882;
    wire N__69879;
    wire N__69876;
    wire N__69873;
    wire N__69868;
    wire N__69863;
    wire N__69860;
    wire N__69855;
    wire N__69852;
    wire N__69849;
    wire N__69846;
    wire N__69839;
    wire N__69836;
    wire N__69833;
    wire N__69830;
    wire N__69827;
    wire N__69822;
    wire N__69819;
    wire N__69812;
    wire N__69803;
    wire N__69800;
    wire N__69799;
    wire N__69798;
    wire N__69791;
    wire N__69790;
    wire N__69789;
    wire N__69786;
    wire N__69783;
    wire N__69780;
    wire N__69773;
    wire N__69770;
    wire N__69767;
    wire N__69766;
    wire N__69763;
    wire N__69760;
    wire N__69757;
    wire N__69752;
    wire N__69749;
    wire N__69748;
    wire N__69747;
    wire N__69746;
    wire N__69745;
    wire N__69744;
    wire N__69739;
    wire N__69736;
    wire N__69733;
    wire N__69730;
    wire N__69729;
    wire N__69726;
    wire N__69723;
    wire N__69720;
    wire N__69717;
    wire N__69716;
    wire N__69715;
    wire N__69712;
    wire N__69707;
    wire N__69700;
    wire N__69699;
    wire N__69698;
    wire N__69697;
    wire N__69694;
    wire N__69691;
    wire N__69690;
    wire N__69689;
    wire N__69684;
    wire N__69681;
    wire N__69680;
    wire N__69679;
    wire N__69678;
    wire N__69675;
    wire N__69672;
    wire N__69667;
    wire N__69666;
    wire N__69661;
    wire N__69658;
    wire N__69655;
    wire N__69652;
    wire N__69651;
    wire N__69648;
    wire N__69647;
    wire N__69646;
    wire N__69645;
    wire N__69642;
    wire N__69641;
    wire N__69640;
    wire N__69637;
    wire N__69634;
    wire N__69631;
    wire N__69628;
    wire N__69627;
    wire N__69624;
    wire N__69621;
    wire N__69618;
    wire N__69613;
    wire N__69610;
    wire N__69603;
    wire N__69596;
    wire N__69593;
    wire N__69590;
    wire N__69583;
    wire N__69580;
    wire N__69577;
    wire N__69574;
    wire N__69563;
    wire N__69560;
    wire N__69555;
    wire N__69552;
    wire N__69547;
    wire N__69544;
    wire N__69539;
    wire N__69530;
    wire N__69529;
    wire N__69526;
    wire N__69523;
    wire N__69520;
    wire N__69519;
    wire N__69514;
    wire N__69513;
    wire N__69512;
    wire N__69509;
    wire N__69506;
    wire N__69503;
    wire N__69500;
    wire N__69497;
    wire N__69496;
    wire N__69493;
    wire N__69490;
    wire N__69487;
    wire N__69484;
    wire N__69481;
    wire N__69478;
    wire N__69473;
    wire N__69470;
    wire N__69467;
    wire N__69458;
    wire N__69455;
    wire N__69454;
    wire N__69453;
    wire N__69452;
    wire N__69451;
    wire N__69450;
    wire N__69449;
    wire N__69446;
    wire N__69443;
    wire N__69440;
    wire N__69437;
    wire N__69434;
    wire N__69431;
    wire N__69428;
    wire N__69425;
    wire N__69422;
    wire N__69419;
    wire N__69416;
    wire N__69413;
    wire N__69408;
    wire N__69405;
    wire N__69402;
    wire N__69399;
    wire N__69396;
    wire N__69393;
    wire N__69390;
    wire N__69387;
    wire N__69382;
    wire N__69379;
    wire N__69376;
    wire N__69373;
    wire N__69370;
    wire N__69359;
    wire N__69356;
    wire N__69353;
    wire N__69350;
    wire N__69347;
    wire N__69344;
    wire N__69341;
    wire N__69338;
    wire N__69337;
    wire N__69334;
    wire N__69333;
    wire N__69332;
    wire N__69331;
    wire N__69324;
    wire N__69319;
    wire N__69318;
    wire N__69317;
    wire N__69312;
    wire N__69309;
    wire N__69306;
    wire N__69303;
    wire N__69298;
    wire N__69295;
    wire N__69292;
    wire N__69289;
    wire N__69284;
    wire N__69283;
    wire N__69282;
    wire N__69281;
    wire N__69276;
    wire N__69271;
    wire N__69270;
    wire N__69267;
    wire N__69264;
    wire N__69261;
    wire N__69258;
    wire N__69255;
    wire N__69248;
    wire N__69245;
    wire N__69244;
    wire N__69243;
    wire N__69240;
    wire N__69237;
    wire N__69234;
    wire N__69231;
    wire N__69228;
    wire N__69225;
    wire N__69222;
    wire N__69219;
    wire N__69216;
    wire N__69213;
    wire N__69210;
    wire N__69207;
    wire N__69204;
    wire N__69201;
    wire N__69198;
    wire N__69195;
    wire N__69188;
    wire N__69185;
    wire N__69182;
    wire N__69179;
    wire N__69176;
    wire N__69173;
    wire N__69170;
    wire N__69169;
    wire N__69168;
    wire N__69165;
    wire N__69162;
    wire N__69161;
    wire N__69160;
    wire N__69157;
    wire N__69156;
    wire N__69151;
    wire N__69150;
    wire N__69149;
    wire N__69146;
    wire N__69143;
    wire N__69140;
    wire N__69137;
    wire N__69134;
    wire N__69131;
    wire N__69128;
    wire N__69121;
    wire N__69118;
    wire N__69117;
    wire N__69112;
    wire N__69107;
    wire N__69106;
    wire N__69103;
    wire N__69100;
    wire N__69095;
    wire N__69092;
    wire N__69089;
    wire N__69084;
    wire N__69077;
    wire N__69074;
    wire N__69071;
    wire N__69070;
    wire N__69067;
    wire N__69064;
    wire N__69061;
    wire N__69058;
    wire N__69057;
    wire N__69054;
    wire N__69051;
    wire N__69048;
    wire N__69045;
    wire N__69042;
    wire N__69039;
    wire N__69036;
    wire N__69033;
    wire N__69030;
    wire N__69027;
    wire N__69024;
    wire N__69021;
    wire N__69014;
    wire N__69013;
    wire N__69012;
    wire N__69011;
    wire N__69010;
    wire N__69009;
    wire N__69006;
    wire N__69003;
    wire N__69002;
    wire N__68999;
    wire N__68996;
    wire N__68993;
    wire N__68990;
    wire N__68989;
    wire N__68986;
    wire N__68983;
    wire N__68980;
    wire N__68977;
    wire N__68970;
    wire N__68967;
    wire N__68962;
    wire N__68955;
    wire N__68950;
    wire N__68945;
    wire N__68944;
    wire N__68943;
    wire N__68942;
    wire N__68941;
    wire N__68940;
    wire N__68939;
    wire N__68936;
    wire N__68935;
    wire N__68934;
    wire N__68933;
    wire N__68932;
    wire N__68931;
    wire N__68930;
    wire N__68929;
    wire N__68928;
    wire N__68927;
    wire N__68926;
    wire N__68925;
    wire N__68924;
    wire N__68923;
    wire N__68922;
    wire N__68921;
    wire N__68920;
    wire N__68919;
    wire N__68918;
    wire N__68917;
    wire N__68914;
    wire N__68911;
    wire N__68910;
    wire N__68909;
    wire N__68908;
    wire N__68901;
    wire N__68898;
    wire N__68897;
    wire N__68896;
    wire N__68895;
    wire N__68894;
    wire N__68891;
    wire N__68886;
    wire N__68883;
    wire N__68880;
    wire N__68875;
    wire N__68872;
    wire N__68867;
    wire N__68860;
    wire N__68855;
    wire N__68852;
    wire N__68847;
    wire N__68846;
    wire N__68845;
    wire N__68844;
    wire N__68843;
    wire N__68842;
    wire N__68841;
    wire N__68836;
    wire N__68831;
    wire N__68826;
    wire N__68825;
    wire N__68824;
    wire N__68823;
    wire N__68822;
    wire N__68819;
    wire N__68816;
    wire N__68813;
    wire N__68812;
    wire N__68811;
    wire N__68810;
    wire N__68809;
    wire N__68804;
    wire N__68799;
    wire N__68796;
    wire N__68791;
    wire N__68790;
    wire N__68789;
    wire N__68786;
    wire N__68783;
    wire N__68774;
    wire N__68769;
    wire N__68762;
    wire N__68755;
    wire N__68752;
    wire N__68747;
    wire N__68746;
    wire N__68745;
    wire N__68744;
    wire N__68741;
    wire N__68734;
    wire N__68733;
    wire N__68730;
    wire N__68729;
    wire N__68728;
    wire N__68727;
    wire N__68722;
    wire N__68721;
    wire N__68720;
    wire N__68719;
    wire N__68712;
    wire N__68709;
    wire N__68706;
    wire N__68703;
    wire N__68698;
    wire N__68693;
    wire N__68690;
    wire N__68679;
    wire N__68674;
    wire N__68667;
    wire N__68662;
    wire N__68661;
    wire N__68660;
    wire N__68659;
    wire N__68658;
    wire N__68655;
    wire N__68652;
    wire N__68649;
    wire N__68646;
    wire N__68643;
    wire N__68640;
    wire N__68637;
    wire N__68632;
    wire N__68619;
    wire N__68614;
    wire N__68607;
    wire N__68600;
    wire N__68595;
    wire N__68588;
    wire N__68567;
    wire N__68566;
    wire N__68565;
    wire N__68560;
    wire N__68557;
    wire N__68556;
    wire N__68553;
    wire N__68550;
    wire N__68547;
    wire N__68544;
    wire N__68541;
    wire N__68538;
    wire N__68531;
    wire N__68530;
    wire N__68529;
    wire N__68528;
    wire N__68527;
    wire N__68526;
    wire N__68525;
    wire N__68524;
    wire N__68523;
    wire N__68522;
    wire N__68521;
    wire N__68518;
    wire N__68517;
    wire N__68516;
    wire N__68515;
    wire N__68512;
    wire N__68511;
    wire N__68510;
    wire N__68509;
    wire N__68508;
    wire N__68507;
    wire N__68506;
    wire N__68505;
    wire N__68502;
    wire N__68499;
    wire N__68494;
    wire N__68491;
    wire N__68490;
    wire N__68485;
    wire N__68484;
    wire N__68483;
    wire N__68482;
    wire N__68481;
    wire N__68480;
    wire N__68479;
    wire N__68472;
    wire N__68469;
    wire N__68468;
    wire N__68465;
    wire N__68464;
    wire N__68461;
    wire N__68460;
    wire N__68459;
    wire N__68458;
    wire N__68455;
    wire N__68452;
    wire N__68445;
    wire N__68442;
    wire N__68441;
    wire N__68440;
    wire N__68439;
    wire N__68438;
    wire N__68435;
    wire N__68432;
    wire N__68431;
    wire N__68426;
    wire N__68423;
    wire N__68420;
    wire N__68417;
    wire N__68414;
    wire N__68411;
    wire N__68404;
    wire N__68399;
    wire N__68396;
    wire N__68395;
    wire N__68394;
    wire N__68391;
    wire N__68388;
    wire N__68385;
    wire N__68382;
    wire N__68379;
    wire N__68378;
    wire N__68375;
    wire N__68374;
    wire N__68371;
    wire N__68368;
    wire N__68359;
    wire N__68352;
    wire N__68349;
    wire N__68346;
    wire N__68343;
    wire N__68340;
    wire N__68329;
    wire N__68322;
    wire N__68319;
    wire N__68316;
    wire N__68315;
    wire N__68312;
    wire N__68309;
    wire N__68306;
    wire N__68299;
    wire N__68292;
    wire N__68285;
    wire N__68282;
    wire N__68281;
    wire N__68280;
    wire N__68271;
    wire N__68270;
    wire N__68267;
    wire N__68260;
    wire N__68257;
    wire N__68256;
    wire N__68253;
    wire N__68240;
    wire N__68237;
    wire N__68234;
    wire N__68233;
    wire N__68232;
    wire N__68231;
    wire N__68230;
    wire N__68229;
    wire N__68228;
    wire N__68225;
    wire N__68222;
    wire N__68215;
    wire N__68212;
    wire N__68205;
    wire N__68196;
    wire N__68189;
    wire N__68174;
    wire N__68171;
    wire N__68168;
    wire N__68167;
    wire N__68166;
    wire N__68163;
    wire N__68158;
    wire N__68153;
    wire N__68150;
    wire N__68147;
    wire N__68144;
    wire N__68141;
    wire N__68140;
    wire N__68139;
    wire N__68138;
    wire N__68137;
    wire N__68136;
    wire N__68133;
    wire N__68130;
    wire N__68127;
    wire N__68124;
    wire N__68123;
    wire N__68122;
    wire N__68119;
    wire N__68116;
    wire N__68109;
    wire N__68106;
    wire N__68103;
    wire N__68100;
    wire N__68087;
    wire N__68086;
    wire N__68083;
    wire N__68080;
    wire N__68079;
    wire N__68078;
    wire N__68077;
    wire N__68076;
    wire N__68071;
    wire N__68068;
    wire N__68065;
    wire N__68062;
    wire N__68059;
    wire N__68058;
    wire N__68057;
    wire N__68054;
    wire N__68049;
    wire N__68046;
    wire N__68043;
    wire N__68040;
    wire N__68037;
    wire N__68034;
    wire N__68023;
    wire N__68020;
    wire N__68017;
    wire N__68012;
    wire N__68011;
    wire N__68008;
    wire N__68005;
    wire N__68004;
    wire N__68003;
    wire N__68002;
    wire N__68001;
    wire N__68000;
    wire N__67997;
    wire N__67994;
    wire N__67991;
    wire N__67988;
    wire N__67985;
    wire N__67982;
    wire N__67979;
    wire N__67964;
    wire N__67963;
    wire N__67960;
    wire N__67957;
    wire N__67952;
    wire N__67949;
    wire N__67946;
    wire N__67943;
    wire N__67942;
    wire N__67939;
    wire N__67938;
    wire N__67935;
    wire N__67932;
    wire N__67931;
    wire N__67928;
    wire N__67925;
    wire N__67922;
    wire N__67921;
    wire N__67918;
    wire N__67915;
    wire N__67912;
    wire N__67909;
    wire N__67906;
    wire N__67903;
    wire N__67900;
    wire N__67897;
    wire N__67894;
    wire N__67891;
    wire N__67888;
    wire N__67885;
    wire N__67880;
    wire N__67871;
    wire N__67868;
    wire N__67865;
    wire N__67864;
    wire N__67861;
    wire N__67860;
    wire N__67857;
    wire N__67854;
    wire N__67851;
    wire N__67848;
    wire N__67845;
    wire N__67842;
    wire N__67839;
    wire N__67836;
    wire N__67833;
    wire N__67830;
    wire N__67827;
    wire N__67820;
    wire N__67817;
    wire N__67814;
    wire N__67811;
    wire N__67808;
    wire N__67805;
    wire N__67802;
    wire N__67799;
    wire N__67796;
    wire N__67793;
    wire N__67790;
    wire N__67787;
    wire N__67784;
    wire N__67783;
    wire N__67780;
    wire N__67777;
    wire N__67774;
    wire N__67771;
    wire N__67766;
    wire N__67763;
    wire N__67760;
    wire N__67757;
    wire N__67756;
    wire N__67755;
    wire N__67754;
    wire N__67753;
    wire N__67750;
    wire N__67747;
    wire N__67744;
    wire N__67743;
    wire N__67742;
    wire N__67741;
    wire N__67738;
    wire N__67735;
    wire N__67732;
    wire N__67729;
    wire N__67726;
    wire N__67723;
    wire N__67720;
    wire N__67717;
    wire N__67712;
    wire N__67707;
    wire N__67704;
    wire N__67691;
    wire N__67688;
    wire N__67687;
    wire N__67686;
    wire N__67685;
    wire N__67682;
    wire N__67679;
    wire N__67676;
    wire N__67673;
    wire N__67672;
    wire N__67669;
    wire N__67668;
    wire N__67665;
    wire N__67662;
    wire N__67659;
    wire N__67656;
    wire N__67655;
    wire N__67654;
    wire N__67651;
    wire N__67648;
    wire N__67639;
    wire N__67636;
    wire N__67633;
    wire N__67622;
    wire N__67621;
    wire N__67618;
    wire N__67617;
    wire N__67614;
    wire N__67611;
    wire N__67610;
    wire N__67607;
    wire N__67604;
    wire N__67603;
    wire N__67602;
    wire N__67599;
    wire N__67596;
    wire N__67595;
    wire N__67590;
    wire N__67587;
    wire N__67584;
    wire N__67581;
    wire N__67578;
    wire N__67575;
    wire N__67570;
    wire N__67567;
    wire N__67556;
    wire N__67553;
    wire N__67550;
    wire N__67549;
    wire N__67546;
    wire N__67543;
    wire N__67538;
    wire N__67535;
    wire N__67532;
    wire N__67529;
    wire N__67526;
    wire N__67523;
    wire N__67520;
    wire N__67517;
    wire N__67516;
    wire N__67513;
    wire N__67512;
    wire N__67509;
    wire N__67508;
    wire N__67505;
    wire N__67504;
    wire N__67501;
    wire N__67498;
    wire N__67495;
    wire N__67494;
    wire N__67493;
    wire N__67490;
    wire N__67487;
    wire N__67484;
    wire N__67479;
    wire N__67476;
    wire N__67473;
    wire N__67460;
    wire N__67459;
    wire N__67456;
    wire N__67455;
    wire N__67452;
    wire N__67451;
    wire N__67450;
    wire N__67449;
    wire N__67446;
    wire N__67443;
    wire N__67442;
    wire N__67439;
    wire N__67436;
    wire N__67433;
    wire N__67432;
    wire N__67429;
    wire N__67424;
    wire N__67421;
    wire N__67414;
    wire N__67411;
    wire N__67400;
    wire N__67399;
    wire N__67396;
    wire N__67393;
    wire N__67392;
    wire N__67391;
    wire N__67390;
    wire N__67389;
    wire N__67388;
    wire N__67385;
    wire N__67382;
    wire N__67379;
    wire N__67376;
    wire N__67373;
    wire N__67370;
    wire N__67367;
    wire N__67352;
    wire N__67349;
    wire N__67348;
    wire N__67345;
    wire N__67342;
    wire N__67339;
    wire N__67336;
    wire N__67333;
    wire N__67330;
    wire N__67327;
    wire N__67324;
    wire N__67321;
    wire N__67316;
    wire N__67313;
    wire N__67312;
    wire N__67309;
    wire N__67306;
    wire N__67303;
    wire N__67300;
    wire N__67297;
    wire N__67294;
    wire N__67289;
    wire N__67286;
    wire N__67283;
    wire N__67282;
    wire N__67277;
    wire N__67274;
    wire N__67273;
    wire N__67272;
    wire N__67271;
    wire N__67270;
    wire N__67269;
    wire N__67268;
    wire N__67267;
    wire N__67266;
    wire N__67263;
    wire N__67256;
    wire N__67255;
    wire N__67254;
    wire N__67253;
    wire N__67252;
    wire N__67251;
    wire N__67250;
    wire N__67249;
    wire N__67248;
    wire N__67245;
    wire N__67244;
    wire N__67243;
    wire N__67242;
    wire N__67239;
    wire N__67236;
    wire N__67233;
    wire N__67232;
    wire N__67231;
    wire N__67230;
    wire N__67227;
    wire N__67226;
    wire N__67225;
    wire N__67220;
    wire N__67219;
    wire N__67218;
    wire N__67217;
    wire N__67216;
    wire N__67215;
    wire N__67214;
    wire N__67213;
    wire N__67212;
    wire N__67209;
    wire N__67208;
    wire N__67207;
    wire N__67206;
    wire N__67205;
    wire N__67204;
    wire N__67197;
    wire N__67184;
    wire N__67183;
    wire N__67180;
    wire N__67179;
    wire N__67176;
    wire N__67173;
    wire N__67170;
    wire N__67165;
    wire N__67164;
    wire N__67161;
    wire N__67158;
    wire N__67151;
    wire N__67148;
    wire N__67145;
    wire N__67138;
    wire N__67135;
    wire N__67130;
    wire N__67123;
    wire N__67116;
    wire N__67115;
    wire N__67112;
    wire N__67107;
    wire N__67100;
    wire N__67097;
    wire N__67090;
    wire N__67087;
    wire N__67066;
    wire N__67065;
    wire N__67064;
    wire N__67061;
    wire N__67060;
    wire N__67057;
    wire N__67054;
    wire N__67053;
    wire N__67052;
    wire N__67051;
    wire N__67048;
    wire N__67047;
    wire N__67046;
    wire N__67045;
    wire N__67044;
    wire N__67043;
    wire N__67042;
    wire N__67039;
    wire N__67036;
    wire N__67033;
    wire N__67030;
    wire N__67027;
    wire N__67020;
    wire N__67017;
    wire N__67014;
    wire N__67007;
    wire N__67004;
    wire N__66997;
    wire N__66994;
    wire N__66991;
    wire N__66988;
    wire N__66985;
    wire N__66982;
    wire N__66977;
    wire N__66976;
    wire N__66973;
    wire N__66970;
    wire N__66963;
    wire N__66958;
    wire N__66951;
    wire N__66948;
    wire N__66945;
    wire N__66942;
    wire N__66939;
    wire N__66930;
    wire N__66927;
    wire N__66920;
    wire N__66915;
    wire N__66910;
    wire N__66907;
    wire N__66902;
    wire N__66901;
    wire N__66898;
    wire N__66897;
    wire N__66896;
    wire N__66891;
    wire N__66888;
    wire N__66885;
    wire N__66882;
    wire N__66879;
    wire N__66876;
    wire N__66873;
    wire N__66870;
    wire N__66865;
    wire N__66860;
    wire N__66857;
    wire N__66856;
    wire N__66853;
    wire N__66850;
    wire N__66845;
    wire N__66844;
    wire N__66843;
    wire N__66840;
    wire N__66837;
    wire N__66834;
    wire N__66833;
    wire N__66832;
    wire N__66831;
    wire N__66828;
    wire N__66827;
    wire N__66822;
    wire N__66819;
    wire N__66816;
    wire N__66813;
    wire N__66810;
    wire N__66807;
    wire N__66806;
    wire N__66801;
    wire N__66796;
    wire N__66791;
    wire N__66788;
    wire N__66785;
    wire N__66778;
    wire N__66773;
    wire N__66772;
    wire N__66769;
    wire N__66768;
    wire N__66767;
    wire N__66766;
    wire N__66765;
    wire N__66764;
    wire N__66763;
    wire N__66762;
    wire N__66761;
    wire N__66758;
    wire N__66757;
    wire N__66756;
    wire N__66755;
    wire N__66754;
    wire N__66753;
    wire N__66750;
    wire N__66747;
    wire N__66746;
    wire N__66743;
    wire N__66742;
    wire N__66737;
    wire N__66736;
    wire N__66735;
    wire N__66734;
    wire N__66733;
    wire N__66730;
    wire N__66727;
    wire N__66722;
    wire N__66721;
    wire N__66720;
    wire N__66719;
    wire N__66718;
    wire N__66717;
    wire N__66716;
    wire N__66715;
    wire N__66714;
    wire N__66713;
    wire N__66710;
    wire N__66705;
    wire N__66704;
    wire N__66703;
    wire N__66702;
    wire N__66701;
    wire N__66700;
    wire N__66699;
    wire N__66698;
    wire N__66697;
    wire N__66696;
    wire N__66693;
    wire N__66690;
    wire N__66687;
    wire N__66686;
    wire N__66685;
    wire N__66684;
    wire N__66683;
    wire N__66682;
    wire N__66677;
    wire N__66672;
    wire N__66669;
    wire N__66666;
    wire N__66663;
    wire N__66662;
    wire N__66659;
    wire N__66654;
    wire N__66653;
    wire N__66652;
    wire N__66647;
    wire N__66644;
    wire N__66641;
    wire N__66634;
    wire N__66631;
    wire N__66630;
    wire N__66629;
    wire N__66626;
    wire N__66623;
    wire N__66618;
    wire N__66615;
    wire N__66612;
    wire N__66609;
    wire N__66604;
    wire N__66603;
    wire N__66602;
    wire N__66601;
    wire N__66600;
    wire N__66599;
    wire N__66598;
    wire N__66597;
    wire N__66596;
    wire N__66591;
    wire N__66586;
    wire N__66583;
    wire N__66582;
    wire N__66581;
    wire N__66580;
    wire N__66579;
    wire N__66578;
    wire N__66577;
    wire N__66574;
    wire N__66571;
    wire N__66570;
    wire N__66569;
    wire N__66564;
    wire N__66559;
    wire N__66552;
    wire N__66547;
    wire N__66540;
    wire N__66537;
    wire N__66532;
    wire N__66529;
    wire N__66526;
    wire N__66523;
    wire N__66516;
    wire N__66513;
    wire N__66508;
    wire N__66501;
    wire N__66492;
    wire N__66487;
    wire N__66482;
    wire N__66473;
    wire N__66468;
    wire N__66465;
    wire N__66462;
    wire N__66451;
    wire N__66448;
    wire N__66445;
    wire N__66442;
    wire N__66441;
    wire N__66438;
    wire N__66435;
    wire N__66426;
    wire N__66421;
    wire N__66418;
    wire N__66415;
    wire N__66410;
    wire N__66401;
    wire N__66394;
    wire N__66385;
    wire N__66378;
    wire N__66377;
    wire N__66376;
    wire N__66375;
    wire N__66372;
    wire N__66369;
    wire N__66362;
    wire N__66355;
    wire N__66350;
    wire N__66345;
    wire N__66340;
    wire N__66337;
    wire N__66320;
    wire N__66317;
    wire N__66316;
    wire N__66315;
    wire N__66314;
    wire N__66313;
    wire N__66312;
    wire N__66309;
    wire N__66304;
    wire N__66303;
    wire N__66300;
    wire N__66299;
    wire N__66298;
    wire N__66297;
    wire N__66296;
    wire N__66293;
    wire N__66292;
    wire N__66289;
    wire N__66288;
    wire N__66287;
    wire N__66284;
    wire N__66281;
    wire N__66278;
    wire N__66275;
    wire N__66272;
    wire N__66271;
    wire N__66270;
    wire N__66269;
    wire N__66266;
    wire N__66263;
    wire N__66260;
    wire N__66257;
    wire N__66254;
    wire N__66253;
    wire N__66252;
    wire N__66251;
    wire N__66250;
    wire N__66249;
    wire N__66248;
    wire N__66245;
    wire N__66242;
    wire N__66241;
    wire N__66240;
    wire N__66237;
    wire N__66230;
    wire N__66229;
    wire N__66228;
    wire N__66225;
    wire N__66222;
    wire N__66215;
    wire N__66208;
    wire N__66203;
    wire N__66198;
    wire N__66195;
    wire N__66188;
    wire N__66183;
    wire N__66180;
    wire N__66177;
    wire N__66176;
    wire N__66175;
    wire N__66174;
    wire N__66169;
    wire N__66164;
    wire N__66161;
    wire N__66154;
    wire N__66151;
    wire N__66140;
    wire N__66137;
    wire N__66134;
    wire N__66131;
    wire N__66128;
    wire N__66127;
    wire N__66124;
    wire N__66117;
    wire N__66112;
    wire N__66103;
    wire N__66100;
    wire N__66089;
    wire N__66086;
    wire N__66085;
    wire N__66084;
    wire N__66083;
    wire N__66082;
    wire N__66081;
    wire N__66080;
    wire N__66079;
    wire N__66078;
    wire N__66077;
    wire N__66076;
    wire N__66075;
    wire N__66074;
    wire N__66073;
    wire N__66068;
    wire N__66067;
    wire N__66066;
    wire N__66065;
    wire N__66064;
    wire N__66063;
    wire N__66062;
    wire N__66061;
    wire N__66060;
    wire N__66059;
    wire N__66058;
    wire N__66055;
    wire N__66052;
    wire N__66051;
    wire N__66050;
    wire N__66049;
    wire N__66048;
    wire N__66047;
    wire N__66046;
    wire N__66045;
    wire N__66040;
    wire N__66037;
    wire N__66030;
    wire N__66029;
    wire N__66028;
    wire N__66027;
    wire N__66026;
    wire N__66023;
    wire N__66020;
    wire N__66015;
    wire N__66014;
    wire N__66013;
    wire N__66012;
    wire N__66011;
    wire N__66010;
    wire N__66007;
    wire N__66000;
    wire N__65991;
    wire N__65990;
    wire N__65989;
    wire N__65986;
    wire N__65981;
    wire N__65978;
    wire N__65969;
    wire N__65968;
    wire N__65967;
    wire N__65966;
    wire N__65965;
    wire N__65964;
    wire N__65963;
    wire N__65962;
    wire N__65959;
    wire N__65958;
    wire N__65957;
    wire N__65956;
    wire N__65955;
    wire N__65954;
    wire N__65953;
    wire N__65952;
    wire N__65951;
    wire N__65944;
    wire N__65937;
    wire N__65936;
    wire N__65935;
    wire N__65932;
    wire N__65931;
    wire N__65930;
    wire N__65929;
    wire N__65928;
    wire N__65927;
    wire N__65926;
    wire N__65921;
    wire N__65918;
    wire N__65911;
    wire N__65906;
    wire N__65905;
    wire N__65904;
    wire N__65903;
    wire N__65902;
    wire N__65899;
    wire N__65896;
    wire N__65893;
    wire N__65890;
    wire N__65887;
    wire N__65884;
    wire N__65881;
    wire N__65878;
    wire N__65873;
    wire N__65868;
    wire N__65861;
    wire N__65852;
    wire N__65849;
    wire N__65840;
    wire N__65837;
    wire N__65834;
    wire N__65829;
    wire N__65828;
    wire N__65827;
    wire N__65826;
    wire N__65823;
    wire N__65820;
    wire N__65817;
    wire N__65814;
    wire N__65811;
    wire N__65808;
    wire N__65805;
    wire N__65802;
    wire N__65799;
    wire N__65794;
    wire N__65789;
    wire N__65784;
    wire N__65779;
    wire N__65774;
    wire N__65771;
    wire N__65766;
    wire N__65759;
    wire N__65756;
    wire N__65755;
    wire N__65754;
    wire N__65753;
    wire N__65750;
    wire N__65743;
    wire N__65740;
    wire N__65737;
    wire N__65734;
    wire N__65727;
    wire N__65724;
    wire N__65721;
    wire N__65720;
    wire N__65719;
    wire N__65718;
    wire N__65717;
    wire N__65716;
    wire N__65715;
    wire N__65712;
    wire N__65711;
    wire N__65710;
    wire N__65701;
    wire N__65698;
    wire N__65695;
    wire N__65690;
    wire N__65687;
    wire N__65676;
    wire N__65667;
    wire N__65660;
    wire N__65655;
    wire N__65652;
    wire N__65647;
    wire N__65642;
    wire N__65635;
    wire N__65628;
    wire N__65619;
    wire N__65610;
    wire N__65585;
    wire N__65584;
    wire N__65581;
    wire N__65576;
    wire N__65575;
    wire N__65574;
    wire N__65571;
    wire N__65570;
    wire N__65569;
    wire N__65566;
    wire N__65565;
    wire N__65564;
    wire N__65563;
    wire N__65562;
    wire N__65559;
    wire N__65558;
    wire N__65557;
    wire N__65556;
    wire N__65553;
    wire N__65552;
    wire N__65551;
    wire N__65550;
    wire N__65547;
    wire N__65546;
    wire N__65545;
    wire N__65544;
    wire N__65543;
    wire N__65542;
    wire N__65541;
    wire N__65540;
    wire N__65539;
    wire N__65538;
    wire N__65537;
    wire N__65536;
    wire N__65531;
    wire N__65528;
    wire N__65527;
    wire N__65526;
    wire N__65523;
    wire N__65522;
    wire N__65521;
    wire N__65520;
    wire N__65517;
    wire N__65514;
    wire N__65511;
    wire N__65508;
    wire N__65505;
    wire N__65502;
    wire N__65499;
    wire N__65494;
    wire N__65493;
    wire N__65490;
    wire N__65487;
    wire N__65484;
    wire N__65483;
    wire N__65482;
    wire N__65481;
    wire N__65480;
    wire N__65479;
    wire N__65474;
    wire N__65469;
    wire N__65464;
    wire N__65461;
    wire N__65458;
    wire N__65455;
    wire N__65452;
    wire N__65447;
    wire N__65446;
    wire N__65445;
    wire N__65444;
    wire N__65439;
    wire N__65434;
    wire N__65431;
    wire N__65428;
    wire N__65423;
    wire N__65418;
    wire N__65409;
    wire N__65408;
    wire N__65407;
    wire N__65404;
    wire N__65399;
    wire N__65386;
    wire N__65379;
    wire N__65374;
    wire N__65369;
    wire N__65366;
    wire N__65359;
    wire N__65352;
    wire N__65351;
    wire N__65348;
    wire N__65343;
    wire N__65340;
    wire N__65335;
    wire N__65326;
    wire N__65319;
    wire N__65316;
    wire N__65313;
    wire N__65310;
    wire N__65305;
    wire N__65298;
    wire N__65285;
    wire N__65282;
    wire N__65279;
    wire N__65276;
    wire N__65273;
    wire N__65272;
    wire N__65269;
    wire N__65266;
    wire N__65263;
    wire N__65260;
    wire N__65255;
    wire N__65252;
    wire N__65249;
    wire N__65246;
    wire N__65243;
    wire N__65240;
    wire N__65237;
    wire N__65236;
    wire N__65233;
    wire N__65228;
    wire N__65225;
    wire N__65222;
    wire N__65219;
    wire N__65216;
    wire N__65213;
    wire N__65210;
    wire N__65207;
    wire N__65204;
    wire N__65201;
    wire N__65198;
    wire N__65195;
    wire N__65192;
    wire N__65189;
    wire N__65186;
    wire N__65183;
    wire N__65180;
    wire N__65177;
    wire N__65174;
    wire N__65171;
    wire N__65168;
    wire N__65165;
    wire N__65162;
    wire N__65159;
    wire N__65156;
    wire N__65153;
    wire N__65150;
    wire N__65149;
    wire N__65146;
    wire N__65143;
    wire N__65140;
    wire N__65137;
    wire N__65134;
    wire N__65131;
    wire N__65126;
    wire N__65123;
    wire N__65120;
    wire N__65117;
    wire N__65114;
    wire N__65111;
    wire N__65108;
    wire N__65105;
    wire N__65102;
    wire N__65099;
    wire N__65096;
    wire N__65093;
    wire N__65090;
    wire N__65089;
    wire N__65086;
    wire N__65083;
    wire N__65078;
    wire N__65075;
    wire N__65072;
    wire N__65069;
    wire N__65066;
    wire N__65063;
    wire N__65060;
    wire N__65057;
    wire N__65056;
    wire N__65053;
    wire N__65050;
    wire N__65047;
    wire N__65044;
    wire N__65041;
    wire N__65038;
    wire N__65033;
    wire N__65030;
    wire N__65029;
    wire N__65026;
    wire N__65023;
    wire N__65020;
    wire N__65017;
    wire N__65014;
    wire N__65013;
    wire N__65010;
    wire N__65007;
    wire N__65004;
    wire N__65001;
    wire N__64998;
    wire N__64995;
    wire N__64992;
    wire N__64989;
    wire N__64984;
    wire N__64981;
    wire N__64976;
    wire N__64973;
    wire N__64970;
    wire N__64967;
    wire N__64966;
    wire N__64965;
    wire N__64964;
    wire N__64961;
    wire N__64958;
    wire N__64955;
    wire N__64952;
    wire N__64949;
    wire N__64946;
    wire N__64941;
    wire N__64940;
    wire N__64933;
    wire N__64930;
    wire N__64925;
    wire N__64922;
    wire N__64919;
    wire N__64916;
    wire N__64913;
    wire N__64910;
    wire N__64907;
    wire N__64904;
    wire N__64901;
    wire N__64900;
    wire N__64897;
    wire N__64894;
    wire N__64891;
    wire N__64888;
    wire N__64885;
    wire N__64882;
    wire N__64877;
    wire N__64876;
    wire N__64875;
    wire N__64872;
    wire N__64871;
    wire N__64870;
    wire N__64867;
    wire N__64864;
    wire N__64863;
    wire N__64862;
    wire N__64861;
    wire N__64858;
    wire N__64855;
    wire N__64852;
    wire N__64849;
    wire N__64844;
    wire N__64841;
    wire N__64838;
    wire N__64837;
    wire N__64834;
    wire N__64831;
    wire N__64828;
    wire N__64825;
    wire N__64822;
    wire N__64819;
    wire N__64814;
    wire N__64809;
    wire N__64804;
    wire N__64793;
    wire N__64790;
    wire N__64789;
    wire N__64786;
    wire N__64783;
    wire N__64778;
    wire N__64775;
    wire N__64772;
    wire N__64769;
    wire N__64766;
    wire N__64763;
    wire N__64760;
    wire N__64757;
    wire N__64754;
    wire N__64751;
    wire N__64748;
    wire N__64747;
    wire N__64742;
    wire N__64741;
    wire N__64740;
    wire N__64737;
    wire N__64734;
    wire N__64731;
    wire N__64728;
    wire N__64725;
    wire N__64722;
    wire N__64715;
    wire N__64712;
    wire N__64711;
    wire N__64710;
    wire N__64705;
    wire N__64702;
    wire N__64699;
    wire N__64698;
    wire N__64695;
    wire N__64694;
    wire N__64693;
    wire N__64692;
    wire N__64689;
    wire N__64686;
    wire N__64683;
    wire N__64680;
    wire N__64675;
    wire N__64664;
    wire N__64663;
    wire N__64662;
    wire N__64659;
    wire N__64656;
    wire N__64655;
    wire N__64652;
    wire N__64649;
    wire N__64646;
    wire N__64643;
    wire N__64642;
    wire N__64641;
    wire N__64638;
    wire N__64635;
    wire N__64632;
    wire N__64629;
    wire N__64626;
    wire N__64623;
    wire N__64620;
    wire N__64619;
    wire N__64616;
    wire N__64611;
    wire N__64608;
    wire N__64605;
    wire N__64602;
    wire N__64599;
    wire N__64598;
    wire N__64597;
    wire N__64596;
    wire N__64595;
    wire N__64594;
    wire N__64591;
    wire N__64588;
    wire N__64583;
    wire N__64580;
    wire N__64577;
    wire N__64574;
    wire N__64569;
    wire N__64566;
    wire N__64563;
    wire N__64544;
    wire N__64541;
    wire N__64538;
    wire N__64535;
    wire N__64532;
    wire N__64531;
    wire N__64528;
    wire N__64525;
    wire N__64524;
    wire N__64521;
    wire N__64518;
    wire N__64515;
    wire N__64512;
    wire N__64509;
    wire N__64506;
    wire N__64503;
    wire N__64500;
    wire N__64497;
    wire N__64492;
    wire N__64487;
    wire N__64486;
    wire N__64485;
    wire N__64482;
    wire N__64479;
    wire N__64476;
    wire N__64473;
    wire N__64470;
    wire N__64467;
    wire N__64466;
    wire N__64465;
    wire N__64462;
    wire N__64459;
    wire N__64456;
    wire N__64451;
    wire N__64442;
    wire N__64439;
    wire N__64436;
    wire N__64433;
    wire N__64430;
    wire N__64427;
    wire N__64424;
    wire N__64421;
    wire N__64418;
    wire N__64415;
    wire N__64412;
    wire N__64409;
    wire N__64406;
    wire N__64403;
    wire N__64400;
    wire N__64397;
    wire N__64396;
    wire N__64393;
    wire N__64390;
    wire N__64387;
    wire N__64382;
    wire N__64379;
    wire N__64376;
    wire N__64373;
    wire N__64370;
    wire N__64367;
    wire N__64364;
    wire N__64361;
    wire N__64358;
    wire N__64355;
    wire N__64352;
    wire N__64349;
    wire N__64346;
    wire N__64343;
    wire N__64340;
    wire N__64337;
    wire N__64334;
    wire N__64331;
    wire N__64328;
    wire N__64325;
    wire N__64324;
    wire N__64323;
    wire N__64320;
    wire N__64317;
    wire N__64314;
    wire N__64311;
    wire N__64308;
    wire N__64305;
    wire N__64298;
    wire N__64295;
    wire N__64292;
    wire N__64289;
    wire N__64286;
    wire N__64283;
    wire N__64280;
    wire N__64277;
    wire N__64274;
    wire N__64271;
    wire N__64268;
    wire N__64265;
    wire N__64262;
    wire N__64261;
    wire N__64258;
    wire N__64255;
    wire N__64254;
    wire N__64251;
    wire N__64250;
    wire N__64247;
    wire N__64246;
    wire N__64245;
    wire N__64242;
    wire N__64239;
    wire N__64236;
    wire N__64235;
    wire N__64232;
    wire N__64229;
    wire N__64226;
    wire N__64223;
    wire N__64218;
    wire N__64215;
    wire N__64202;
    wire N__64199;
    wire N__64196;
    wire N__64193;
    wire N__64190;
    wire N__64187;
    wire N__64184;
    wire N__64181;
    wire N__64178;
    wire N__64175;
    wire N__64172;
    wire N__64169;
    wire N__64166;
    wire N__64163;
    wire N__64160;
    wire N__64157;
    wire N__64154;
    wire N__64151;
    wire N__64148;
    wire N__64145;
    wire N__64142;
    wire N__64139;
    wire N__64136;
    wire N__64133;
    wire N__64130;
    wire N__64127;
    wire N__64124;
    wire N__64123;
    wire N__64120;
    wire N__64117;
    wire N__64112;
    wire N__64109;
    wire N__64108;
    wire N__64107;
    wire N__64106;
    wire N__64105;
    wire N__64102;
    wire N__64099;
    wire N__64092;
    wire N__64085;
    wire N__64084;
    wire N__64083;
    wire N__64080;
    wire N__64075;
    wire N__64070;
    wire N__64067;
    wire N__64064;
    wire N__64061;
    wire N__64058;
    wire N__64057;
    wire N__64054;
    wire N__64049;
    wire N__64046;
    wire N__64043;
    wire N__64040;
    wire N__64037;
    wire N__64034;
    wire N__64031;
    wire N__64028;
    wire N__64025;
    wire N__64022;
    wire N__64019;
    wire N__64018;
    wire N__64017;
    wire N__64014;
    wire N__64011;
    wire N__64008;
    wire N__64007;
    wire N__64004;
    wire N__64001;
    wire N__63998;
    wire N__63995;
    wire N__63992;
    wire N__63987;
    wire N__63984;
    wire N__63981;
    wire N__63978;
    wire N__63975;
    wire N__63968;
    wire N__63967;
    wire N__63964;
    wire N__63959;
    wire N__63956;
    wire N__63953;
    wire N__63950;
    wire N__63947;
    wire N__63944;
    wire N__63941;
    wire N__63938;
    wire N__63935;
    wire N__63932;
    wire N__63929;
    wire N__63926;
    wire N__63923;
    wire N__63920;
    wire N__63917;
    wire N__63914;
    wire N__63911;
    wire N__63908;
    wire N__63905;
    wire N__63902;
    wire N__63899;
    wire N__63896;
    wire N__63893;
    wire N__63890;
    wire N__63887;
    wire N__63884;
    wire N__63881;
    wire N__63878;
    wire N__63875;
    wire N__63872;
    wire N__63869;
    wire N__63866;
    wire N__63863;
    wire N__63860;
    wire N__63857;
    wire N__63854;
    wire N__63853;
    wire N__63852;
    wire N__63849;
    wire N__63848;
    wire N__63847;
    wire N__63844;
    wire N__63843;
    wire N__63842;
    wire N__63839;
    wire N__63836;
    wire N__63835;
    wire N__63832;
    wire N__63829;
    wire N__63826;
    wire N__63823;
    wire N__63820;
    wire N__63819;
    wire N__63816;
    wire N__63813;
    wire N__63810;
    wire N__63809;
    wire N__63806;
    wire N__63803;
    wire N__63802;
    wire N__63797;
    wire N__63794;
    wire N__63791;
    wire N__63788;
    wire N__63783;
    wire N__63780;
    wire N__63779;
    wire N__63778;
    wire N__63775;
    wire N__63774;
    wire N__63771;
    wire N__63768;
    wire N__63763;
    wire N__63760;
    wire N__63753;
    wire N__63748;
    wire N__63745;
    wire N__63742;
    wire N__63739;
    wire N__63734;
    wire N__63731;
    wire N__63728;
    wire N__63721;
    wire N__63716;
    wire N__63711;
    wire N__63706;
    wire N__63701;
    wire N__63700;
    wire N__63699;
    wire N__63694;
    wire N__63691;
    wire N__63688;
    wire N__63683;
    wire N__63680;
    wire N__63677;
    wire N__63674;
    wire N__63671;
    wire N__63670;
    wire N__63669;
    wire N__63668;
    wire N__63665;
    wire N__63662;
    wire N__63659;
    wire N__63658;
    wire N__63655;
    wire N__63652;
    wire N__63649;
    wire N__63646;
    wire N__63645;
    wire N__63644;
    wire N__63641;
    wire N__63640;
    wire N__63639;
    wire N__63638;
    wire N__63635;
    wire N__63628;
    wire N__63625;
    wire N__63622;
    wire N__63619;
    wire N__63616;
    wire N__63615;
    wire N__63614;
    wire N__63613;
    wire N__63612;
    wire N__63607;
    wire N__63598;
    wire N__63595;
    wire N__63594;
    wire N__63593;
    wire N__63592;
    wire N__63589;
    wire N__63586;
    wire N__63583;
    wire N__63582;
    wire N__63579;
    wire N__63576;
    wire N__63571;
    wire N__63568;
    wire N__63561;
    wire N__63558;
    wire N__63555;
    wire N__63548;
    wire N__63545;
    wire N__63542;
    wire N__63537;
    wire N__63524;
    wire N__63523;
    wire N__63520;
    wire N__63517;
    wire N__63516;
    wire N__63513;
    wire N__63512;
    wire N__63509;
    wire N__63506;
    wire N__63503;
    wire N__63500;
    wire N__63497;
    wire N__63488;
    wire N__63485;
    wire N__63482;
    wire N__63481;
    wire N__63478;
    wire N__63475;
    wire N__63472;
    wire N__63469;
    wire N__63464;
    wire N__63463;
    wire N__63462;
    wire N__63461;
    wire N__63460;
    wire N__63459;
    wire N__63456;
    wire N__63453;
    wire N__63448;
    wire N__63443;
    wire N__63442;
    wire N__63435;
    wire N__63432;
    wire N__63429;
    wire N__63426;
    wire N__63423;
    wire N__63418;
    wire N__63415;
    wire N__63414;
    wire N__63411;
    wire N__63408;
    wire N__63405;
    wire N__63402;
    wire N__63399;
    wire N__63392;
    wire N__63389;
    wire N__63386;
    wire N__63383;
    wire N__63380;
    wire N__63377;
    wire N__63374;
    wire N__63371;
    wire N__63370;
    wire N__63367;
    wire N__63364;
    wire N__63361;
    wire N__63360;
    wire N__63357;
    wire N__63354;
    wire N__63351;
    wire N__63348;
    wire N__63343;
    wire N__63340;
    wire N__63337;
    wire N__63334;
    wire N__63331;
    wire N__63328;
    wire N__63325;
    wire N__63320;
    wire N__63319;
    wire N__63314;
    wire N__63311;
    wire N__63308;
    wire N__63305;
    wire N__63302;
    wire N__63301;
    wire N__63300;
    wire N__63299;
    wire N__63298;
    wire N__63297;
    wire N__63294;
    wire N__63293;
    wire N__63292;
    wire N__63291;
    wire N__63290;
    wire N__63289;
    wire N__63280;
    wire N__63277;
    wire N__63276;
    wire N__63275;
    wire N__63274;
    wire N__63273;
    wire N__63270;
    wire N__63269;
    wire N__63266;
    wire N__63265;
    wire N__63262;
    wire N__63261;
    wire N__63260;
    wire N__63257;
    wire N__63256;
    wire N__63255;
    wire N__63254;
    wire N__63253;
    wire N__63250;
    wire N__63249;
    wire N__63248;
    wire N__63247;
    wire N__63246;
    wire N__63243;
    wire N__63242;
    wire N__63241;
    wire N__63240;
    wire N__63239;
    wire N__63238;
    wire N__63235;
    wire N__63232;
    wire N__63229;
    wire N__63226;
    wire N__63225;
    wire N__63222;
    wire N__63219;
    wire N__63218;
    wire N__63217;
    wire N__63214;
    wire N__63209;
    wire N__63204;
    wire N__63199;
    wire N__63196;
    wire N__63193;
    wire N__63188;
    wire N__63185;
    wire N__63178;
    wire N__63173;
    wire N__63170;
    wire N__63163;
    wire N__63158;
    wire N__63151;
    wire N__63150;
    wire N__63147;
    wire N__63142;
    wire N__63135;
    wire N__63132;
    wire N__63125;
    wire N__63122;
    wire N__63117;
    wire N__63116;
    wire N__63115;
    wire N__63114;
    wire N__63113;
    wire N__63112;
    wire N__63109;
    wire N__63106;
    wire N__63103;
    wire N__63100;
    wire N__63093;
    wire N__63090;
    wire N__63087;
    wire N__63082;
    wire N__63077;
    wire N__63076;
    wire N__63075;
    wire N__63070;
    wire N__63067;
    wire N__63062;
    wire N__63059;
    wire N__63056;
    wire N__63053;
    wire N__63050;
    wire N__63047;
    wire N__63044;
    wire N__63041;
    wire N__63036;
    wire N__63031;
    wire N__63030;
    wire N__63027;
    wire N__63026;
    wire N__63023;
    wire N__63022;
    wire N__63009;
    wire N__63004;
    wire N__63001;
    wire N__62998;
    wire N__62993;
    wire N__62986;
    wire N__62981;
    wire N__62978;
    wire N__62973;
    wire N__62968;
    wire N__62957;
    wire N__62956;
    wire N__62953;
    wire N__62950;
    wire N__62949;
    wire N__62946;
    wire N__62943;
    wire N__62940;
    wire N__62939;
    wire N__62936;
    wire N__62933;
    wire N__62928;
    wire N__62927;
    wire N__62922;
    wire N__62919;
    wire N__62916;
    wire N__62913;
    wire N__62910;
    wire N__62907;
    wire N__62904;
    wire N__62899;
    wire N__62894;
    wire N__62891;
    wire N__62890;
    wire N__62889;
    wire N__62888;
    wire N__62887;
    wire N__62886;
    wire N__62885;
    wire N__62884;
    wire N__62883;
    wire N__62882;
    wire N__62881;
    wire N__62878;
    wire N__62875;
    wire N__62874;
    wire N__62873;
    wire N__62872;
    wire N__62871;
    wire N__62868;
    wire N__62863;
    wire N__62860;
    wire N__62859;
    wire N__62856;
    wire N__62849;
    wire N__62846;
    wire N__62845;
    wire N__62842;
    wire N__62839;
    wire N__62836;
    wire N__62833;
    wire N__62830;
    wire N__62829;
    wire N__62826;
    wire N__62821;
    wire N__62820;
    wire N__62819;
    wire N__62818;
    wire N__62815;
    wire N__62812;
    wire N__62811;
    wire N__62806;
    wire N__62805;
    wire N__62802;
    wire N__62801;
    wire N__62798;
    wire N__62793;
    wire N__62786;
    wire N__62785;
    wire N__62782;
    wire N__62777;
    wire N__62774;
    wire N__62769;
    wire N__62766;
    wire N__62765;
    wire N__62764;
    wire N__62761;
    wire N__62758;
    wire N__62755;
    wire N__62752;
    wire N__62749;
    wire N__62746;
    wire N__62739;
    wire N__62736;
    wire N__62733;
    wire N__62726;
    wire N__62723;
    wire N__62718;
    wire N__62709;
    wire N__62704;
    wire N__62701;
    wire N__62698;
    wire N__62693;
    wire N__62688;
    wire N__62685;
    wire N__62672;
    wire N__62669;
    wire N__62666;
    wire N__62663;
    wire N__62660;
    wire N__62657;
    wire N__62656;
    wire N__62655;
    wire N__62652;
    wire N__62649;
    wire N__62648;
    wire N__62645;
    wire N__62642;
    wire N__62639;
    wire N__62636;
    wire N__62627;
    wire N__62624;
    wire N__62621;
    wire N__62618;
    wire N__62615;
    wire N__62612;
    wire N__62609;
    wire N__62608;
    wire N__62603;
    wire N__62600;
    wire N__62597;
    wire N__62594;
    wire N__62591;
    wire N__62588;
    wire N__62587;
    wire N__62586;
    wire N__62585;
    wire N__62584;
    wire N__62583;
    wire N__62580;
    wire N__62579;
    wire N__62576;
    wire N__62573;
    wire N__62572;
    wire N__62571;
    wire N__62570;
    wire N__62567;
    wire N__62564;
    wire N__62559;
    wire N__62558;
    wire N__62557;
    wire N__62556;
    wire N__62553;
    wire N__62552;
    wire N__62551;
    wire N__62550;
    wire N__62547;
    wire N__62544;
    wire N__62541;
    wire N__62538;
    wire N__62535;
    wire N__62530;
    wire N__62527;
    wire N__62524;
    wire N__62523;
    wire N__62520;
    wire N__62519;
    wire N__62518;
    wire N__62515;
    wire N__62512;
    wire N__62507;
    wire N__62506;
    wire N__62505;
    wire N__62504;
    wire N__62503;
    wire N__62502;
    wire N__62499;
    wire N__62496;
    wire N__62493;
    wire N__62490;
    wire N__62487;
    wire N__62482;
    wire N__62479;
    wire N__62476;
    wire N__62473;
    wire N__62468;
    wire N__62465;
    wire N__62462;
    wire N__62459;
    wire N__62456;
    wire N__62447;
    wire N__62444;
    wire N__62441;
    wire N__62436;
    wire N__62433;
    wire N__62430;
    wire N__62427;
    wire N__62422;
    wire N__62417;
    wire N__62414;
    wire N__62411;
    wire N__62402;
    wire N__62399;
    wire N__62392;
    wire N__62389;
    wire N__62382;
    wire N__62377;
    wire N__62366;
    wire N__62363;
    wire N__62360;
    wire N__62357;
    wire N__62354;
    wire N__62351;
    wire N__62348;
    wire N__62345;
    wire N__62342;
    wire N__62339;
    wire N__62338;
    wire N__62335;
    wire N__62332;
    wire N__62327;
    wire N__62324;
    wire N__62321;
    wire N__62320;
    wire N__62317;
    wire N__62316;
    wire N__62315;
    wire N__62314;
    wire N__62311;
    wire N__62308;
    wire N__62307;
    wire N__62306;
    wire N__62303;
    wire N__62302;
    wire N__62299;
    wire N__62298;
    wire N__62295;
    wire N__62292;
    wire N__62289;
    wire N__62286;
    wire N__62285;
    wire N__62282;
    wire N__62281;
    wire N__62278;
    wire N__62275;
    wire N__62274;
    wire N__62273;
    wire N__62272;
    wire N__62271;
    wire N__62270;
    wire N__62269;
    wire N__62266;
    wire N__62265;
    wire N__62262;
    wire N__62261;
    wire N__62256;
    wire N__62251;
    wire N__62244;
    wire N__62241;
    wire N__62238;
    wire N__62235;
    wire N__62234;
    wire N__62233;
    wire N__62232;
    wire N__62223;
    wire N__62220;
    wire N__62219;
    wire N__62216;
    wire N__62213;
    wire N__62210;
    wire N__62209;
    wire N__62206;
    wire N__62199;
    wire N__62192;
    wire N__62191;
    wire N__62190;
    wire N__62187;
    wire N__62186;
    wire N__62185;
    wire N__62182;
    wire N__62179;
    wire N__62176;
    wire N__62173;
    wire N__62170;
    wire N__62165;
    wire N__62162;
    wire N__62159;
    wire N__62158;
    wire N__62157;
    wire N__62156;
    wire N__62151;
    wire N__62148;
    wire N__62143;
    wire N__62138;
    wire N__62135;
    wire N__62132;
    wire N__62125;
    wire N__62122;
    wire N__62119;
    wire N__62114;
    wire N__62107;
    wire N__62100;
    wire N__62095;
    wire N__62090;
    wire N__62087;
    wire N__62084;
    wire N__62079;
    wire N__62076;
    wire N__62071;
    wire N__62060;
    wire N__62057;
    wire N__62054;
    wire N__62051;
    wire N__62048;
    wire N__62047;
    wire N__62044;
    wire N__62041;
    wire N__62038;
    wire N__62035;
    wire N__62030;
    wire N__62027;
    wire N__62026;
    wire N__62025;
    wire N__62024;
    wire N__62023;
    wire N__62022;
    wire N__62021;
    wire N__62018;
    wire N__62017;
    wire N__62014;
    wire N__62011;
    wire N__62010;
    wire N__62007;
    wire N__62004;
    wire N__62001;
    wire N__62000;
    wire N__61997;
    wire N__61994;
    wire N__61991;
    wire N__61984;
    wire N__61983;
    wire N__61982;
    wire N__61979;
    wire N__61978;
    wire N__61977;
    wire N__61976;
    wire N__61975;
    wire N__61972;
    wire N__61969;
    wire N__61966;
    wire N__61963;
    wire N__61960;
    wire N__61955;
    wire N__61952;
    wire N__61949;
    wire N__61948;
    wire N__61947;
    wire N__61944;
    wire N__61939;
    wire N__61936;
    wire N__61935;
    wire N__61932;
    wire N__61931;
    wire N__61930;
    wire N__61925;
    wire N__61922;
    wire N__61919;
    wire N__61914;
    wire N__61911;
    wire N__61908;
    wire N__61905;
    wire N__61902;
    wire N__61901;
    wire N__61896;
    wire N__61893;
    wire N__61890;
    wire N__61887;
    wire N__61882;
    wire N__61881;
    wire N__61878;
    wire N__61869;
    wire N__61866;
    wire N__61863;
    wire N__61860;
    wire N__61857;
    wire N__61852;
    wire N__61849;
    wire N__61846;
    wire N__61843;
    wire N__61840;
    wire N__61837;
    wire N__61836;
    wire N__61833;
    wire N__61830;
    wire N__61827;
    wire N__61820;
    wire N__61817;
    wire N__61812;
    wire N__61807;
    wire N__61804;
    wire N__61799;
    wire N__61794;
    wire N__61781;
    wire N__61778;
    wire N__61775;
    wire N__61772;
    wire N__61769;
    wire N__61766;
    wire N__61763;
    wire N__61760;
    wire N__61757;
    wire N__61754;
    wire N__61753;
    wire N__61750;
    wire N__61747;
    wire N__61742;
    wire N__61739;
    wire N__61736;
    wire N__61733;
    wire N__61730;
    wire N__61727;
    wire N__61724;
    wire N__61721;
    wire N__61718;
    wire N__61717;
    wire N__61716;
    wire N__61715;
    wire N__61714;
    wire N__61711;
    wire N__61710;
    wire N__61707;
    wire N__61704;
    wire N__61703;
    wire N__61702;
    wire N__61701;
    wire N__61698;
    wire N__61697;
    wire N__61692;
    wire N__61689;
    wire N__61686;
    wire N__61683;
    wire N__61682;
    wire N__61681;
    wire N__61676;
    wire N__61675;
    wire N__61672;
    wire N__61669;
    wire N__61668;
    wire N__61667;
    wire N__61666;
    wire N__61663;
    wire N__61662;
    wire N__61661;
    wire N__61658;
    wire N__61655;
    wire N__61650;
    wire N__61647;
    wire N__61644;
    wire N__61641;
    wire N__61640;
    wire N__61637;
    wire N__61636;
    wire N__61633;
    wire N__61630;
    wire N__61627;
    wire N__61624;
    wire N__61621;
    wire N__61618;
    wire N__61613;
    wire N__61610;
    wire N__61607;
    wire N__61604;
    wire N__61599;
    wire N__61596;
    wire N__61593;
    wire N__61588;
    wire N__61583;
    wire N__61580;
    wire N__61577;
    wire N__61574;
    wire N__61571;
    wire N__61568;
    wire N__61565;
    wire N__61562;
    wire N__61559;
    wire N__61556;
    wire N__61553;
    wire N__61546;
    wire N__61541;
    wire N__61536;
    wire N__61533;
    wire N__61526;
    wire N__61521;
    wire N__61516;
    wire N__61505;
    wire N__61502;
    wire N__61499;
    wire N__61496;
    wire N__61493;
    wire N__61492;
    wire N__61489;
    wire N__61486;
    wire N__61483;
    wire N__61478;
    wire N__61475;
    wire N__61474;
    wire N__61473;
    wire N__61472;
    wire N__61471;
    wire N__61470;
    wire N__61467;
    wire N__61466;
    wire N__61465;
    wire N__61464;
    wire N__61463;
    wire N__61462;
    wire N__61461;
    wire N__61460;
    wire N__61457;
    wire N__61454;
    wire N__61447;
    wire N__61446;
    wire N__61443;
    wire N__61440;
    wire N__61439;
    wire N__61436;
    wire N__61435;
    wire N__61434;
    wire N__61433;
    wire N__61428;
    wire N__61427;
    wire N__61426;
    wire N__61425;
    wire N__61422;
    wire N__61417;
    wire N__61410;
    wire N__61407;
    wire N__61404;
    wire N__61401;
    wire N__61398;
    wire N__61395;
    wire N__61390;
    wire N__61387;
    wire N__61384;
    wire N__61381;
    wire N__61378;
    wire N__61375;
    wire N__61372;
    wire N__61365;
    wire N__61364;
    wire N__61353;
    wire N__61350;
    wire N__61347;
    wire N__61344;
    wire N__61341;
    wire N__61334;
    wire N__61331;
    wire N__61328;
    wire N__61325;
    wire N__61322;
    wire N__61317;
    wire N__61314;
    wire N__61309;
    wire N__61298;
    wire N__61295;
    wire N__61292;
    wire N__61289;
    wire N__61286;
    wire N__61283;
    wire N__61280;
    wire N__61277;
    wire N__61276;
    wire N__61273;
    wire N__61270;
    wire N__61267;
    wire N__61264;
    wire N__61261;
    wire N__61258;
    wire N__61255;
    wire N__61252;
    wire N__61247;
    wire N__61244;
    wire N__61241;
    wire N__61238;
    wire N__61235;
    wire N__61232;
    wire N__61229;
    wire N__61226;
    wire N__61225;
    wire N__61224;
    wire N__61221;
    wire N__61218;
    wire N__61217;
    wire N__61216;
    wire N__61213;
    wire N__61212;
    wire N__61211;
    wire N__61210;
    wire N__61207;
    wire N__61204;
    wire N__61203;
    wire N__61200;
    wire N__61199;
    wire N__61196;
    wire N__61195;
    wire N__61194;
    wire N__61193;
    wire N__61190;
    wire N__61187;
    wire N__61184;
    wire N__61181;
    wire N__61176;
    wire N__61171;
    wire N__61170;
    wire N__61167;
    wire N__61164;
    wire N__61161;
    wire N__61158;
    wire N__61157;
    wire N__61156;
    wire N__61153;
    wire N__61152;
    wire N__61151;
    wire N__61148;
    wire N__61143;
    wire N__61140;
    wire N__61135;
    wire N__61132;
    wire N__61129;
    wire N__61126;
    wire N__61123;
    wire N__61120;
    wire N__61115;
    wire N__61112;
    wire N__61107;
    wire N__61104;
    wire N__61101;
    wire N__61094;
    wire N__61091;
    wire N__61082;
    wire N__61079;
    wire N__61076;
    wire N__61071;
    wire N__61068;
    wire N__61063;
    wire N__61058;
    wire N__61053;
    wire N__61050;
    wire N__61043;
    wire N__61042;
    wire N__61037;
    wire N__61034;
    wire N__61031;
    wire N__61028;
    wire N__61025;
    wire N__61022;
    wire N__61019;
    wire N__61018;
    wire N__61015;
    wire N__61014;
    wire N__61013;
    wire N__61012;
    wire N__61011;
    wire N__61010;
    wire N__61009;
    wire N__61008;
    wire N__61005;
    wire N__61002;
    wire N__60999;
    wire N__60996;
    wire N__60995;
    wire N__60994;
    wire N__60991;
    wire N__60990;
    wire N__60987;
    wire N__60984;
    wire N__60979;
    wire N__60972;
    wire N__60969;
    wire N__60966;
    wire N__60965;
    wire N__60964;
    wire N__60961;
    wire N__60958;
    wire N__60955;
    wire N__60954;
    wire N__60953;
    wire N__60950;
    wire N__60947;
    wire N__60944;
    wire N__60941;
    wire N__60940;
    wire N__60939;
    wire N__60938;
    wire N__60933;
    wire N__60928;
    wire N__60925;
    wire N__60920;
    wire N__60917;
    wire N__60914;
    wire N__60911;
    wire N__60906;
    wire N__60903;
    wire N__60896;
    wire N__60893;
    wire N__60890;
    wire N__60887;
    wire N__60884;
    wire N__60879;
    wire N__60870;
    wire N__60867;
    wire N__60864;
    wire N__60861;
    wire N__60858;
    wire N__60853;
    wire N__60848;
    wire N__60839;
    wire N__60836;
    wire N__60835;
    wire N__60832;
    wire N__60829;
    wire N__60826;
    wire N__60823;
    wire N__60818;
    wire N__60815;
    wire N__60814;
    wire N__60813;
    wire N__60812;
    wire N__60809;
    wire N__60806;
    wire N__60805;
    wire N__60802;
    wire N__60799;
    wire N__60796;
    wire N__60793;
    wire N__60790;
    wire N__60787;
    wire N__60784;
    wire N__60781;
    wire N__60780;
    wire N__60777;
    wire N__60774;
    wire N__60769;
    wire N__60766;
    wire N__60763;
    wire N__60760;
    wire N__60755;
    wire N__60752;
    wire N__60743;
    wire N__60740;
    wire N__60737;
    wire N__60736;
    wire N__60735;
    wire N__60734;
    wire N__60731;
    wire N__60730;
    wire N__60727;
    wire N__60724;
    wire N__60723;
    wire N__60720;
    wire N__60717;
    wire N__60714;
    wire N__60711;
    wire N__60708;
    wire N__60705;
    wire N__60702;
    wire N__60701;
    wire N__60696;
    wire N__60693;
    wire N__60686;
    wire N__60683;
    wire N__60682;
    wire N__60679;
    wire N__60676;
    wire N__60673;
    wire N__60668;
    wire N__60663;
    wire N__60660;
    wire N__60653;
    wire N__60650;
    wire N__60647;
    wire N__60644;
    wire N__60641;
    wire N__60638;
    wire N__60635;
    wire N__60632;
    wire N__60629;
    wire N__60628;
    wire N__60627;
    wire N__60626;
    wire N__60625;
    wire N__60624;
    wire N__60621;
    wire N__60618;
    wire N__60617;
    wire N__60616;
    wire N__60613;
    wire N__60610;
    wire N__60609;
    wire N__60606;
    wire N__60603;
    wire N__60602;
    wire N__60599;
    wire N__60598;
    wire N__60595;
    wire N__60594;
    wire N__60593;
    wire N__60590;
    wire N__60589;
    wire N__60586;
    wire N__60585;
    wire N__60580;
    wire N__60579;
    wire N__60576;
    wire N__60575;
    wire N__60574;
    wire N__60573;
    wire N__60572;
    wire N__60569;
    wire N__60568;
    wire N__60567;
    wire N__60566;
    wire N__60563;
    wire N__60560;
    wire N__60557;
    wire N__60554;
    wire N__60551;
    wire N__60546;
    wire N__60545;
    wire N__60544;
    wire N__60543;
    wire N__60542;
    wire N__60541;
    wire N__60540;
    wire N__60539;
    wire N__60536;
    wire N__60533;
    wire N__60530;
    wire N__60527;
    wire N__60524;
    wire N__60521;
    wire N__60518;
    wire N__60513;
    wire N__60508;
    wire N__60505;
    wire N__60500;
    wire N__60497;
    wire N__60492;
    wire N__60485;
    wire N__60482;
    wire N__60471;
    wire N__60466;
    wire N__60461;
    wire N__60454;
    wire N__60451;
    wire N__60448;
    wire N__60445;
    wire N__60438;
    wire N__60433;
    wire N__60430;
    wire N__60427;
    wire N__60418;
    wire N__60415;
    wire N__60412;
    wire N__60407;
    wire N__60402;
    wire N__60397;
    wire N__60386;
    wire N__60383;
    wire N__60380;
    wire N__60377;
    wire N__60374;
    wire N__60371;
    wire N__60368;
    wire N__60365;
    wire N__60362;
    wire N__60359;
    wire N__60358;
    wire N__60355;
    wire N__60352;
    wire N__60347;
    wire N__60344;
    wire N__60341;
    wire N__60338;
    wire N__60335;
    wire N__60332;
    wire N__60329;
    wire N__60326;
    wire N__60323;
    wire N__60320;
    wire N__60319;
    wire N__60316;
    wire N__60313;
    wire N__60308;
    wire N__60305;
    wire N__60302;
    wire N__60299;
    wire N__60296;
    wire N__60293;
    wire N__60290;
    wire N__60287;
    wire N__60284;
    wire N__60281;
    wire N__60280;
    wire N__60277;
    wire N__60274;
    wire N__60269;
    wire N__60266;
    wire N__60265;
    wire N__60264;
    wire N__60263;
    wire N__60262;
    wire N__60261;
    wire N__60260;
    wire N__60257;
    wire N__60254;
    wire N__60251;
    wire N__60248;
    wire N__60247;
    wire N__60246;
    wire N__60245;
    wire N__60242;
    wire N__60241;
    wire N__60238;
    wire N__60237;
    wire N__60236;
    wire N__60233;
    wire N__60228;
    wire N__60227;
    wire N__60224;
    wire N__60221;
    wire N__60220;
    wire N__60219;
    wire N__60218;
    wire N__60215;
    wire N__60214;
    wire N__60213;
    wire N__60210;
    wire N__60209;
    wire N__60208;
    wire N__60207;
    wire N__60206;
    wire N__60205;
    wire N__60202;
    wire N__60199;
    wire N__60198;
    wire N__60197;
    wire N__60196;
    wire N__60193;
    wire N__60192;
    wire N__60191;
    wire N__60190;
    wire N__60189;
    wire N__60188;
    wire N__60187;
    wire N__60184;
    wire N__60181;
    wire N__60178;
    wire N__60173;
    wire N__60170;
    wire N__60165;
    wire N__60162;
    wire N__60159;
    wire N__60158;
    wire N__60157;
    wire N__60152;
    wire N__60147;
    wire N__60144;
    wire N__60139;
    wire N__60134;
    wire N__60133;
    wire N__60130;
    wire N__60127;
    wire N__60124;
    wire N__60119;
    wire N__60118;
    wire N__60109;
    wire N__60102;
    wire N__60101;
    wire N__60100;
    wire N__60099;
    wire N__60096;
    wire N__60093;
    wire N__60090;
    wire N__60087;
    wire N__60084;
    wire N__60079;
    wire N__60074;
    wire N__60069;
    wire N__60066;
    wire N__60057;
    wire N__60052;
    wire N__60045;
    wire N__60042;
    wire N__60037;
    wire N__60030;
    wire N__60027;
    wire N__60024;
    wire N__60017;
    wire N__60010;
    wire N__60007;
    wire N__60004;
    wire N__59999;
    wire N__59992;
    wire N__59989;
    wire N__59986;
    wire N__59983;
    wire N__59980;
    wire N__59975;
    wire N__59970;
    wire N__59957;
    wire N__59954;
    wire N__59951;
    wire N__59948;
    wire N__59945;
    wire N__59942;
    wire N__59939;
    wire N__59936;
    wire N__59933;
    wire N__59930;
    wire N__59929;
    wire N__59926;
    wire N__59923;
    wire N__59920;
    wire N__59915;
    wire N__59912;
    wire N__59911;
    wire N__59910;
    wire N__59907;
    wire N__59904;
    wire N__59903;
    wire N__59902;
    wire N__59899;
    wire N__59898;
    wire N__59895;
    wire N__59894;
    wire N__59891;
    wire N__59888;
    wire N__59885;
    wire N__59884;
    wire N__59883;
    wire N__59882;
    wire N__59881;
    wire N__59878;
    wire N__59875;
    wire N__59874;
    wire N__59873;
    wire N__59870;
    wire N__59867;
    wire N__59866;
    wire N__59865;
    wire N__59864;
    wire N__59861;
    wire N__59858;
    wire N__59853;
    wire N__59850;
    wire N__59849;
    wire N__59846;
    wire N__59843;
    wire N__59842;
    wire N__59841;
    wire N__59840;
    wire N__59837;
    wire N__59834;
    wire N__59833;
    wire N__59830;
    wire N__59827;
    wire N__59824;
    wire N__59821;
    wire N__59818;
    wire N__59817;
    wire N__59814;
    wire N__59811;
    wire N__59806;
    wire N__59803;
    wire N__59802;
    wire N__59801;
    wire N__59800;
    wire N__59797;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59785;
    wire N__59780;
    wire N__59775;
    wire N__59772;
    wire N__59769;
    wire N__59766;
    wire N__59761;
    wire N__59756;
    wire N__59747;
    wire N__59742;
    wire N__59739;
    wire N__59732;
    wire N__59725;
    wire N__59718;
    wire N__59713;
    wire N__59708;
    wire N__59693;
    wire N__59690;
    wire N__59687;
    wire N__59684;
    wire N__59681;
    wire N__59678;
    wire N__59675;
    wire N__59672;
    wire N__59669;
    wire N__59666;
    wire N__59665;
    wire N__59662;
    wire N__59659;
    wire N__59656;
    wire N__59653;
    wire N__59648;
    wire N__59645;
    wire N__59644;
    wire N__59641;
    wire N__59640;
    wire N__59639;
    wire N__59638;
    wire N__59637;
    wire N__59634;
    wire N__59629;
    wire N__59626;
    wire N__59625;
    wire N__59624;
    wire N__59621;
    wire N__59620;
    wire N__59619;
    wire N__59618;
    wire N__59615;
    wire N__59612;
    wire N__59609;
    wire N__59606;
    wire N__59603;
    wire N__59602;
    wire N__59601;
    wire N__59600;
    wire N__59599;
    wire N__59596;
    wire N__59595;
    wire N__59592;
    wire N__59589;
    wire N__59588;
    wire N__59587;
    wire N__59586;
    wire N__59585;
    wire N__59584;
    wire N__59583;
    wire N__59582;
    wire N__59577;
    wire N__59574;
    wire N__59567;
    wire N__59564;
    wire N__59557;
    wire N__59554;
    wire N__59551;
    wire N__59550;
    wire N__59549;
    wire N__59546;
    wire N__59541;
    wire N__59540;
    wire N__59537;
    wire N__59534;
    wire N__59531;
    wire N__59528;
    wire N__59521;
    wire N__59518;
    wire N__59515;
    wire N__59512;
    wire N__59507;
    wire N__59504;
    wire N__59503;
    wire N__59500;
    wire N__59497;
    wire N__59494;
    wire N__59491;
    wire N__59488;
    wire N__59487;
    wire N__59486;
    wire N__59485;
    wire N__59484;
    wire N__59483;
    wire N__59480;
    wire N__59479;
    wire N__59478;
    wire N__59477;
    wire N__59476;
    wire N__59473;
    wire N__59470;
    wire N__59463;
    wire N__59454;
    wire N__59451;
    wire N__59448;
    wire N__59439;
    wire N__59436;
    wire N__59431;
    wire N__59424;
    wire N__59413;
    wire N__59406;
    wire N__59403;
    wire N__59384;
    wire N__59381;
    wire N__59378;
    wire N__59375;
    wire N__59372;
    wire N__59369;
    wire N__59366;
    wire N__59363;
    wire N__59360;
    wire N__59357;
    wire N__59354;
    wire N__59353;
    wire N__59350;
    wire N__59347;
    wire N__59342;
    wire N__59339;
    wire N__59338;
    wire N__59335;
    wire N__59332;
    wire N__59329;
    wire N__59328;
    wire N__59325;
    wire N__59322;
    wire N__59319;
    wire N__59316;
    wire N__59313;
    wire N__59306;
    wire N__59305;
    wire N__59302;
    wire N__59299;
    wire N__59298;
    wire N__59297;
    wire N__59296;
    wire N__59295;
    wire N__59292;
    wire N__59291;
    wire N__59290;
    wire N__59289;
    wire N__59288;
    wire N__59287;
    wire N__59286;
    wire N__59283;
    wire N__59282;
    wire N__59281;
    wire N__59276;
    wire N__59271;
    wire N__59268;
    wire N__59267;
    wire N__59266;
    wire N__59263;
    wire N__59262;
    wire N__59259;
    wire N__59250;
    wire N__59249;
    wire N__59248;
    wire N__59245;
    wire N__59240;
    wire N__59235;
    wire N__59232;
    wire N__59229;
    wire N__59226;
    wire N__59223;
    wire N__59220;
    wire N__59215;
    wire N__59212;
    wire N__59209;
    wire N__59202;
    wire N__59195;
    wire N__59188;
    wire N__59177;
    wire N__59176;
    wire N__59173;
    wire N__59170;
    wire N__59169;
    wire N__59166;
    wire N__59163;
    wire N__59160;
    wire N__59159;
    wire N__59158;
    wire N__59151;
    wire N__59146;
    wire N__59145;
    wire N__59144;
    wire N__59143;
    wire N__59142;
    wire N__59141;
    wire N__59140;
    wire N__59139;
    wire N__59138;
    wire N__59137;
    wire N__59136;
    wire N__59133;
    wire N__59130;
    wire N__59125;
    wire N__59124;
    wire N__59121;
    wire N__59120;
    wire N__59117;
    wire N__59114;
    wire N__59111;
    wire N__59108;
    wire N__59107;
    wire N__59106;
    wire N__59103;
    wire N__59102;
    wire N__59101;
    wire N__59100;
    wire N__59095;
    wire N__59088;
    wire N__59085;
    wire N__59082;
    wire N__59079;
    wire N__59076;
    wire N__59073;
    wire N__59070;
    wire N__59067;
    wire N__59066;
    wire N__59059;
    wire N__59056;
    wire N__59051;
    wire N__59050;
    wire N__59049;
    wire N__59048;
    wire N__59045;
    wire N__59044;
    wire N__59043;
    wire N__59042;
    wire N__59037;
    wire N__59034;
    wire N__59031;
    wire N__59024;
    wire N__59021;
    wire N__59018;
    wire N__59013;
    wire N__59010;
    wire N__59009;
    wire N__59006;
    wire N__59005;
    wire N__59002;
    wire N__59001;
    wire N__58998;
    wire N__58995;
    wire N__58988;
    wire N__58987;
    wire N__58984;
    wire N__58981;
    wire N__58976;
    wire N__58971;
    wire N__58968;
    wire N__58965;
    wire N__58958;
    wire N__58951;
    wire N__58946;
    wire N__58943;
    wire N__58940;
    wire N__58933;
    wire N__58930;
    wire N__58927;
    wire N__58920;
    wire N__58915;
    wire N__58910;
    wire N__58907;
    wire N__58904;
    wire N__58899;
    wire N__58894;
    wire N__58889;
    wire N__58888;
    wire N__58887;
    wire N__58886;
    wire N__58885;
    wire N__58884;
    wire N__58881;
    wire N__58878;
    wire N__58877;
    wire N__58874;
    wire N__58871;
    wire N__58868;
    wire N__58865;
    wire N__58864;
    wire N__58861;
    wire N__58858;
    wire N__58855;
    wire N__58850;
    wire N__58845;
    wire N__58842;
    wire N__58839;
    wire N__58836;
    wire N__58831;
    wire N__58828;
    wire N__58817;
    wire N__58816;
    wire N__58813;
    wire N__58812;
    wire N__58809;
    wire N__58808;
    wire N__58805;
    wire N__58802;
    wire N__58801;
    wire N__58800;
    wire N__58799;
    wire N__58796;
    wire N__58793;
    wire N__58790;
    wire N__58787;
    wire N__58784;
    wire N__58781;
    wire N__58778;
    wire N__58773;
    wire N__58768;
    wire N__58757;
    wire N__58756;
    wire N__58753;
    wire N__58752;
    wire N__58749;
    wire N__58746;
    wire N__58745;
    wire N__58742;
    wire N__58741;
    wire N__58740;
    wire N__58739;
    wire N__58736;
    wire N__58733;
    wire N__58730;
    wire N__58727;
    wire N__58724;
    wire N__58721;
    wire N__58718;
    wire N__58717;
    wire N__58714;
    wire N__58709;
    wire N__58706;
    wire N__58699;
    wire N__58696;
    wire N__58691;
    wire N__58684;
    wire N__58679;
    wire N__58678;
    wire N__58677;
    wire N__58676;
    wire N__58673;
    wire N__58670;
    wire N__58667;
    wire N__58666;
    wire N__58665;
    wire N__58664;
    wire N__58663;
    wire N__58660;
    wire N__58657;
    wire N__58654;
    wire N__58651;
    wire N__58648;
    wire N__58645;
    wire N__58642;
    wire N__58639;
    wire N__58636;
    wire N__58633;
    wire N__58630;
    wire N__58627;
    wire N__58610;
    wire N__58607;
    wire N__58606;
    wire N__58603;
    wire N__58602;
    wire N__58599;
    wire N__58596;
    wire N__58593;
    wire N__58590;
    wire N__58585;
    wire N__58582;
    wire N__58579;
    wire N__58576;
    wire N__58573;
    wire N__58570;
    wire N__58565;
    wire N__58564;
    wire N__58563;
    wire N__58562;
    wire N__58559;
    wire N__58556;
    wire N__58553;
    wire N__58552;
    wire N__58551;
    wire N__58548;
    wire N__58547;
    wire N__58544;
    wire N__58541;
    wire N__58538;
    wire N__58535;
    wire N__58534;
    wire N__58533;
    wire N__58530;
    wire N__58527;
    wire N__58526;
    wire N__58525;
    wire N__58524;
    wire N__58521;
    wire N__58516;
    wire N__58511;
    wire N__58510;
    wire N__58505;
    wire N__58502;
    wire N__58499;
    wire N__58498;
    wire N__58497;
    wire N__58496;
    wire N__58495;
    wire N__58494;
    wire N__58491;
    wire N__58488;
    wire N__58485;
    wire N__58482;
    wire N__58479;
    wire N__58476;
    wire N__58473;
    wire N__58470;
    wire N__58465;
    wire N__58462;
    wire N__58457;
    wire N__58456;
    wire N__58455;
    wire N__58452;
    wire N__58449;
    wire N__58444;
    wire N__58439;
    wire N__58434;
    wire N__58431;
    wire N__58428;
    wire N__58423;
    wire N__58420;
    wire N__58417;
    wire N__58414;
    wire N__58409;
    wire N__58406;
    wire N__58403;
    wire N__58396;
    wire N__58393;
    wire N__58390;
    wire N__58373;
    wire N__58372;
    wire N__58371;
    wire N__58370;
    wire N__58367;
    wire N__58366;
    wire N__58365;
    wire N__58362;
    wire N__58359;
    wire N__58356;
    wire N__58353;
    wire N__58350;
    wire N__58347;
    wire N__58344;
    wire N__58343;
    wire N__58340;
    wire N__58337;
    wire N__58330;
    wire N__58327;
    wire N__58324;
    wire N__58321;
    wire N__58318;
    wire N__58315;
    wire N__58312;
    wire N__58301;
    wire N__58300;
    wire N__58299;
    wire N__58296;
    wire N__58295;
    wire N__58294;
    wire N__58291;
    wire N__58288;
    wire N__58285;
    wire N__58284;
    wire N__58283;
    wire N__58280;
    wire N__58277;
    wire N__58274;
    wire N__58271;
    wire N__58268;
    wire N__58265;
    wire N__58262;
    wire N__58255;
    wire N__58250;
    wire N__58241;
    wire N__58238;
    wire N__58235;
    wire N__58234;
    wire N__58231;
    wire N__58228;
    wire N__58227;
    wire N__58222;
    wire N__58219;
    wire N__58216;
    wire N__58213;
    wire N__58210;
    wire N__58207;
    wire N__58202;
    wire N__58199;
    wire N__58196;
    wire N__58195;
    wire N__58194;
    wire N__58191;
    wire N__58190;
    wire N__58189;
    wire N__58188;
    wire N__58185;
    wire N__58184;
    wire N__58181;
    wire N__58178;
    wire N__58175;
    wire N__58172;
    wire N__58169;
    wire N__58166;
    wire N__58165;
    wire N__58162;
    wire N__58159;
    wire N__58150;
    wire N__58147;
    wire N__58144;
    wire N__58139;
    wire N__58134;
    wire N__58127;
    wire N__58126;
    wire N__58123;
    wire N__58120;
    wire N__58119;
    wire N__58118;
    wire N__58115;
    wire N__58112;
    wire N__58111;
    wire N__58110;
    wire N__58109;
    wire N__58108;
    wire N__58105;
    wire N__58102;
    wire N__58099;
    wire N__58096;
    wire N__58093;
    wire N__58090;
    wire N__58087;
    wire N__58084;
    wire N__58081;
    wire N__58076;
    wire N__58073;
    wire N__58058;
    wire N__58057;
    wire N__58056;
    wire N__58053;
    wire N__58052;
    wire N__58051;
    wire N__58050;
    wire N__58049;
    wire N__58046;
    wire N__58043;
    wire N__58040;
    wire N__58037;
    wire N__58034;
    wire N__58031;
    wire N__58028;
    wire N__58025;
    wire N__58022;
    wire N__58019;
    wire N__58004;
    wire N__58001;
    wire N__57998;
    wire N__57997;
    wire N__57994;
    wire N__57991;
    wire N__57988;
    wire N__57985;
    wire N__57982;
    wire N__57981;
    wire N__57978;
    wire N__57975;
    wire N__57972;
    wire N__57969;
    wire N__57964;
    wire N__57961;
    wire N__57958;
    wire N__57955;
    wire N__57950;
    wire N__57947;
    wire N__57946;
    wire N__57943;
    wire N__57940;
    wire N__57935;
    wire N__57934;
    wire N__57931;
    wire N__57928;
    wire N__57925;
    wire N__57922;
    wire N__57917;
    wire N__57914;
    wire N__57911;
    wire N__57908;
    wire N__57905;
    wire N__57902;
    wire N__57899;
    wire N__57896;
    wire N__57893;
    wire N__57892;
    wire N__57891;
    wire N__57888;
    wire N__57885;
    wire N__57882;
    wire N__57877;
    wire N__57872;
    wire N__57869;
    wire N__57866;
    wire N__57863;
    wire N__57860;
    wire N__57859;
    wire N__57856;
    wire N__57853;
    wire N__57852;
    wire N__57849;
    wire N__57846;
    wire N__57843;
    wire N__57840;
    wire N__57835;
    wire N__57830;
    wire N__57827;
    wire N__57824;
    wire N__57821;
    wire N__57820;
    wire N__57819;
    wire N__57816;
    wire N__57813;
    wire N__57810;
    wire N__57809;
    wire N__57808;
    wire N__57805;
    wire N__57802;
    wire N__57801;
    wire N__57798;
    wire N__57793;
    wire N__57792;
    wire N__57791;
    wire N__57788;
    wire N__57785;
    wire N__57782;
    wire N__57777;
    wire N__57774;
    wire N__57771;
    wire N__57768;
    wire N__57765;
    wire N__57762;
    wire N__57761;
    wire N__57758;
    wire N__57755;
    wire N__57752;
    wire N__57751;
    wire N__57748;
    wire N__57743;
    wire N__57740;
    wire N__57737;
    wire N__57732;
    wire N__57729;
    wire N__57728;
    wire N__57725;
    wire N__57722;
    wire N__57715;
    wire N__57712;
    wire N__57709;
    wire N__57706;
    wire N__57703;
    wire N__57700;
    wire N__57697;
    wire N__57686;
    wire N__57685;
    wire N__57682;
    wire N__57679;
    wire N__57676;
    wire N__57675;
    wire N__57672;
    wire N__57669;
    wire N__57666;
    wire N__57661;
    wire N__57658;
    wire N__57655;
    wire N__57652;
    wire N__57649;
    wire N__57646;
    wire N__57643;
    wire N__57638;
    wire N__57635;
    wire N__57632;
    wire N__57631;
    wire N__57628;
    wire N__57625;
    wire N__57622;
    wire N__57621;
    wire N__57616;
    wire N__57613;
    wire N__57610;
    wire N__57607;
    wire N__57604;
    wire N__57601;
    wire N__57598;
    wire N__57593;
    wire N__57590;
    wire N__57587;
    wire N__57586;
    wire N__57583;
    wire N__57582;
    wire N__57579;
    wire N__57576;
    wire N__57573;
    wire N__57570;
    wire N__57567;
    wire N__57564;
    wire N__57561;
    wire N__57558;
    wire N__57555;
    wire N__57552;
    wire N__57549;
    wire N__57546;
    wire N__57543;
    wire N__57540;
    wire N__57537;
    wire N__57534;
    wire N__57527;
    wire N__57524;
    wire N__57523;
    wire N__57518;
    wire N__57515;
    wire N__57514;
    wire N__57511;
    wire N__57508;
    wire N__57503;
    wire N__57500;
    wire N__57497;
    wire N__57494;
    wire N__57491;
    wire N__57488;
    wire N__57485;
    wire N__57482;
    wire N__57479;
    wire N__57476;
    wire N__57473;
    wire N__57470;
    wire N__57467;
    wire N__57464;
    wire N__57461;
    wire N__57458;
    wire N__57455;
    wire N__57454;
    wire N__57451;
    wire N__57448;
    wire N__57445;
    wire N__57442;
    wire N__57439;
    wire N__57436;
    wire N__57433;
    wire N__57430;
    wire N__57427;
    wire N__57422;
    wire N__57421;
    wire N__57420;
    wire N__57419;
    wire N__57416;
    wire N__57413;
    wire N__57412;
    wire N__57407;
    wire N__57406;
    wire N__57405;
    wire N__57400;
    wire N__57397;
    wire N__57396;
    wire N__57393;
    wire N__57390;
    wire N__57389;
    wire N__57388;
    wire N__57385;
    wire N__57384;
    wire N__57383;
    wire N__57382;
    wire N__57379;
    wire N__57378;
    wire N__57373;
    wire N__57372;
    wire N__57371;
    wire N__57368;
    wire N__57365;
    wire N__57360;
    wire N__57355;
    wire N__57352;
    wire N__57351;
    wire N__57350;
    wire N__57349;
    wire N__57346;
    wire N__57343;
    wire N__57340;
    wire N__57337;
    wire N__57332;
    wire N__57329;
    wire N__57322;
    wire N__57321;
    wire N__57316;
    wire N__57311;
    wire N__57300;
    wire N__57295;
    wire N__57292;
    wire N__57285;
    wire N__57282;
    wire N__57279;
    wire N__57276;
    wire N__57273;
    wire N__57270;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57258;
    wire N__57255;
    wire N__57248;
    wire N__57245;
    wire N__57242;
    wire N__57239;
    wire N__57238;
    wire N__57235;
    wire N__57232;
    wire N__57231;
    wire N__57228;
    wire N__57227;
    wire N__57224;
    wire N__57221;
    wire N__57218;
    wire N__57215;
    wire N__57212;
    wire N__57209;
    wire N__57204;
    wire N__57199;
    wire N__57196;
    wire N__57193;
    wire N__57190;
    wire N__57185;
    wire N__57182;
    wire N__57179;
    wire N__57176;
    wire N__57173;
    wire N__57170;
    wire N__57167;
    wire N__57166;
    wire N__57163;
    wire N__57160;
    wire N__57157;
    wire N__57154;
    wire N__57151;
    wire N__57148;
    wire N__57145;
    wire N__57142;
    wire N__57137;
    wire N__57134;
    wire N__57131;
    wire N__57128;
    wire N__57125;
    wire N__57122;
    wire N__57121;
    wire N__57118;
    wire N__57113;
    wire N__57110;
    wire N__57109;
    wire N__57104;
    wire N__57101;
    wire N__57098;
    wire N__57095;
    wire N__57094;
    wire N__57091;
    wire N__57088;
    wire N__57085;
    wire N__57082;
    wire N__57077;
    wire N__57074;
    wire N__57073;
    wire N__57068;
    wire N__57065;
    wire N__57062;
    wire N__57059;
    wire N__57056;
    wire N__57053;
    wire N__57050;
    wire N__57047;
    wire N__57046;
    wire N__57043;
    wire N__57040;
    wire N__57039;
    wire N__57034;
    wire N__57033;
    wire N__57032;
    wire N__57031;
    wire N__57030;
    wire N__57029;
    wire N__57028;
    wire N__57025;
    wire N__57024;
    wire N__57021;
    wire N__57016;
    wire N__57015;
    wire N__57012;
    wire N__57009;
    wire N__57006;
    wire N__57003;
    wire N__57000;
    wire N__56997;
    wire N__56994;
    wire N__56991;
    wire N__56988;
    wire N__56987;
    wire N__56984;
    wire N__56977;
    wire N__56974;
    wire N__56971;
    wire N__56966;
    wire N__56963;
    wire N__56960;
    wire N__56955;
    wire N__56942;
    wire N__56939;
    wire N__56936;
    wire N__56933;
    wire N__56930;
    wire N__56929;
    wire N__56928;
    wire N__56925;
    wire N__56920;
    wire N__56917;
    wire N__56914;
    wire N__56911;
    wire N__56910;
    wire N__56909;
    wire N__56906;
    wire N__56905;
    wire N__56904;
    wire N__56901;
    wire N__56900;
    wire N__56895;
    wire N__56892;
    wire N__56889;
    wire N__56886;
    wire N__56883;
    wire N__56880;
    wire N__56877;
    wire N__56870;
    wire N__56865;
    wire N__56862;
    wire N__56859;
    wire N__56852;
    wire N__56849;
    wire N__56846;
    wire N__56843;
    wire N__56840;
    wire N__56839;
    wire N__56836;
    wire N__56833;
    wire N__56830;
    wire N__56829;
    wire N__56828;
    wire N__56825;
    wire N__56824;
    wire N__56823;
    wire N__56820;
    wire N__56815;
    wire N__56812;
    wire N__56809;
    wire N__56806;
    wire N__56805;
    wire N__56804;
    wire N__56799;
    wire N__56796;
    wire N__56793;
    wire N__56788;
    wire N__56787;
    wire N__56784;
    wire N__56781;
    wire N__56778;
    wire N__56773;
    wire N__56768;
    wire N__56759;
    wire N__56756;
    wire N__56753;
    wire N__56750;
    wire N__56749;
    wire N__56748;
    wire N__56745;
    wire N__56742;
    wire N__56741;
    wire N__56738;
    wire N__56737;
    wire N__56734;
    wire N__56731;
    wire N__56728;
    wire N__56723;
    wire N__56720;
    wire N__56719;
    wire N__56718;
    wire N__56713;
    wire N__56710;
    wire N__56707;
    wire N__56702;
    wire N__56699;
    wire N__56696;
    wire N__56693;
    wire N__56688;
    wire N__56685;
    wire N__56678;
    wire N__56675;
    wire N__56672;
    wire N__56669;
    wire N__56666;
    wire N__56663;
    wire N__56660;
    wire N__56657;
    wire N__56656;
    wire N__56651;
    wire N__56648;
    wire N__56647;
    wire N__56644;
    wire N__56641;
    wire N__56638;
    wire N__56635;
    wire N__56632;
    wire N__56627;
    wire N__56624;
    wire N__56623;
    wire N__56622;
    wire N__56621;
    wire N__56618;
    wire N__56615;
    wire N__56610;
    wire N__56607;
    wire N__56604;
    wire N__56603;
    wire N__56600;
    wire N__56595;
    wire N__56592;
    wire N__56589;
    wire N__56586;
    wire N__56583;
    wire N__56580;
    wire N__56577;
    wire N__56574;
    wire N__56573;
    wire N__56570;
    wire N__56567;
    wire N__56564;
    wire N__56561;
    wire N__56558;
    wire N__56555;
    wire N__56552;
    wire N__56543;
    wire N__56542;
    wire N__56539;
    wire N__56536;
    wire N__56533;
    wire N__56532;
    wire N__56529;
    wire N__56526;
    wire N__56523;
    wire N__56520;
    wire N__56517;
    wire N__56514;
    wire N__56511;
    wire N__56506;
    wire N__56503;
    wire N__56500;
    wire N__56495;
    wire N__56492;
    wire N__56491;
    wire N__56490;
    wire N__56487;
    wire N__56482;
    wire N__56479;
    wire N__56474;
    wire N__56473;
    wire N__56472;
    wire N__56469;
    wire N__56466;
    wire N__56465;
    wire N__56462;
    wire N__56459;
    wire N__56456;
    wire N__56453;
    wire N__56450;
    wire N__56445;
    wire N__56442;
    wire N__56439;
    wire N__56434;
    wire N__56431;
    wire N__56426;
    wire N__56423;
    wire N__56420;
    wire N__56417;
    wire N__56416;
    wire N__56415;
    wire N__56414;
    wire N__56413;
    wire N__56410;
    wire N__56407;
    wire N__56402;
    wire N__56401;
    wire N__56398;
    wire N__56395;
    wire N__56394;
    wire N__56391;
    wire N__56388;
    wire N__56385;
    wire N__56382;
    wire N__56379;
    wire N__56378;
    wire N__56377;
    wire N__56374;
    wire N__56371;
    wire N__56366;
    wire N__56361;
    wire N__56360;
    wire N__56359;
    wire N__56358;
    wire N__56357;
    wire N__56352;
    wire N__56347;
    wire N__56346;
    wire N__56345;
    wire N__56342;
    wire N__56339;
    wire N__56336;
    wire N__56329;
    wire N__56328;
    wire N__56327;
    wire N__56326;
    wire N__56321;
    wire N__56316;
    wire N__56313;
    wire N__56306;
    wire N__56303;
    wire N__56298;
    wire N__56285;
    wire N__56282;
    wire N__56279;
    wire N__56276;
    wire N__56273;
    wire N__56272;
    wire N__56269;
    wire N__56268;
    wire N__56267;
    wire N__56266;
    wire N__56263;
    wire N__56260;
    wire N__56259;
    wire N__56256;
    wire N__56253;
    wire N__56250;
    wire N__56247;
    wire N__56244;
    wire N__56241;
    wire N__56240;
    wire N__56239;
    wire N__56236;
    wire N__56233;
    wire N__56230;
    wire N__56229;
    wire N__56228;
    wire N__56225;
    wire N__56224;
    wire N__56223;
    wire N__56218;
    wire N__56213;
    wire N__56206;
    wire N__56203;
    wire N__56202;
    wire N__56201;
    wire N__56200;
    wire N__56197;
    wire N__56196;
    wire N__56193;
    wire N__56188;
    wire N__56185;
    wire N__56182;
    wire N__56179;
    wire N__56168;
    wire N__56165;
    wire N__56150;
    wire N__56147;
    wire N__56144;
    wire N__56141;
    wire N__56138;
    wire N__56135;
    wire N__56132;
    wire N__56131;
    wire N__56130;
    wire N__56127;
    wire N__56124;
    wire N__56121;
    wire N__56120;
    wire N__56117;
    wire N__56116;
    wire N__56115;
    wire N__56112;
    wire N__56109;
    wire N__56106;
    wire N__56103;
    wire N__56100;
    wire N__56097;
    wire N__56096;
    wire N__56093;
    wire N__56090;
    wire N__56087;
    wire N__56086;
    wire N__56083;
    wire N__56082;
    wire N__56079;
    wire N__56078;
    wire N__56077;
    wire N__56076;
    wire N__56073;
    wire N__56070;
    wire N__56069;
    wire N__56068;
    wire N__56065;
    wire N__56060;
    wire N__56057;
    wire N__56054;
    wire N__56051;
    wire N__56048;
    wire N__56043;
    wire N__56040;
    wire N__56037;
    wire N__56032;
    wire N__56029;
    wire N__56022;
    wire N__56003;
    wire N__56000;
    wire N__55997;
    wire N__55994;
    wire N__55993;
    wire N__55992;
    wire N__55991;
    wire N__55990;
    wire N__55989;
    wire N__55986;
    wire N__55985;
    wire N__55984;
    wire N__55979;
    wire N__55976;
    wire N__55973;
    wire N__55970;
    wire N__55967;
    wire N__55964;
    wire N__55961;
    wire N__55960;
    wire N__55959;
    wire N__55958;
    wire N__55957;
    wire N__55954;
    wire N__55953;
    wire N__55950;
    wire N__55949;
    wire N__55946;
    wire N__55941;
    wire N__55938;
    wire N__55931;
    wire N__55928;
    wire N__55925;
    wire N__55922;
    wire N__55919;
    wire N__55916;
    wire N__55913;
    wire N__55904;
    wire N__55901;
    wire N__55898;
    wire N__55893;
    wire N__55888;
    wire N__55887;
    wire N__55886;
    wire N__55885;
    wire N__55882;
    wire N__55879;
    wire N__55876;
    wire N__55875;
    wire N__55872;
    wire N__55869;
    wire N__55862;
    wire N__55859;
    wire N__55854;
    wire N__55851;
    wire N__55848;
    wire N__55835;
    wire N__55832;
    wire N__55829;
    wire N__55826;
    wire N__55823;
    wire N__55822;
    wire N__55821;
    wire N__55818;
    wire N__55817;
    wire N__55816;
    wire N__55813;
    wire N__55812;
    wire N__55811;
    wire N__55808;
    wire N__55805;
    wire N__55802;
    wire N__55801;
    wire N__55800;
    wire N__55799;
    wire N__55796;
    wire N__55793;
    wire N__55788;
    wire N__55783;
    wire N__55780;
    wire N__55777;
    wire N__55772;
    wire N__55769;
    wire N__55768;
    wire N__55767;
    wire N__55764;
    wire N__55761;
    wire N__55752;
    wire N__55749;
    wire N__55746;
    wire N__55743;
    wire N__55740;
    wire N__55737;
    wire N__55734;
    wire N__55727;
    wire N__55726;
    wire N__55725;
    wire N__55724;
    wire N__55721;
    wire N__55716;
    wire N__55713;
    wire N__55706;
    wire N__55697;
    wire N__55694;
    wire N__55691;
    wire N__55688;
    wire N__55687;
    wire N__55686;
    wire N__55685;
    wire N__55682;
    wire N__55681;
    wire N__55678;
    wire N__55675;
    wire N__55674;
    wire N__55671;
    wire N__55670;
    wire N__55665;
    wire N__55662;
    wire N__55661;
    wire N__55660;
    wire N__55657;
    wire N__55654;
    wire N__55651;
    wire N__55648;
    wire N__55647;
    wire N__55644;
    wire N__55641;
    wire N__55638;
    wire N__55635;
    wire N__55628;
    wire N__55625;
    wire N__55622;
    wire N__55619;
    wire N__55612;
    wire N__55609;
    wire N__55598;
    wire N__55595;
    wire N__55592;
    wire N__55589;
    wire N__55586;
    wire N__55585;
    wire N__55582;
    wire N__55579;
    wire N__55578;
    wire N__55577;
    wire N__55576;
    wire N__55573;
    wire N__55570;
    wire N__55565;
    wire N__55562;
    wire N__55559;
    wire N__55558;
    wire N__55555;
    wire N__55550;
    wire N__55549;
    wire N__55548;
    wire N__55547;
    wire N__55546;
    wire N__55543;
    wire N__55540;
    wire N__55535;
    wire N__55526;
    wire N__55517;
    wire N__55514;
    wire N__55511;
    wire N__55508;
    wire N__55505;
    wire N__55502;
    wire N__55499;
    wire N__55496;
    wire N__55493;
    wire N__55490;
    wire N__55487;
    wire N__55484;
    wire N__55481;
    wire N__55478;
    wire N__55475;
    wire N__55474;
    wire N__55473;
    wire N__55472;
    wire N__55471;
    wire N__55470;
    wire N__55467;
    wire N__55466;
    wire N__55465;
    wire N__55462;
    wire N__55457;
    wire N__55456;
    wire N__55455;
    wire N__55454;
    wire N__55453;
    wire N__55452;
    wire N__55451;
    wire N__55448;
    wire N__55445;
    wire N__55444;
    wire N__55441;
    wire N__55436;
    wire N__55431;
    wire N__55424;
    wire N__55423;
    wire N__55422;
    wire N__55421;
    wire N__55418;
    wire N__55413;
    wire N__55408;
    wire N__55405;
    wire N__55400;
    wire N__55399;
    wire N__55396;
    wire N__55393;
    wire N__55386;
    wire N__55381;
    wire N__55376;
    wire N__55373;
    wire N__55370;
    wire N__55365;
    wire N__55360;
    wire N__55357;
    wire N__55354;
    wire N__55351;
    wire N__55346;
    wire N__55343;
    wire N__55334;
    wire N__55333;
    wire N__55330;
    wire N__55327;
    wire N__55324;
    wire N__55321;
    wire N__55318;
    wire N__55315;
    wire N__55312;
    wire N__55309;
    wire N__55306;
    wire N__55301;
    wire N__55298;
    wire N__55295;
    wire N__55294;
    wire N__55291;
    wire N__55288;
    wire N__55283;
    wire N__55280;
    wire N__55277;
    wire N__55274;
    wire N__55271;
    wire N__55268;
    wire N__55265;
    wire N__55262;
    wire N__55259;
    wire N__55256;
    wire N__55253;
    wire N__55250;
    wire N__55247;
    wire N__55244;
    wire N__55241;
    wire N__55238;
    wire N__55235;
    wire N__55232;
    wire N__55229;
    wire N__55226;
    wire N__55223;
    wire N__55222;
    wire N__55221;
    wire N__55218;
    wire N__55215;
    wire N__55212;
    wire N__55205;
    wire N__55202;
    wire N__55199;
    wire N__55196;
    wire N__55193;
    wire N__55190;
    wire N__55187;
    wire N__55184;
    wire N__55183;
    wire N__55180;
    wire N__55177;
    wire N__55174;
    wire N__55169;
    wire N__55168;
    wire N__55167;
    wire N__55164;
    wire N__55159;
    wire N__55156;
    wire N__55155;
    wire N__55152;
    wire N__55149;
    wire N__55146;
    wire N__55139;
    wire N__55138;
    wire N__55137;
    wire N__55134;
    wire N__55131;
    wire N__55128;
    wire N__55125;
    wire N__55124;
    wire N__55123;
    wire N__55122;
    wire N__55121;
    wire N__55120;
    wire N__55119;
    wire N__55118;
    wire N__55115;
    wire N__55112;
    wire N__55109;
    wire N__55104;
    wire N__55099;
    wire N__55092;
    wire N__55079;
    wire N__55078;
    wire N__55077;
    wire N__55074;
    wire N__55071;
    wire N__55068;
    wire N__55065;
    wire N__55064;
    wire N__55059;
    wire N__55058;
    wire N__55057;
    wire N__55056;
    wire N__55055;
    wire N__55054;
    wire N__55053;
    wire N__55050;
    wire N__55047;
    wire N__55044;
    wire N__55041;
    wire N__55036;
    wire N__55033;
    wire N__55028;
    wire N__55013;
    wire N__55010;
    wire N__55007;
    wire N__55004;
    wire N__55001;
    wire N__54998;
    wire N__54995;
    wire N__54992;
    wire N__54989;
    wire N__54986;
    wire N__54983;
    wire N__54980;
    wire N__54977;
    wire N__54974;
    wire N__54971;
    wire N__54968;
    wire N__54965;
    wire N__54962;
    wire N__54959;
    wire N__54956;
    wire N__54953;
    wire N__54950;
    wire N__54947;
    wire N__54944;
    wire N__54941;
    wire N__54938;
    wire N__54935;
    wire N__54932;
    wire N__54929;
    wire N__54926;
    wire N__54923;
    wire N__54922;
    wire N__54919;
    wire N__54916;
    wire N__54913;
    wire N__54908;
    wire N__54905;
    wire N__54902;
    wire N__54901;
    wire N__54898;
    wire N__54895;
    wire N__54890;
    wire N__54889;
    wire N__54884;
    wire N__54881;
    wire N__54878;
    wire N__54875;
    wire N__54872;
    wire N__54869;
    wire N__54866;
    wire N__54863;
    wire N__54860;
    wire N__54857;
    wire N__54854;
    wire N__54851;
    wire N__54848;
    wire N__54845;
    wire N__54842;
    wire N__54839;
    wire N__54836;
    wire N__54833;
    wire N__54830;
    wire N__54827;
    wire N__54824;
    wire N__54821;
    wire N__54818;
    wire N__54815;
    wire N__54814;
    wire N__54811;
    wire N__54808;
    wire N__54803;
    wire N__54802;
    wire N__54799;
    wire N__54796;
    wire N__54791;
    wire N__54788;
    wire N__54785;
    wire N__54782;
    wire N__54779;
    wire N__54776;
    wire N__54773;
    wire N__54770;
    wire N__54767;
    wire N__54766;
    wire N__54763;
    wire N__54760;
    wire N__54757;
    wire N__54752;
    wire N__54751;
    wire N__54750;
    wire N__54747;
    wire N__54746;
    wire N__54741;
    wire N__54738;
    wire N__54735;
    wire N__54732;
    wire N__54729;
    wire N__54726;
    wire N__54723;
    wire N__54720;
    wire N__54719;
    wire N__54716;
    wire N__54711;
    wire N__54708;
    wire N__54707;
    wire N__54702;
    wire N__54699;
    wire N__54696;
    wire N__54689;
    wire N__54688;
    wire N__54687;
    wire N__54686;
    wire N__54685;
    wire N__54682;
    wire N__54681;
    wire N__54680;
    wire N__54679;
    wire N__54678;
    wire N__54677;
    wire N__54674;
    wire N__54671;
    wire N__54670;
    wire N__54669;
    wire N__54668;
    wire N__54665;
    wire N__54662;
    wire N__54661;
    wire N__54660;
    wire N__54659;
    wire N__54658;
    wire N__54657;
    wire N__54656;
    wire N__54655;
    wire N__54654;
    wire N__54653;
    wire N__54652;
    wire N__54651;
    wire N__54648;
    wire N__54641;
    wire N__54636;
    wire N__54635;
    wire N__54634;
    wire N__54633;
    wire N__54632;
    wire N__54627;
    wire N__54620;
    wire N__54615;
    wire N__54612;
    wire N__54609;
    wire N__54602;
    wire N__54599;
    wire N__54596;
    wire N__54593;
    wire N__54588;
    wire N__54587;
    wire N__54586;
    wire N__54585;
    wire N__54584;
    wire N__54583;
    wire N__54582;
    wire N__54581;
    wire N__54580;
    wire N__54579;
    wire N__54576;
    wire N__54575;
    wire N__54574;
    wire N__54573;
    wire N__54572;
    wire N__54571;
    wire N__54570;
    wire N__54569;
    wire N__54568;
    wire N__54563;
    wire N__54560;
    wire N__54553;
    wire N__54550;
    wire N__54545;
    wire N__54544;
    wire N__54543;
    wire N__54542;
    wire N__54541;
    wire N__54540;
    wire N__54539;
    wire N__54536;
    wire N__54531;
    wire N__54528;
    wire N__54519;
    wire N__54514;
    wire N__54511;
    wire N__54506;
    wire N__54501;
    wire N__54494;
    wire N__54491;
    wire N__54486;
    wire N__54477;
    wire N__54474;
    wire N__54469;
    wire N__54466;
    wire N__54461;
    wire N__54458;
    wire N__54453;
    wire N__54446;
    wire N__54435;
    wire N__54426;
    wire N__54401;
    wire N__54398;
    wire N__54395;
    wire N__54392;
    wire N__54389;
    wire N__54386;
    wire N__54383;
    wire N__54380;
    wire N__54377;
    wire N__54374;
    wire N__54371;
    wire N__54368;
    wire N__54365;
    wire N__54362;
    wire N__54359;
    wire N__54358;
    wire N__54357;
    wire N__54356;
    wire N__54355;
    wire N__54352;
    wire N__54343;
    wire N__54338;
    wire N__54335;
    wire N__54332;
    wire N__54329;
    wire N__54328;
    wire N__54323;
    wire N__54320;
    wire N__54317;
    wire N__54314;
    wire N__54311;
    wire N__54308;
    wire N__54305;
    wire N__54304;
    wire N__54303;
    wire N__54300;
    wire N__54299;
    wire N__54298;
    wire N__54297;
    wire N__54296;
    wire N__54295;
    wire N__54294;
    wire N__54293;
    wire N__54292;
    wire N__54289;
    wire N__54286;
    wire N__54285;
    wire N__54284;
    wire N__54281;
    wire N__54276;
    wire N__54271;
    wire N__54266;
    wire N__54261;
    wire N__54258;
    wire N__54255;
    wire N__54250;
    wire N__54249;
    wire N__54244;
    wire N__54237;
    wire N__54236;
    wire N__54235;
    wire N__54234;
    wire N__54231;
    wire N__54228;
    wire N__54225;
    wire N__54222;
    wire N__54217;
    wire N__54212;
    wire N__54209;
    wire N__54194;
    wire N__54191;
    wire N__54188;
    wire N__54187;
    wire N__54186;
    wire N__54183;
    wire N__54178;
    wire N__54175;
    wire N__54172;
    wire N__54169;
    wire N__54166;
    wire N__54161;
    wire N__54158;
    wire N__54155;
    wire N__54152;
    wire N__54149;
    wire N__54146;
    wire N__54143;
    wire N__54142;
    wire N__54141;
    wire N__54140;
    wire N__54139;
    wire N__54138;
    wire N__54135;
    wire N__54134;
    wire N__54131;
    wire N__54130;
    wire N__54129;
    wire N__54128;
    wire N__54125;
    wire N__54122;
    wire N__54119;
    wire N__54118;
    wire N__54115;
    wire N__54114;
    wire N__54113;
    wire N__54112;
    wire N__54111;
    wire N__54110;
    wire N__54107;
    wire N__54104;
    wire N__54101;
    wire N__54098;
    wire N__54093;
    wire N__54090;
    wire N__54085;
    wire N__54082;
    wire N__54079;
    wire N__54074;
    wire N__54069;
    wire N__54066;
    wire N__54063;
    wire N__54062;
    wire N__54061;
    wire N__54060;
    wire N__54059;
    wire N__54056;
    wire N__54047;
    wire N__54042;
    wire N__54041;
    wire N__54034;
    wire N__54029;
    wire N__54022;
    wire N__54019;
    wire N__54012;
    wire N__54009;
    wire N__54006;
    wire N__54001;
    wire N__53990;
    wire N__53987;
    wire N__53984;
    wire N__53981;
    wire N__53978;
    wire N__53975;
    wire N__53972;
    wire N__53969;
    wire N__53968;
    wire N__53967;
    wire N__53966;
    wire N__53965;
    wire N__53964;
    wire N__53963;
    wire N__53962;
    wire N__53961;
    wire N__53958;
    wire N__53957;
    wire N__53956;
    wire N__53953;
    wire N__53952;
    wire N__53951;
    wire N__53946;
    wire N__53943;
    wire N__53942;
    wire N__53941;
    wire N__53940;
    wire N__53939;
    wire N__53938;
    wire N__53937;
    wire N__53936;
    wire N__53931;
    wire N__53924;
    wire N__53919;
    wire N__53916;
    wire N__53911;
    wire N__53910;
    wire N__53909;
    wire N__53904;
    wire N__53899;
    wire N__53898;
    wire N__53895;
    wire N__53890;
    wire N__53889;
    wire N__53888;
    wire N__53887;
    wire N__53882;
    wire N__53879;
    wire N__53876;
    wire N__53873;
    wire N__53870;
    wire N__53867;
    wire N__53862;
    wire N__53861;
    wire N__53860;
    wire N__53859;
    wire N__53856;
    wire N__53853;
    wire N__53848;
    wire N__53845;
    wire N__53842;
    wire N__53837;
    wire N__53828;
    wire N__53823;
    wire N__53820;
    wire N__53817;
    wire N__53812;
    wire N__53805;
    wire N__53796;
    wire N__53783;
    wire N__53780;
    wire N__53777;
    wire N__53774;
    wire N__53771;
    wire N__53768;
    wire N__53765;
    wire N__53762;
    wire N__53759;
    wire N__53758;
    wire N__53757;
    wire N__53754;
    wire N__53749;
    wire N__53744;
    wire N__53741;
    wire N__53738;
    wire N__53735;
    wire N__53732;
    wire N__53729;
    wire N__53726;
    wire N__53723;
    wire N__53720;
    wire N__53719;
    wire N__53718;
    wire N__53717;
    wire N__53714;
    wire N__53709;
    wire N__53706;
    wire N__53705;
    wire N__53704;
    wire N__53701;
    wire N__53698;
    wire N__53691;
    wire N__53690;
    wire N__53689;
    wire N__53682;
    wire N__53677;
    wire N__53674;
    wire N__53669;
    wire N__53668;
    wire N__53667;
    wire N__53666;
    wire N__53663;
    wire N__53662;
    wire N__53661;
    wire N__53658;
    wire N__53653;
    wire N__53650;
    wire N__53645;
    wire N__53642;
    wire N__53639;
    wire N__53636;
    wire N__53627;
    wire N__53624;
    wire N__53621;
    wire N__53618;
    wire N__53615;
    wire N__53612;
    wire N__53611;
    wire N__53608;
    wire N__53605;
    wire N__53602;
    wire N__53599;
    wire N__53596;
    wire N__53593;
    wire N__53588;
    wire N__53585;
    wire N__53584;
    wire N__53583;
    wire N__53580;
    wire N__53575;
    wire N__53574;
    wire N__53573;
    wire N__53572;
    wire N__53571;
    wire N__53570;
    wire N__53567;
    wire N__53564;
    wire N__53561;
    wire N__53558;
    wire N__53555;
    wire N__53550;
    wire N__53545;
    wire N__53534;
    wire N__53531;
    wire N__53530;
    wire N__53527;
    wire N__53524;
    wire N__53521;
    wire N__53518;
    wire N__53517;
    wire N__53514;
    wire N__53511;
    wire N__53508;
    wire N__53505;
    wire N__53502;
    wire N__53499;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53485;
    wire N__53480;
    wire N__53479;
    wire N__53478;
    wire N__53477;
    wire N__53474;
    wire N__53471;
    wire N__53468;
    wire N__53467;
    wire N__53466;
    wire N__53463;
    wire N__53458;
    wire N__53455;
    wire N__53450;
    wire N__53445;
    wire N__53438;
    wire N__53435;
    wire N__53434;
    wire N__53431;
    wire N__53430;
    wire N__53429;
    wire N__53426;
    wire N__53425;
    wire N__53422;
    wire N__53417;
    wire N__53414;
    wire N__53411;
    wire N__53410;
    wire N__53407;
    wire N__53406;
    wire N__53405;
    wire N__53402;
    wire N__53401;
    wire N__53400;
    wire N__53395;
    wire N__53392;
    wire N__53389;
    wire N__53384;
    wire N__53381;
    wire N__53376;
    wire N__53363;
    wire N__53360;
    wire N__53357;
    wire N__53354;
    wire N__53351;
    wire N__53348;
    wire N__53345;
    wire N__53342;
    wire N__53339;
    wire N__53336;
    wire N__53333;
    wire N__53332;
    wire N__53329;
    wire N__53326;
    wire N__53323;
    wire N__53320;
    wire N__53317;
    wire N__53314;
    wire N__53309;
    wire N__53306;
    wire N__53305;
    wire N__53304;
    wire N__53303;
    wire N__53302;
    wire N__53301;
    wire N__53300;
    wire N__53299;
    wire N__53298;
    wire N__53297;
    wire N__53296;
    wire N__53295;
    wire N__53294;
    wire N__53293;
    wire N__53292;
    wire N__53291;
    wire N__53290;
    wire N__53289;
    wire N__53288;
    wire N__53285;
    wire N__53282;
    wire N__53275;
    wire N__53272;
    wire N__53267;
    wire N__53264;
    wire N__53259;
    wire N__53250;
    wire N__53249;
    wire N__53246;
    wire N__53245;
    wire N__53242;
    wire N__53239;
    wire N__53238;
    wire N__53237;
    wire N__53234;
    wire N__53233;
    wire N__53232;
    wire N__53231;
    wire N__53226;
    wire N__53223;
    wire N__53220;
    wire N__53217;
    wire N__53216;
    wire N__53209;
    wire N__53206;
    wire N__53205;
    wire N__53204;
    wire N__53201;
    wire N__53198;
    wire N__53195;
    wire N__53192;
    wire N__53187;
    wire N__53184;
    wire N__53181;
    wire N__53178;
    wire N__53177;
    wire N__53174;
    wire N__53171;
    wire N__53166;
    wire N__53165;
    wire N__53162;
    wire N__53161;
    wire N__53158;
    wire N__53155;
    wire N__53152;
    wire N__53147;
    wire N__53146;
    wire N__53145;
    wire N__53144;
    wire N__53141;
    wire N__53138;
    wire N__53133;
    wire N__53130;
    wire N__53127;
    wire N__53122;
    wire N__53119;
    wire N__53112;
    wire N__53109;
    wire N__53106;
    wire N__53103;
    wire N__53094;
    wire N__53089;
    wire N__53086;
    wire N__53079;
    wire N__53072;
    wire N__53067;
    wire N__53048;
    wire N__53045;
    wire N__53042;
    wire N__53039;
    wire N__53036;
    wire N__53033;
    wire N__53030;
    wire N__53027;
    wire N__53024;
    wire N__53021;
    wire N__53018;
    wire N__53015;
    wire N__53012;
    wire N__53011;
    wire N__53010;
    wire N__53009;
    wire N__53008;
    wire N__53007;
    wire N__53006;
    wire N__53003;
    wire N__53000;
    wire N__52997;
    wire N__52994;
    wire N__52991;
    wire N__52988;
    wire N__52987;
    wire N__52984;
    wire N__52981;
    wire N__52974;
    wire N__52971;
    wire N__52968;
    wire N__52965;
    wire N__52958;
    wire N__52953;
    wire N__52950;
    wire N__52947;
    wire N__52942;
    wire N__52937;
    wire N__52936;
    wire N__52935;
    wire N__52934;
    wire N__52933;
    wire N__52932;
    wire N__52931;
    wire N__52928;
    wire N__52925;
    wire N__52922;
    wire N__52919;
    wire N__52916;
    wire N__52913;
    wire N__52910;
    wire N__52905;
    wire N__52902;
    wire N__52889;
    wire N__52886;
    wire N__52883;
    wire N__52880;
    wire N__52879;
    wire N__52878;
    wire N__52875;
    wire N__52872;
    wire N__52871;
    wire N__52870;
    wire N__52867;
    wire N__52866;
    wire N__52863;
    wire N__52860;
    wire N__52857;
    wire N__52856;
    wire N__52853;
    wire N__52850;
    wire N__52847;
    wire N__52844;
    wire N__52839;
    wire N__52836;
    wire N__52833;
    wire N__52830;
    wire N__52825;
    wire N__52822;
    wire N__52813;
    wire N__52808;
    wire N__52807;
    wire N__52806;
    wire N__52805;
    wire N__52802;
    wire N__52801;
    wire N__52798;
    wire N__52795;
    wire N__52792;
    wire N__52789;
    wire N__52788;
    wire N__52787;
    wire N__52786;
    wire N__52783;
    wire N__52780;
    wire N__52777;
    wire N__52772;
    wire N__52769;
    wire N__52766;
    wire N__52763;
    wire N__52754;
    wire N__52745;
    wire N__52744;
    wire N__52741;
    wire N__52738;
    wire N__52735;
    wire N__52732;
    wire N__52729;
    wire N__52726;
    wire N__52723;
    wire N__52720;
    wire N__52717;
    wire N__52714;
    wire N__52709;
    wire N__52706;
    wire N__52705;
    wire N__52702;
    wire N__52699;
    wire N__52696;
    wire N__52691;
    wire N__52688;
    wire N__52685;
    wire N__52684;
    wire N__52683;
    wire N__52680;
    wire N__52679;
    wire N__52678;
    wire N__52675;
    wire N__52672;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52660;
    wire N__52657;
    wire N__52654;
    wire N__52645;
    wire N__52640;
    wire N__52637;
    wire N__52636;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52628;
    wire N__52627;
    wire N__52624;
    wire N__52623;
    wire N__52620;
    wire N__52619;
    wire N__52616;
    wire N__52613;
    wire N__52612;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52600;
    wire N__52597;
    wire N__52592;
    wire N__52589;
    wire N__52586;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52572;
    wire N__52565;
    wire N__52562;
    wire N__52559;
    wire N__52556;
    wire N__52553;
    wire N__52548;
    wire N__52541;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52531;
    wire N__52528;
    wire N__52527;
    wire N__52524;
    wire N__52521;
    wire N__52518;
    wire N__52515;
    wire N__52510;
    wire N__52507;
    wire N__52504;
    wire N__52499;
    wire N__52496;
    wire N__52493;
    wire N__52490;
    wire N__52487;
    wire N__52484;
    wire N__52481;
    wire N__52478;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52462;
    wire N__52459;
    wire N__52456;
    wire N__52451;
    wire N__52448;
    wire N__52447;
    wire N__52444;
    wire N__52441;
    wire N__52438;
    wire N__52435;
    wire N__52432;
    wire N__52429;
    wire N__52426;
    wire N__52423;
    wire N__52420;
    wire N__52417;
    wire N__52412;
    wire N__52411;
    wire N__52410;
    wire N__52407;
    wire N__52404;
    wire N__52401;
    wire N__52398;
    wire N__52395;
    wire N__52392;
    wire N__52389;
    wire N__52386;
    wire N__52383;
    wire N__52380;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52366;
    wire N__52363;
    wire N__52358;
    wire N__52357;
    wire N__52354;
    wire N__52351;
    wire N__52350;
    wire N__52347;
    wire N__52344;
    wire N__52341;
    wire N__52338;
    wire N__52335;
    wire N__52332;
    wire N__52329;
    wire N__52326;
    wire N__52323;
    wire N__52320;
    wire N__52315;
    wire N__52312;
    wire N__52307;
    wire N__52304;
    wire N__52301;
    wire N__52298;
    wire N__52295;
    wire N__52292;
    wire N__52291;
    wire N__52288;
    wire N__52285;
    wire N__52284;
    wire N__52281;
    wire N__52278;
    wire N__52275;
    wire N__52270;
    wire N__52267;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52252;
    wire N__52247;
    wire N__52246;
    wire N__52245;
    wire N__52242;
    wire N__52241;
    wire N__52240;
    wire N__52237;
    wire N__52236;
    wire N__52233;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52223;
    wire N__52220;
    wire N__52217;
    wire N__52214;
    wire N__52211;
    wire N__52206;
    wire N__52205;
    wire N__52202;
    wire N__52199;
    wire N__52196;
    wire N__52189;
    wire N__52186;
    wire N__52183;
    wire N__52178;
    wire N__52175;
    wire N__52166;
    wire N__52165;
    wire N__52162;
    wire N__52159;
    wire N__52156;
    wire N__52153;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52141;
    wire N__52138;
    wire N__52135;
    wire N__52132;
    wire N__52129;
    wire N__52124;
    wire N__52123;
    wire N__52122;
    wire N__52119;
    wire N__52118;
    wire N__52117;
    wire N__52114;
    wire N__52111;
    wire N__52108;
    wire N__52105;
    wire N__52102;
    wire N__52097;
    wire N__52096;
    wire N__52093;
    wire N__52090;
    wire N__52087;
    wire N__52084;
    wire N__52081;
    wire N__52080;
    wire N__52077;
    wire N__52072;
    wire N__52067;
    wire N__52064;
    wire N__52055;
    wire N__52054;
    wire N__52053;
    wire N__52052;
    wire N__52051;
    wire N__52050;
    wire N__52049;
    wire N__52046;
    wire N__52043;
    wire N__52040;
    wire N__52037;
    wire N__52034;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52024;
    wire N__52021;
    wire N__52014;
    wire N__52011;
    wire N__52008;
    wire N__52005;
    wire N__52002;
    wire N__51999;
    wire N__51996;
    wire N__51989;
    wire N__51986;
    wire N__51981;
    wire N__51978;
    wire N__51971;
    wire N__51968;
    wire N__51967;
    wire N__51964;
    wire N__51961;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51949;
    wire N__51946;
    wire N__51941;
    wire N__51938;
    wire N__51937;
    wire N__51934;
    wire N__51933;
    wire N__51932;
    wire N__51931;
    wire N__51930;
    wire N__51929;
    wire N__51926;
    wire N__51923;
    wire N__51920;
    wire N__51917;
    wire N__51914;
    wire N__51911;
    wire N__51908;
    wire N__51905;
    wire N__51904;
    wire N__51901;
    wire N__51898;
    wire N__51893;
    wire N__51886;
    wire N__51883;
    wire N__51880;
    wire N__51875;
    wire N__51872;
    wire N__51863;
    wire N__51862;
    wire N__51859;
    wire N__51858;
    wire N__51857;
    wire N__51854;
    wire N__51853;
    wire N__51852;
    wire N__51851;
    wire N__51848;
    wire N__51845;
    wire N__51842;
    wire N__51839;
    wire N__51836;
    wire N__51833;
    wire N__51830;
    wire N__51827;
    wire N__51824;
    wire N__51819;
    wire N__51806;
    wire N__51805;
    wire N__51802;
    wire N__51799;
    wire N__51794;
    wire N__51791;
    wire N__51788;
    wire N__51785;
    wire N__51784;
    wire N__51783;
    wire N__51780;
    wire N__51779;
    wire N__51778;
    wire N__51777;
    wire N__51776;
    wire N__51775;
    wire N__51772;
    wire N__51769;
    wire N__51766;
    wire N__51763;
    wire N__51760;
    wire N__51757;
    wire N__51754;
    wire N__51751;
    wire N__51748;
    wire N__51743;
    wire N__51728;
    wire N__51727;
    wire N__51724;
    wire N__51723;
    wire N__51722;
    wire N__51721;
    wire N__51720;
    wire N__51717;
    wire N__51714;
    wire N__51711;
    wire N__51708;
    wire N__51705;
    wire N__51704;
    wire N__51703;
    wire N__51700;
    wire N__51695;
    wire N__51692;
    wire N__51689;
    wire N__51686;
    wire N__51683;
    wire N__51680;
    wire N__51677;
    wire N__51674;
    wire N__51669;
    wire N__51660;
    wire N__51657;
    wire N__51654;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51638;
    wire N__51637;
    wire N__51636;
    wire N__51635;
    wire N__51634;
    wire N__51633;
    wire N__51632;
    wire N__51629;
    wire N__51626;
    wire N__51623;
    wire N__51620;
    wire N__51617;
    wire N__51614;
    wire N__51611;
    wire N__51608;
    wire N__51605;
    wire N__51602;
    wire N__51587;
    wire N__51584;
    wire N__51581;
    wire N__51580;
    wire N__51577;
    wire N__51574;
    wire N__51571;
    wire N__51568;
    wire N__51565;
    wire N__51562;
    wire N__51559;
    wire N__51554;
    wire N__51551;
    wire N__51548;
    wire N__51545;
    wire N__51542;
    wire N__51541;
    wire N__51538;
    wire N__51535;
    wire N__51532;
    wire N__51529;
    wire N__51526;
    wire N__51523;
    wire N__51520;
    wire N__51515;
    wire N__51512;
    wire N__51509;
    wire N__51506;
    wire N__51503;
    wire N__51502;
    wire N__51499;
    wire N__51496;
    wire N__51491;
    wire N__51490;
    wire N__51487;
    wire N__51484;
    wire N__51481;
    wire N__51478;
    wire N__51475;
    wire N__51472;
    wire N__51469;
    wire N__51466;
    wire N__51461;
    wire N__51458;
    wire N__51455;
    wire N__51452;
    wire N__51449;
    wire N__51446;
    wire N__51443;
    wire N__51440;
    wire N__51437;
    wire N__51434;
    wire N__51431;
    wire N__51428;
    wire N__51425;
    wire N__51422;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51406;
    wire N__51403;
    wire N__51400;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51388;
    wire N__51385;
    wire N__51382;
    wire N__51377;
    wire N__51374;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51356;
    wire N__51353;
    wire N__51350;
    wire N__51347;
    wire N__51344;
    wire N__51341;
    wire N__51338;
    wire N__51335;
    wire N__51334;
    wire N__51331;
    wire N__51328;
    wire N__51323;
    wire N__51322;
    wire N__51319;
    wire N__51316;
    wire N__51313;
    wire N__51310;
    wire N__51307;
    wire N__51304;
    wire N__51301;
    wire N__51296;
    wire N__51295;
    wire N__51292;
    wire N__51289;
    wire N__51286;
    wire N__51283;
    wire N__51280;
    wire N__51277;
    wire N__51272;
    wire N__51269;
    wire N__51266;
    wire N__51263;
    wire N__51262;
    wire N__51259;
    wire N__51256;
    wire N__51253;
    wire N__51248;
    wire N__51245;
    wire N__51242;
    wire N__51239;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51223;
    wire N__51220;
    wire N__51217;
    wire N__51214;
    wire N__51211;
    wire N__51206;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51182;
    wire N__51179;
    wire N__51176;
    wire N__51173;
    wire N__51170;
    wire N__51167;
    wire N__51164;
    wire N__51161;
    wire N__51158;
    wire N__51155;
    wire N__51152;
    wire N__51149;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51133;
    wire N__51130;
    wire N__51125;
    wire N__51122;
    wire N__51121;
    wire N__51118;
    wire N__51115;
    wire N__51110;
    wire N__51107;
    wire N__51104;
    wire N__51101;
    wire N__51098;
    wire N__51095;
    wire N__51092;
    wire N__51089;
    wire N__51086;
    wire N__51083;
    wire N__51080;
    wire N__51077;
    wire N__51074;
    wire N__51071;
    wire N__51068;
    wire N__51065;
    wire N__51064;
    wire N__51059;
    wire N__51056;
    wire N__51053;
    wire N__51050;
    wire N__51047;
    wire N__51044;
    wire N__51041;
    wire N__51038;
    wire N__51035;
    wire N__51032;
    wire N__51029;
    wire N__51026;
    wire N__51023;
    wire N__51020;
    wire N__51017;
    wire N__51014;
    wire N__51011;
    wire N__51008;
    wire N__51005;
    wire N__51002;
    wire N__50999;
    wire N__50996;
    wire N__50993;
    wire N__50990;
    wire N__50987;
    wire N__50986;
    wire N__50983;
    wire N__50980;
    wire N__50977;
    wire N__50974;
    wire N__50969;
    wire N__50966;
    wire N__50963;
    wire N__50962;
    wire N__50959;
    wire N__50956;
    wire N__50955;
    wire N__50952;
    wire N__50949;
    wire N__50948;
    wire N__50947;
    wire N__50944;
    wire N__50941;
    wire N__50938;
    wire N__50935;
    wire N__50932;
    wire N__50921;
    wire N__50918;
    wire N__50915;
    wire N__50912;
    wire N__50909;
    wire N__50906;
    wire N__50905;
    wire N__50904;
    wire N__50903;
    wire N__50900;
    wire N__50899;
    wire N__50898;
    wire N__50893;
    wire N__50890;
    wire N__50887;
    wire N__50884;
    wire N__50881;
    wire N__50876;
    wire N__50873;
    wire N__50872;
    wire N__50871;
    wire N__50866;
    wire N__50863;
    wire N__50860;
    wire N__50855;
    wire N__50850;
    wire N__50843;
    wire N__50842;
    wire N__50841;
    wire N__50838;
    wire N__50837;
    wire N__50836;
    wire N__50835;
    wire N__50834;
    wire N__50831;
    wire N__50830;
    wire N__50827;
    wire N__50822;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50808;
    wire N__50805;
    wire N__50800;
    wire N__50797;
    wire N__50794;
    wire N__50791;
    wire N__50788;
    wire N__50785;
    wire N__50782;
    wire N__50775;
    wire N__50772;
    wire N__50767;
    wire N__50764;
    wire N__50759;
    wire N__50756;
    wire N__50753;
    wire N__50750;
    wire N__50747;
    wire N__50744;
    wire N__50741;
    wire N__50738;
    wire N__50735;
    wire N__50732;
    wire N__50729;
    wire N__50726;
    wire N__50723;
    wire N__50720;
    wire N__50717;
    wire N__50714;
    wire N__50713;
    wire N__50710;
    wire N__50707;
    wire N__50704;
    wire N__50701;
    wire N__50696;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50684;
    wire N__50681;
    wire N__50678;
    wire N__50675;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50662;
    wire N__50659;
    wire N__50656;
    wire N__50651;
    wire N__50648;
    wire N__50645;
    wire N__50642;
    wire N__50639;
    wire N__50636;
    wire N__50633;
    wire N__50630;
    wire N__50627;
    wire N__50624;
    wire N__50621;
    wire N__50620;
    wire N__50617;
    wire N__50612;
    wire N__50609;
    wire N__50606;
    wire N__50603;
    wire N__50600;
    wire N__50597;
    wire N__50594;
    wire N__50591;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50579;
    wire N__50576;
    wire N__50573;
    wire N__50572;
    wire N__50569;
    wire N__50566;
    wire N__50561;
    wire N__50558;
    wire N__50555;
    wire N__50552;
    wire N__50549;
    wire N__50546;
    wire N__50543;
    wire N__50542;
    wire N__50541;
    wire N__50538;
    wire N__50537;
    wire N__50532;
    wire N__50527;
    wire N__50524;
    wire N__50521;
    wire N__50516;
    wire N__50513;
    wire N__50512;
    wire N__50507;
    wire N__50504;
    wire N__50501;
    wire N__50498;
    wire N__50495;
    wire N__50494;
    wire N__50491;
    wire N__50488;
    wire N__50487;
    wire N__50486;
    wire N__50477;
    wire N__50474;
    wire N__50471;
    wire N__50470;
    wire N__50467;
    wire N__50464;
    wire N__50461;
    wire N__50458;
    wire N__50455;
    wire N__50452;
    wire N__50447;
    wire N__50444;
    wire N__50441;
    wire N__50438;
    wire N__50435;
    wire N__50432;
    wire N__50431;
    wire N__50430;
    wire N__50427;
    wire N__50422;
    wire N__50417;
    wire N__50414;
    wire N__50411;
    wire N__50408;
    wire N__50405;
    wire N__50404;
    wire N__50401;
    wire N__50400;
    wire N__50397;
    wire N__50394;
    wire N__50389;
    wire N__50386;
    wire N__50383;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50354;
    wire N__50351;
    wire N__50348;
    wire N__50345;
    wire N__50342;
    wire N__50341;
    wire N__50338;
    wire N__50337;
    wire N__50334;
    wire N__50331;
    wire N__50328;
    wire N__50327;
    wire N__50326;
    wire N__50325;
    wire N__50324;
    wire N__50321;
    wire N__50318;
    wire N__50315;
    wire N__50312;
    wire N__50309;
    wire N__50306;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50298;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50280;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50266;
    wire N__50259;
    wire N__50256;
    wire N__50243;
    wire N__50240;
    wire N__50237;
    wire N__50234;
    wire N__50231;
    wire N__50228;
    wire N__50225;
    wire N__50224;
    wire N__50223;
    wire N__50222;
    wire N__50221;
    wire N__50220;
    wire N__50219;
    wire N__50218;
    wire N__50217;
    wire N__50216;
    wire N__50215;
    wire N__50214;
    wire N__50213;
    wire N__50204;
    wire N__50203;
    wire N__50202;
    wire N__50201;
    wire N__50200;
    wire N__50199;
    wire N__50198;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50190;
    wire N__50187;
    wire N__50186;
    wire N__50183;
    wire N__50178;
    wire N__50175;
    wire N__50172;
    wire N__50169;
    wire N__50168;
    wire N__50165;
    wire N__50158;
    wire N__50157;
    wire N__50156;
    wire N__50155;
    wire N__50154;
    wire N__50153;
    wire N__50152;
    wire N__50149;
    wire N__50148;
    wire N__50147;
    wire N__50144;
    wire N__50143;
    wire N__50138;
    wire N__50133;
    wire N__50132;
    wire N__50131;
    wire N__50128;
    wire N__50127;
    wire N__50126;
    wire N__50125;
    wire N__50124;
    wire N__50123;
    wire N__50120;
    wire N__50117;
    wire N__50114;
    wire N__50113;
    wire N__50112;
    wire N__50111;
    wire N__50108;
    wire N__50107;
    wire N__50106;
    wire N__50105;
    wire N__50104;
    wire N__50103;
    wire N__50102;
    wire N__50095;
    wire N__50092;
    wire N__50087;
    wire N__50084;
    wire N__50077;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50063;
    wire N__50060;
    wire N__50057;
    wire N__50052;
    wire N__50047;
    wire N__50044;
    wire N__50041;
    wire N__50032;
    wire N__50029;
    wire N__50026;
    wire N__50023;
    wire N__50022;
    wire N__50021;
    wire N__50020;
    wire N__50019;
    wire N__50012;
    wire N__50011;
    wire N__50010;
    wire N__50009;
    wire N__50008;
    wire N__50007;
    wire N__50006;
    wire N__50005;
    wire N__50004;
    wire N__50003;
    wire N__50000;
    wire N__49991;
    wire N__49986;
    wire N__49979;
    wire N__49974;
    wire N__49969;
    wire N__49956;
    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49946;
    wire N__49945;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49939;
    wire N__49934;
    wire N__49925;
    wire N__49922;
    wire N__49911;
    wire N__49902;
    wire N__49893;
    wire N__49888;
    wire N__49883;
    wire N__49880;
    wire N__49867;
    wire N__49844;
    wire N__49841;
    wire N__49838;
    wire N__49835;
    wire N__49832;
    wire N__49831;
    wire N__49830;
    wire N__49829;
    wire N__49826;
    wire N__49825;
    wire N__49824;
    wire N__49819;
    wire N__49818;
    wire N__49817;
    wire N__49816;
    wire N__49815;
    wire N__49812;
    wire N__49811;
    wire N__49810;
    wire N__49807;
    wire N__49806;
    wire N__49803;
    wire N__49802;
    wire N__49799;
    wire N__49798;
    wire N__49797;
    wire N__49794;
    wire N__49793;
    wire N__49790;
    wire N__49787;
    wire N__49786;
    wire N__49785;
    wire N__49780;
    wire N__49777;
    wire N__49774;
    wire N__49771;
    wire N__49768;
    wire N__49765;
    wire N__49762;
    wire N__49759;
    wire N__49758;
    wire N__49755;
    wire N__49752;
    wire N__49749;
    wire N__49746;
    wire N__49743;
    wire N__49742;
    wire N__49739;
    wire N__49736;
    wire N__49733;
    wire N__49730;
    wire N__49727;
    wire N__49724;
    wire N__49719;
    wire N__49712;
    wire N__49711;
    wire N__49710;
    wire N__49709;
    wire N__49706;
    wire N__49703;
    wire N__49700;
    wire N__49697;
    wire N__49690;
    wire N__49687;
    wire N__49684;
    wire N__49681;
    wire N__49678;
    wire N__49675;
    wire N__49666;
    wire N__49659;
    wire N__49652;
    wire N__49647;
    wire N__49628;
    wire N__49625;
    wire N__49622;
    wire N__49619;
    wire N__49616;
    wire N__49613;
    wire N__49610;
    wire N__49607;
    wire N__49606;
    wire N__49605;
    wire N__49604;
    wire N__49601;
    wire N__49600;
    wire N__49597;
    wire N__49596;
    wire N__49595;
    wire N__49594;
    wire N__49593;
    wire N__49592;
    wire N__49589;
    wire N__49588;
    wire N__49587;
    wire N__49584;
    wire N__49583;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49579;
    wire N__49578;
    wire N__49577;
    wire N__49576;
    wire N__49575;
    wire N__49574;
    wire N__49573;
    wire N__49572;
    wire N__49569;
    wire N__49564;
    wire N__49563;
    wire N__49562;
    wire N__49561;
    wire N__49554;
    wire N__49553;
    wire N__49552;
    wire N__49547;
    wire N__49546;
    wire N__49545;
    wire N__49544;
    wire N__49541;
    wire N__49538;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49529;
    wire N__49528;
    wire N__49525;
    wire N__49524;
    wire N__49523;
    wire N__49520;
    wire N__49519;
    wire N__49516;
    wire N__49513;
    wire N__49512;
    wire N__49509;
    wire N__49506;
    wire N__49505;
    wire N__49502;
    wire N__49501;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49493;
    wire N__49486;
    wire N__49481;
    wire N__49478;
    wire N__49475;
    wire N__49472;
    wire N__49469;
    wire N__49464;
    wire N__49461;
    wire N__49456;
    wire N__49453;
    wire N__49450;
    wire N__49445;
    wire N__49438;
    wire N__49435;
    wire N__49432;
    wire N__49431;
    wire N__49428;
    wire N__49423;
    wire N__49418;
    wire N__49413;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49399;
    wire N__49396;
    wire N__49393;
    wire N__49392;
    wire N__49391;
    wire N__49384;
    wire N__49375;
    wire N__49370;
    wire N__49367;
    wire N__49364;
    wire N__49361;
    wire N__49354;
    wire N__49351;
    wire N__49348;
    wire N__49343;
    wire N__49342;
    wire N__49341;
    wire N__49340;
    wire N__49339;
    wire N__49334;
    wire N__49331;
    wire N__49324;
    wire N__49323;
    wire N__49322;
    wire N__49321;
    wire N__49320;
    wire N__49317;
    wire N__49312;
    wire N__49309;
    wire N__49304;
    wire N__49295;
    wire N__49286;
    wire N__49281;
    wire N__49272;
    wire N__49269;
    wire N__49264;
    wire N__49255;
    wire N__49232;
    wire N__49229;
    wire N__49226;
    wire N__49223;
    wire N__49220;
    wire N__49219;
    wire N__49216;
    wire N__49213;
    wire N__49210;
    wire N__49207;
    wire N__49204;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49194;
    wire N__49189;
    wire N__49186;
    wire N__49181;
    wire N__49178;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49168;
    wire N__49165;
    wire N__49164;
    wire N__49159;
    wire N__49156;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49139;
    wire N__49136;
    wire N__49133;
    wire N__49132;
    wire N__49131;
    wire N__49128;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49108;
    wire N__49105;
    wire N__49102;
    wire N__49097;
    wire N__49094;
    wire N__49091;
    wire N__49088;
    wire N__49085;
    wire N__49082;
    wire N__49081;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49071;
    wire N__49068;
    wire N__49063;
    wire N__49058;
    wire N__49055;
    wire N__49052;
    wire N__49049;
    wire N__49046;
    wire N__49045;
    wire N__49044;
    wire N__49041;
    wire N__49038;
    wire N__49035;
    wire N__49030;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49009;
    wire N__49006;
    wire N__49003;
    wire N__48998;
    wire N__48995;
    wire N__48992;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48981;
    wire N__48978;
    wire N__48975;
    wire N__48972;
    wire N__48969;
    wire N__48966;
    wire N__48963;
    wire N__48960;
    wire N__48955;
    wire N__48950;
    wire N__48947;
    wire N__48944;
    wire N__48943;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48933;
    wire N__48928;
    wire N__48925;
    wire N__48920;
    wire N__48917;
    wire N__48914;
    wire N__48911;
    wire N__48908;
    wire N__48905;
    wire N__48902;
    wire N__48901;
    wire N__48900;
    wire N__48897;
    wire N__48894;
    wire N__48891;
    wire N__48886;
    wire N__48883;
    wire N__48878;
    wire N__48875;
    wire N__48872;
    wire N__48871;
    wire N__48868;
    wire N__48867;
    wire N__48864;
    wire N__48861;
    wire N__48858;
    wire N__48855;
    wire N__48852;
    wire N__48849;
    wire N__48846;
    wire N__48843;
    wire N__48838;
    wire N__48833;
    wire N__48832;
    wire N__48829;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48814;
    wire N__48811;
    wire N__48806;
    wire N__48803;
    wire N__48800;
    wire N__48797;
    wire N__48794;
    wire N__48791;
    wire N__48790;
    wire N__48787;
    wire N__48784;
    wire N__48779;
    wire N__48776;
    wire N__48773;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48755;
    wire N__48752;
    wire N__48749;
    wire N__48746;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48727;
    wire N__48724;
    wire N__48719;
    wire N__48716;
    wire N__48713;
    wire N__48710;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48680;
    wire N__48677;
    wire N__48674;
    wire N__48673;
    wire N__48672;
    wire N__48669;
    wire N__48666;
    wire N__48663;
    wire N__48660;
    wire N__48657;
    wire N__48654;
    wire N__48651;
    wire N__48648;
    wire N__48645;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48631;
    wire N__48626;
    wire N__48623;
    wire N__48620;
    wire N__48617;
    wire N__48614;
    wire N__48611;
    wire N__48610;
    wire N__48607;
    wire N__48604;
    wire N__48599;
    wire N__48596;
    wire N__48595;
    wire N__48592;
    wire N__48589;
    wire N__48584;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48554;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48539;
    wire N__48536;
    wire N__48535;
    wire N__48532;
    wire N__48529;
    wire N__48526;
    wire N__48523;
    wire N__48518;
    wire N__48515;
    wire N__48512;
    wire N__48509;
    wire N__48506;
    wire N__48503;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48491;
    wire N__48488;
    wire N__48487;
    wire N__48484;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48468;
    wire N__48465;
    wire N__48464;
    wire N__48463;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48440;
    wire N__48435;
    wire N__48428;
    wire N__48425;
    wire N__48422;
    wire N__48419;
    wire N__48416;
    wire N__48413;
    wire N__48410;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48392;
    wire N__48389;
    wire N__48386;
    wire N__48383;
    wire N__48380;
    wire N__48377;
    wire N__48376;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48364;
    wire N__48361;
    wire N__48358;
    wire N__48353;
    wire N__48350;
    wire N__48347;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48335;
    wire N__48332;
    wire N__48329;
    wire N__48326;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48316;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48290;
    wire N__48287;
    wire N__48284;
    wire N__48281;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48265;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48242;
    wire N__48239;
    wire N__48236;
    wire N__48233;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48212;
    wire N__48209;
    wire N__48206;
    wire N__48203;
    wire N__48200;
    wire N__48197;
    wire N__48194;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48179;
    wire N__48176;
    wire N__48175;
    wire N__48174;
    wire N__48171;
    wire N__48166;
    wire N__48163;
    wire N__48158;
    wire N__48155;
    wire N__48152;
    wire N__48149;
    wire N__48146;
    wire N__48143;
    wire N__48142;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48132;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48097;
    wire N__48092;
    wire N__48089;
    wire N__48086;
    wire N__48083;
    wire N__48082;
    wire N__48079;
    wire N__48076;
    wire N__48073;
    wire N__48068;
    wire N__48065;
    wire N__48062;
    wire N__48059;
    wire N__48058;
    wire N__48055;
    wire N__48052;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48032;
    wire N__48029;
    wire N__48026;
    wire N__48023;
    wire N__48020;
    wire N__48017;
    wire N__48016;
    wire N__48015;
    wire N__48012;
    wire N__48007;
    wire N__48002;
    wire N__47999;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47986;
    wire N__47985;
    wire N__47982;
    wire N__47979;
    wire N__47978;
    wire N__47975;
    wire N__47972;
    wire N__47969;
    wire N__47966;
    wire N__47963;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47949;
    wire N__47942;
    wire N__47939;
    wire N__47936;
    wire N__47933;
    wire N__47930;
    wire N__47927;
    wire N__47924;
    wire N__47921;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47864;
    wire N__47861;
    wire N__47858;
    wire N__47855;
    wire N__47852;
    wire N__47849;
    wire N__47846;
    wire N__47843;
    wire N__47840;
    wire N__47839;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47824;
    wire N__47821;
    wire N__47816;
    wire N__47813;
    wire N__47810;
    wire N__47807;
    wire N__47804;
    wire N__47801;
    wire N__47798;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47786;
    wire N__47783;
    wire N__47780;
    wire N__47777;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47723;
    wire N__47720;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47690;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47680;
    wire N__47677;
    wire N__47674;
    wire N__47669;
    wire N__47666;
    wire N__47663;
    wire N__47660;
    wire N__47657;
    wire N__47654;
    wire N__47651;
    wire N__47648;
    wire N__47645;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47600;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47588;
    wire N__47585;
    wire N__47582;
    wire N__47579;
    wire N__47576;
    wire N__47573;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47552;
    wire N__47549;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47524;
    wire N__47523;
    wire N__47518;
    wire N__47515;
    wire N__47514;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47495;
    wire N__47494;
    wire N__47491;
    wire N__47490;
    wire N__47489;
    wire N__47488;
    wire N__47485;
    wire N__47478;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47456;
    wire N__47453;
    wire N__47450;
    wire N__47447;
    wire N__47442;
    wire N__47437;
    wire N__47434;
    wire N__47429;
    wire N__47426;
    wire N__47423;
    wire N__47420;
    wire N__47417;
    wire N__47414;
    wire N__47411;
    wire N__47408;
    wire N__47407;
    wire N__47404;
    wire N__47403;
    wire N__47400;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47383;
    wire N__47380;
    wire N__47377;
    wire N__47372;
    wire N__47369;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47321;
    wire N__47318;
    wire N__47315;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47296;
    wire N__47293;
    wire N__47288;
    wire N__47285;
    wire N__47284;
    wire N__47281;
    wire N__47278;
    wire N__47277;
    wire N__47276;
    wire N__47275;
    wire N__47274;
    wire N__47273;
    wire N__47272;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47260;
    wire N__47255;
    wire N__47250;
    wire N__47247;
    wire N__47246;
    wire N__47243;
    wire N__47240;
    wire N__47237;
    wire N__47232;
    wire N__47227;
    wire N__47216;
    wire N__47213;
    wire N__47212;
    wire N__47211;
    wire N__47210;
    wire N__47205;
    wire N__47204;
    wire N__47203;
    wire N__47202;
    wire N__47201;
    wire N__47196;
    wire N__47195;
    wire N__47194;
    wire N__47193;
    wire N__47192;
    wire N__47191;
    wire N__47190;
    wire N__47189;
    wire N__47188;
    wire N__47185;
    wire N__47180;
    wire N__47175;
    wire N__47172;
    wire N__47167;
    wire N__47162;
    wire N__47157;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47145;
    wire N__47144;
    wire N__47143;
    wire N__47142;
    wire N__47139;
    wire N__47136;
    wire N__47133;
    wire N__47128;
    wire N__47121;
    wire N__47112;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47084;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47062;
    wire N__47059;
    wire N__47056;
    wire N__47051;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47033;
    wire N__47030;
    wire N__47025;
    wire N__47022;
    wire N__47015;
    wire N__47012;
    wire N__47011;
    wire N__47010;
    wire N__47009;
    wire N__47006;
    wire N__47003;
    wire N__47002;
    wire N__46997;
    wire N__46994;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46984;
    wire N__46981;
    wire N__46974;
    wire N__46971;
    wire N__46964;
    wire N__46961;
    wire N__46958;
    wire N__46955;
    wire N__46952;
    wire N__46949;
    wire N__46946;
    wire N__46945;
    wire N__46944;
    wire N__46943;
    wire N__46942;
    wire N__46939;
    wire N__46936;
    wire N__46935;
    wire N__46932;
    wire N__46927;
    wire N__46926;
    wire N__46925;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46919;
    wire N__46914;
    wire N__46909;
    wire N__46904;
    wire N__46899;
    wire N__46898;
    wire N__46897;
    wire N__46896;
    wire N__46893;
    wire N__46892;
    wire N__46889;
    wire N__46884;
    wire N__46881;
    wire N__46878;
    wire N__46871;
    wire N__46866;
    wire N__46859;
    wire N__46850;
    wire N__46847;
    wire N__46844;
    wire N__46841;
    wire N__46840;
    wire N__46837;
    wire N__46836;
    wire N__46833;
    wire N__46832;
    wire N__46831;
    wire N__46828;
    wire N__46827;
    wire N__46824;
    wire N__46821;
    wire N__46816;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46808;
    wire N__46805;
    wire N__46798;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46782;
    wire N__46781;
    wire N__46780;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46756;
    wire N__46753;
    wire N__46746;
    wire N__46733;
    wire N__46730;
    wire N__46727;
    wire N__46724;
    wire N__46721;
    wire N__46718;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46700;
    wire N__46697;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46685;
    wire N__46684;
    wire N__46679;
    wire N__46676;
    wire N__46673;
    wire N__46670;
    wire N__46667;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46655;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46591;
    wire N__46586;
    wire N__46583;
    wire N__46580;
    wire N__46577;
    wire N__46574;
    wire N__46571;
    wire N__46568;
    wire N__46565;
    wire N__46562;
    wire N__46559;
    wire N__46556;
    wire N__46553;
    wire N__46550;
    wire N__46549;
    wire N__46546;
    wire N__46543;
    wire N__46538;
    wire N__46535;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46511;
    wire N__46508;
    wire N__46505;
    wire N__46502;
    wire N__46501;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46488;
    wire N__46481;
    wire N__46478;
    wire N__46477;
    wire N__46472;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46462;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46433;
    wire N__46430;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46403;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46382;
    wire N__46379;
    wire N__46378;
    wire N__46373;
    wire N__46370;
    wire N__46367;
    wire N__46364;
    wire N__46361;
    wire N__46358;
    wire N__46355;
    wire N__46352;
    wire N__46351;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46339;
    wire N__46334;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46307;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46295;
    wire N__46294;
    wire N__46289;
    wire N__46286;
    wire N__46283;
    wire N__46280;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46238;
    wire N__46237;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46220;
    wire N__46217;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46207;
    wire N__46204;
    wire N__46201;
    wire N__46198;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46147;
    wire N__46144;
    wire N__46139;
    wire N__46136;
    wire N__46133;
    wire N__46130;
    wire N__46127;
    wire N__46124;
    wire N__46121;
    wire N__46118;
    wire N__46117;
    wire N__46114;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46100;
    wire N__46097;
    wire N__46094;
    wire N__46091;
    wire N__46088;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46076;
    wire N__46075;
    wire N__46070;
    wire N__46067;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46055;
    wire N__46052;
    wire N__46049;
    wire N__46046;
    wire N__46043;
    wire N__46040;
    wire N__46039;
    wire N__46036;
    wire N__46033;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45991;
    wire N__45988;
    wire N__45983;
    wire N__45980;
    wire N__45977;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45959;
    wire N__45956;
    wire N__45953;
    wire N__45950;
    wire N__45947;
    wire N__45944;
    wire N__45941;
    wire N__45938;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45887;
    wire N__45884;
    wire N__45881;
    wire N__45878;
    wire N__45875;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45806;
    wire N__45805;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45776;
    wire N__45773;
    wire N__45770;
    wire N__45767;
    wire N__45766;
    wire N__45763;
    wire N__45760;
    wire N__45757;
    wire N__45754;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45740;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45728;
    wire N__45725;
    wire N__45724;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45690;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45673;
    wire N__45670;
    wire N__45667;
    wire N__45662;
    wire N__45659;
    wire N__45658;
    wire N__45655;
    wire N__45652;
    wire N__45649;
    wire N__45646;
    wire N__45641;
    wire N__45638;
    wire N__45635;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45614;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45583;
    wire N__45580;
    wire N__45577;
    wire N__45572;
    wire N__45569;
    wire N__45566;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45516;
    wire N__45515;
    wire N__45510;
    wire N__45509;
    wire N__45506;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45483;
    wire N__45480;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45458;
    wire N__45455;
    wire N__45452;
    wire N__45449;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45421;
    wire N__45410;
    wire N__45407;
    wire N__45404;
    wire N__45403;
    wire N__45402;
    wire N__45401;
    wire N__45398;
    wire N__45393;
    wire N__45392;
    wire N__45391;
    wire N__45390;
    wire N__45387;
    wire N__45382;
    wire N__45375;
    wire N__45368;
    wire N__45365;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45343;
    wire N__45340;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45326;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45316;
    wire N__45313;
    wire N__45310;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45281;
    wire N__45280;
    wire N__45277;
    wire N__45274;
    wire N__45269;
    wire N__45266;
    wire N__45263;
    wire N__45262;
    wire N__45259;
    wire N__45256;
    wire N__45253;
    wire N__45250;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45238;
    wire N__45233;
    wire N__45230;
    wire N__45227;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45188;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45161;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45145;
    wire N__45144;
    wire N__45143;
    wire N__45138;
    wire N__45133;
    wire N__45130;
    wire N__45127;
    wire N__45122;
    wire N__45121;
    wire N__45120;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45098;
    wire N__45095;
    wire N__45092;
    wire N__45089;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45065;
    wire N__45062;
    wire N__45059;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45051;
    wire N__45050;
    wire N__45045;
    wire N__45040;
    wire N__45035;
    wire N__45032;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45020;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45010;
    wire N__45009;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44963;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44945;
    wire N__44942;
    wire N__44939;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44927;
    wire N__44924;
    wire N__44921;
    wire N__44920;
    wire N__44917;
    wire N__44914;
    wire N__44909;
    wire N__44906;
    wire N__44903;
    wire N__44902;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44897;
    wire N__44896;
    wire N__44891;
    wire N__44888;
    wire N__44885;
    wire N__44884;
    wire N__44883;
    wire N__44882;
    wire N__44879;
    wire N__44872;
    wire N__44871;
    wire N__44870;
    wire N__44869;
    wire N__44868;
    wire N__44867;
    wire N__44866;
    wire N__44865;
    wire N__44864;
    wire N__44863;
    wire N__44862;
    wire N__44859;
    wire N__44854;
    wire N__44849;
    wire N__44846;
    wire N__44841;
    wire N__44840;
    wire N__44839;
    wire N__44836;
    wire N__44827;
    wire N__44824;
    wire N__44819;
    wire N__44816;
    wire N__44813;
    wire N__44810;
    wire N__44801;
    wire N__44796;
    wire N__44791;
    wire N__44774;
    wire N__44773;
    wire N__44770;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44759;
    wire N__44756;
    wire N__44753;
    wire N__44750;
    wire N__44749;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44736;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44714;
    wire N__44713;
    wire N__44712;
    wire N__44709;
    wire N__44708;
    wire N__44707;
    wire N__44706;
    wire N__44705;
    wire N__44704;
    wire N__44703;
    wire N__44702;
    wire N__44701;
    wire N__44700;
    wire N__44697;
    wire N__44696;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44680;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44663;
    wire N__44662;
    wire N__44661;
    wire N__44660;
    wire N__44659;
    wire N__44658;
    wire N__44657;
    wire N__44656;
    wire N__44655;
    wire N__44654;
    wire N__44651;
    wire N__44650;
    wire N__44649;
    wire N__44646;
    wire N__44641;
    wire N__44640;
    wire N__44639;
    wire N__44638;
    wire N__44637;
    wire N__44636;
    wire N__44635;
    wire N__44634;
    wire N__44633;
    wire N__44632;
    wire N__44631;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44604;
    wire N__44601;
    wire N__44594;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44565;
    wire N__44560;
    wire N__44549;
    wire N__44546;
    wire N__44541;
    wire N__44530;
    wire N__44523;
    wire N__44498;
    wire N__44497;
    wire N__44496;
    wire N__44495;
    wire N__44490;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44478;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44462;
    wire N__44461;
    wire N__44458;
    wire N__44457;
    wire N__44454;
    wire N__44453;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44435;
    wire N__44434;
    wire N__44429;
    wire N__44426;
    wire N__44419;
    wire N__44416;
    wire N__44415;
    wire N__44412;
    wire N__44407;
    wire N__44402;
    wire N__44399;
    wire N__44398;
    wire N__44397;
    wire N__44396;
    wire N__44393;
    wire N__44390;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44345;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44320;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44308;
    wire N__44307;
    wire N__44304;
    wire N__44299;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44278;
    wire N__44273;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44249;
    wire N__44246;
    wire N__44243;
    wire N__44242;
    wire N__44239;
    wire N__44236;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44195;
    wire N__44192;
    wire N__44189;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44179;
    wire N__44178;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44162;
    wire N__44159;
    wire N__44156;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44101;
    wire N__44098;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44059;
    wire N__44056;
    wire N__44053;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44033;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43999;
    wire N__43998;
    wire N__43997;
    wire N__43992;
    wire N__43987;
    wire N__43984;
    wire N__43983;
    wire N__43982;
    wire N__43981;
    wire N__43980;
    wire N__43979;
    wire N__43976;
    wire N__43975;
    wire N__43974;
    wire N__43971;
    wire N__43964;
    wire N__43959;
    wire N__43956;
    wire N__43951;
    wire N__43948;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43930;
    wire N__43925;
    wire N__43922;
    wire N__43921;
    wire N__43920;
    wire N__43919;
    wire N__43918;
    wire N__43917;
    wire N__43916;
    wire N__43915;
    wire N__43914;
    wire N__43913;
    wire N__43912;
    wire N__43909;
    wire N__43904;
    wire N__43903;
    wire N__43898;
    wire N__43897;
    wire N__43896;
    wire N__43891;
    wire N__43886;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43858;
    wire N__43853;
    wire N__43850;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43826;
    wire N__43823;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43748;
    wire N__43745;
    wire N__43744;
    wire N__43741;
    wire N__43736;
    wire N__43733;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43703;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43679;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43603;
    wire N__43600;
    wire N__43599;
    wire N__43596;
    wire N__43591;
    wire N__43590;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43574;
    wire N__43573;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43535;
    wire N__43532;
    wire N__43531;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43508;
    wire N__43507;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43495;
    wire N__43494;
    wire N__43491;
    wire N__43486;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43386;
    wire N__43383;
    wire N__43380;
    wire N__43377;
    wire N__43374;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43349;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43331;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43309;
    wire N__43308;
    wire N__43307;
    wire N__43306;
    wire N__43305;
    wire N__43304;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43296;
    wire N__43295;
    wire N__43294;
    wire N__43293;
    wire N__43288;
    wire N__43287;
    wire N__43280;
    wire N__43279;
    wire N__43278;
    wire N__43277;
    wire N__43274;
    wire N__43269;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43244;
    wire N__43243;
    wire N__43242;
    wire N__43239;
    wire N__43238;
    wire N__43237;
    wire N__43234;
    wire N__43231;
    wire N__43222;
    wire N__43217;
    wire N__43214;
    wire N__43209;
    wire N__43206;
    wire N__43201;
    wire N__43198;
    wire N__43187;
    wire N__43184;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43169;
    wire N__43166;
    wire N__43165;
    wire N__43164;
    wire N__43161;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43134;
    wire N__43127;
    wire N__43124;
    wire N__43121;
    wire N__43120;
    wire N__43119;
    wire N__43118;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43106;
    wire N__43105;
    wire N__43104;
    wire N__43101;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43086;
    wire N__43075;
    wire N__43072;
    wire N__43067;
    wire N__43066;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43055;
    wire N__43052;
    wire N__43051;
    wire N__43048;
    wire N__43045;
    wire N__43042;
    wire N__43041;
    wire N__43040;
    wire N__43039;
    wire N__43038;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43010;
    wire N__42995;
    wire N__42992;
    wire N__42991;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42983;
    wire N__42982;
    wire N__42979;
    wire N__42978;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42941;
    wire N__42938;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42859;
    wire N__42854;
    wire N__42851;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42811;
    wire N__42810;
    wire N__42807;
    wire N__42802;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42788;
    wire N__42787;
    wire N__42782;
    wire N__42779;
    wire N__42776;
    wire N__42773;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42737;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42719;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42668;
    wire N__42665;
    wire N__42662;
    wire N__42659;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42626;
    wire N__42623;
    wire N__42620;
    wire N__42617;
    wire N__42614;
    wire N__42611;
    wire N__42608;
    wire N__42605;
    wire N__42602;
    wire N__42599;
    wire N__42596;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42584;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42569;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42557;
    wire N__42554;
    wire N__42551;
    wire N__42550;
    wire N__42549;
    wire N__42548;
    wire N__42547;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42536;
    wire N__42533;
    wire N__42530;
    wire N__42529;
    wire N__42526;
    wire N__42523;
    wire N__42520;
    wire N__42517;
    wire N__42514;
    wire N__42509;
    wire N__42506;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42490;
    wire N__42485;
    wire N__42482;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42464;
    wire N__42463;
    wire N__42460;
    wire N__42457;
    wire N__42454;
    wire N__42451;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42437;
    wire N__42434;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42410;
    wire N__42407;
    wire N__42404;
    wire N__42401;
    wire N__42400;
    wire N__42397;
    wire N__42394;
    wire N__42389;
    wire N__42386;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42370;
    wire N__42367;
    wire N__42364;
    wire N__42359;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42344;
    wire N__42341;
    wire N__42338;
    wire N__42335;
    wire N__42334;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42322;
    wire N__42319;
    wire N__42316;
    wire N__42313;
    wire N__42310;
    wire N__42305;
    wire N__42304;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42280;
    wire N__42277;
    wire N__42274;
    wire N__42271;
    wire N__42266;
    wire N__42265;
    wire N__42264;
    wire N__42263;
    wire N__42262;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42245;
    wire N__42244;
    wire N__42241;
    wire N__42236;
    wire N__42235;
    wire N__42232;
    wire N__42225;
    wire N__42222;
    wire N__42221;
    wire N__42220;
    wire N__42217;
    wire N__42216;
    wire N__42213;
    wire N__42212;
    wire N__42209;
    wire N__42208;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42196;
    wire N__42195;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42176;
    wire N__42169;
    wire N__42162;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42110;
    wire N__42107;
    wire N__42104;
    wire N__42101;
    wire N__42098;
    wire N__42095;
    wire N__42092;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42082;
    wire N__42081;
    wire N__42080;
    wire N__42077;
    wire N__42074;
    wire N__42071;
    wire N__42070;
    wire N__42067;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42049;
    wire N__42044;
    wire N__42041;
    wire N__42038;
    wire N__42035;
    wire N__42032;
    wire N__42029;
    wire N__42026;
    wire N__42023;
    wire N__42020;
    wire N__42017;
    wire N__42014;
    wire N__42011;
    wire N__42008;
    wire N__42005;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41986;
    wire N__41983;
    wire N__41982;
    wire N__41981;
    wire N__41978;
    wire N__41977;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41960;
    wire N__41959;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41941;
    wire N__41938;
    wire N__41933;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41923;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41888;
    wire N__41885;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41870;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41846;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41824;
    wire N__41819;
    wire N__41816;
    wire N__41813;
    wire N__41810;
    wire N__41807;
    wire N__41806;
    wire N__41805;
    wire N__41802;
    wire N__41797;
    wire N__41792;
    wire N__41789;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41764;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41747;
    wire N__41744;
    wire N__41741;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41729;
    wire N__41726;
    wire N__41723;
    wire N__41720;
    wire N__41717;
    wire N__41716;
    wire N__41713;
    wire N__41710;
    wire N__41705;
    wire N__41702;
    wire N__41699;
    wire N__41698;
    wire N__41697;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41689;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41671;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41659;
    wire N__41656;
    wire N__41655;
    wire N__41652;
    wire N__41651;
    wire N__41650;
    wire N__41647;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41628;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41602;
    wire N__41597;
    wire N__41596;
    wire N__41595;
    wire N__41594;
    wire N__41591;
    wire N__41586;
    wire N__41583;
    wire N__41582;
    wire N__41581;
    wire N__41580;
    wire N__41577;
    wire N__41576;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41563;
    wire N__41560;
    wire N__41559;
    wire N__41558;
    wire N__41555;
    wire N__41550;
    wire N__41545;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41531;
    wire N__41526;
    wire N__41523;
    wire N__41518;
    wire N__41515;
    wire N__41504;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41489;
    wire N__41488;
    wire N__41485;
    wire N__41480;
    wire N__41477;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41465;
    wire N__41464;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41435;
    wire N__41434;
    wire N__41433;
    wire N__41432;
    wire N__41431;
    wire N__41430;
    wire N__41429;
    wire N__41428;
    wire N__41425;
    wire N__41424;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41416;
    wire N__41415;
    wire N__41412;
    wire N__41409;
    wire N__41408;
    wire N__41405;
    wire N__41398;
    wire N__41397;
    wire N__41396;
    wire N__41395;
    wire N__41394;
    wire N__41393;
    wire N__41392;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41372;
    wire N__41371;
    wire N__41366;
    wire N__41363;
    wire N__41358;
    wire N__41357;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41340;
    wire N__41337;
    wire N__41328;
    wire N__41319;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41289;
    wire N__41284;
    wire N__41277;
    wire N__41264;
    wire N__41261;
    wire N__41260;
    wire N__41259;
    wire N__41258;
    wire N__41257;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41249;
    wire N__41248;
    wire N__41247;
    wire N__41246;
    wire N__41245;
    wire N__41242;
    wire N__41241;
    wire N__41236;
    wire N__41235;
    wire N__41234;
    wire N__41233;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41211;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41203;
    wire N__41202;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41194;
    wire N__41193;
    wire N__41192;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41163;
    wire N__41158;
    wire N__41155;
    wire N__41146;
    wire N__41137;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41101;
    wire N__41100;
    wire N__41097;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41054;
    wire N__41053;
    wire N__41052;
    wire N__41051;
    wire N__41046;
    wire N__41041;
    wire N__41036;
    wire N__41033;
    wire N__41030;
    wire N__41027;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40999;
    wire N__40996;
    wire N__40993;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40963;
    wire N__40962;
    wire N__40959;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40940;
    wire N__40935;
    wire N__40930;
    wire N__40925;
    wire N__40924;
    wire N__40921;
    wire N__40920;
    wire N__40917;
    wire N__40916;
    wire N__40915;
    wire N__40914;
    wire N__40913;
    wire N__40912;
    wire N__40911;
    wire N__40906;
    wire N__40901;
    wire N__40896;
    wire N__40893;
    wire N__40892;
    wire N__40891;
    wire N__40890;
    wire N__40889;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40839;
    wire N__40832;
    wire N__40829;
    wire N__40826;
    wire N__40823;
    wire N__40820;
    wire N__40819;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40802;
    wire N__40801;
    wire N__40800;
    wire N__40797;
    wire N__40796;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40762;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40750;
    wire N__40749;
    wire N__40746;
    wire N__40741;
    wire N__40736;
    wire N__40733;
    wire N__40730;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40715;
    wire N__40712;
    wire N__40709;
    wire N__40706;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40688;
    wire N__40685;
    wire N__40682;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40637;
    wire N__40636;
    wire N__40629;
    wire N__40626;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40601;
    wire N__40598;
    wire N__40595;
    wire N__40594;
    wire N__40593;
    wire N__40592;
    wire N__40589;
    wire N__40586;
    wire N__40585;
    wire N__40582;
    wire N__40581;
    wire N__40580;
    wire N__40577;
    wire N__40576;
    wire N__40571;
    wire N__40568;
    wire N__40565;
    wire N__40560;
    wire N__40555;
    wire N__40550;
    wire N__40541;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40504;
    wire N__40499;
    wire N__40498;
    wire N__40495;
    wire N__40494;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40357;
    wire N__40354;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40325;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40298;
    wire N__40297;
    wire N__40296;
    wire N__40293;
    wire N__40292;
    wire N__40287;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40268;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40227;
    wire N__40220;
    wire N__40219;
    wire N__40216;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40204;
    wire N__40201;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40134;
    wire N__40131;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40108;
    wire N__40105;
    wire N__40102;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40090;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40073;
    wire N__40070;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39998;
    wire N__39995;
    wire N__39992;
    wire N__39989;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39973;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39949;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39923;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39913;
    wire N__39910;
    wire N__39905;
    wire N__39902;
    wire N__39899;
    wire N__39896;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39874;
    wire N__39871;
    wire N__39866;
    wire N__39863;
    wire N__39862;
    wire N__39859;
    wire N__39856;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39841;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39715;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39652;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39607;
    wire N__39606;
    wire N__39605;
    wire N__39604;
    wire N__39603;
    wire N__39600;
    wire N__39599;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39558;
    wire N__39551;
    wire N__39544;
    wire N__39539;
    wire N__39536;
    wire N__39535;
    wire N__39532;
    wire N__39531;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39517;
    wire N__39516;
    wire N__39515;
    wire N__39514;
    wire N__39511;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39479;
    wire N__39476;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39458;
    wire N__39457;
    wire N__39456;
    wire N__39455;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39394;
    wire N__39393;
    wire N__39392;
    wire N__39391;
    wire N__39388;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39335;
    wire N__39330;
    wire N__39323;
    wire N__39322;
    wire N__39321;
    wire N__39320;
    wire N__39319;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39302;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39265;
    wire N__39260;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39233;
    wire N__39230;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39218;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39194;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39100;
    wire N__39097;
    wire N__39096;
    wire N__39095;
    wire N__39092;
    wire N__39091;
    wire N__39090;
    wire N__39089;
    wire N__39088;
    wire N__39087;
    wire N__39086;
    wire N__39083;
    wire N__39078;
    wire N__39075;
    wire N__39068;
    wire N__39061;
    wire N__39058;
    wire N__39047;
    wire N__39046;
    wire N__39045;
    wire N__39044;
    wire N__39041;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39027;
    wire N__39026;
    wire N__39025;
    wire N__39024;
    wire N__39023;
    wire N__39020;
    wire N__39013;
    wire N__39010;
    wire N__39005;
    wire N__38998;
    wire N__38993;
    wire N__38990;
    wire N__38981;
    wire N__38978;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38939;
    wire N__38936;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38869;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38848;
    wire N__38847;
    wire N__38844;
    wire N__38839;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38821;
    wire N__38818;
    wire N__38815;
    wire N__38810;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38800;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38765;
    wire N__38764;
    wire N__38761;
    wire N__38758;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38723;
    wire N__38720;
    wire N__38717;
    wire N__38716;
    wire N__38715;
    wire N__38714;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38700;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38679;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38648;
    wire N__38645;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38596;
    wire N__38595;
    wire N__38588;
    wire N__38585;
    wire N__38584;
    wire N__38583;
    wire N__38582;
    wire N__38581;
    wire N__38580;
    wire N__38579;
    wire N__38576;
    wire N__38571;
    wire N__38568;
    wire N__38567;
    wire N__38566;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38545;
    wire N__38542;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38444;
    wire N__38443;
    wire N__38442;
    wire N__38441;
    wire N__38438;
    wire N__38437;
    wire N__38432;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38415;
    wire N__38412;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38384;
    wire N__38375;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38336;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38265;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38253;
    wire N__38250;
    wire N__38249;
    wire N__38248;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38231;
    wire N__38226;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38210;
    wire N__38209;
    wire N__38206;
    wire N__38205;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38193;
    wire N__38186;
    wire N__38185;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38144;
    wire N__38141;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38127;
    wire N__38126;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38105;
    wire N__38102;
    wire N__38093;
    wire N__38090;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38066;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38058;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38032;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38006;
    wire N__38003;
    wire N__38000;
    wire N__37997;
    wire N__37994;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37981;
    wire N__37978;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37964;
    wire N__37961;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37874;
    wire N__37871;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37802;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37769;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37745;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37702;
    wire N__37699;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37684;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37663;
    wire N__37660;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37645;
    wire N__37642;
    wire N__37637;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37580;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37565;
    wire N__37562;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37549;
    wire N__37548;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37532;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37520;
    wire N__37517;
    wire N__37516;
    wire N__37513;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37495;
    wire N__37492;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37438;
    wire N__37435;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37358;
    wire N__37355;
    wire N__37354;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37342;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37318;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37285;
    wire N__37282;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37261;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37113;
    wire N__37112;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36949;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36918;
    wire N__36915;
    wire N__36910;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36883;
    wire N__36880;
    wire N__36879;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36841;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36817;
    wire N__36814;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36688;
    wire N__36685;
    wire N__36684;
    wire N__36681;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36663;
    wire N__36658;
    wire N__36655;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36625;
    wire N__36622;
    wire N__36621;
    wire N__36618;
    wire N__36613;
    wire N__36610;
    wire N__36609;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36448;
    wire N__36447;
    wire N__36444;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36433;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36370;
    wire N__36365;
    wire N__36364;
    wire N__36363;
    wire N__36362;
    wire N__36361;
    wire N__36358;
    wire N__36353;
    wire N__36348;
    wire N__36341;
    wire N__36340;
    wire N__36339;
    wire N__36338;
    wire N__36333;
    wire N__36328;
    wire N__36327;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36319;
    wire N__36318;
    wire N__36317;
    wire N__36316;
    wire N__36315;
    wire N__36310;
    wire N__36305;
    wire N__36302;
    wire N__36297;
    wire N__36292;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36241;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36206;
    wire N__36205;
    wire N__36200;
    wire N__36197;
    wire N__36196;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36103;
    wire N__36100;
    wire N__36097;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36035;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36008;
    wire N__36005;
    wire N__36004;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35980;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35968;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35930;
    wire N__35929;
    wire N__35928;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35873;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35837;
    wire N__35834;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35798;
    wire N__35797;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35784;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35768;
    wire N__35765;
    wire N__35764;
    wire N__35761;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35731;
    wire N__35728;
    wire N__35723;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35636;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35550;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35222;
    wire N__35219;
    wire N__35216;
    wire N__35213;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35135;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35113;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35102;
    wire N__35101;
    wire N__35100;
    wire N__35099;
    wire N__35098;
    wire N__35097;
    wire N__35090;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35071;
    wire N__35056;
    wire N__35053;
    wire N__35052;
    wire N__35051;
    wire N__35050;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35027;
    wire N__35026;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35008;
    wire N__35007;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34991;
    wire N__34990;
    wire N__34989;
    wire N__34986;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34970;
    wire N__34967;
    wire N__34966;
    wire N__34965;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34954;
    wire N__34951;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34816;
    wire N__34811;
    wire N__34808;
    wire N__34807;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34771;
    wire N__34770;
    wire N__34769;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34757;
    wire N__34754;
    wire N__34753;
    wire N__34750;
    wire N__34743;
    wire N__34740;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34645;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34567;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34553;
    wire N__34548;
    wire N__34543;
    wire N__34542;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34518;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34460;
    wire N__34457;
    wire N__34456;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34432;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34414;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34310;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34243;
    wire N__34242;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34142;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34099;
    wire N__34096;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34083;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34067;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34013;
    wire N__34012;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33997;
    wire N__33994;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33721;
    wire N__33718;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33343;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33306;
    wire N__33301;
    wire N__33298;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33236;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33143;
    wire N__33140;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33058;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33032;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32983;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32938;
    wire N__32937;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32845;
    wire N__32842;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32828;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32816;
    wire N__32811;
    wire N__32810;
    wire N__32809;
    wire N__32806;
    wire N__32801;
    wire N__32796;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32776;
    wire N__32771;
    wire N__32768;
    wire N__32767;
    wire N__32762;
    wire N__32759;
    wire N__32758;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32728;
    wire N__32725;
    wire N__32722;
    wire N__32719;
    wire N__32716;
    wire N__32713;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32689;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32578;
    wire N__32573;
    wire N__32570;
    wire N__32569;
    wire N__32568;
    wire N__32567;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32559;
    wire N__32558;
    wire N__32555;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32544;
    wire N__32531;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32514;
    wire N__32513;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32495;
    wire N__32494;
    wire N__32493;
    wire N__32486;
    wire N__32483;
    wire N__32482;
    wire N__32481;
    wire N__32480;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32468;
    wire N__32465;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32457;
    wire N__32456;
    wire N__32453;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32429;
    wire N__32424;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32392;
    wire N__32389;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32347;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32323;
    wire N__32322;
    wire N__32321;
    wire N__32320;
    wire N__32319;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32308;
    wire N__32307;
    wire N__32304;
    wire N__32303;
    wire N__32302;
    wire N__32301;
    wire N__32300;
    wire N__32299;
    wire N__32296;
    wire N__32295;
    wire N__32290;
    wire N__32287;
    wire N__32282;
    wire N__32277;
    wire N__32274;
    wire N__32265;
    wire N__32264;
    wire N__32263;
    wire N__32262;
    wire N__32261;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32247;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32232;
    wire N__32221;
    wire N__32212;
    wire N__32207;
    wire N__32200;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32012;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31756;
    wire N__31755;
    wire N__31752;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31714;
    wire N__31711;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31277;
    wire N__31276;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31246;
    wire N__31243;
    wire N__31238;
    wire N__31235;
    wire N__31234;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31207;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31169;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31156;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31112;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31085;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30994;
    wire N__30993;
    wire N__30992;
    wire N__30989;
    wire N__30984;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30880;
    wire N__30879;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30793;
    wire N__30792;
    wire N__30791;
    wire N__30790;
    wire N__30789;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30773;
    wire N__30770;
    wire N__30761;
    wire N__30760;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30739;
    wire N__30736;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30542;
    wire N__30541;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30497;
    wire N__30494;
    wire N__30491;
    wire N__30490;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30350;
    wire N__30347;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29842;
    wire N__29839;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29825;
    wire N__29824;
    wire N__29823;
    wire N__29822;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29808;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29726;
    wire N__29723;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29708;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29700;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29456;
    wire N__29455;
    wire N__29452;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29425;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29398;
    wire N__29395;
    wire N__29392;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29173;
    wire N__29170;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29140;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28961;
    wire N__28958;
    wire N__28955;
    wire N__28952;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28922;
    wire N__28921;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28877;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28697;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28537;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28520;
    wire N__28519;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28441;
    wire N__28440;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28123;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28112;
    wire N__28111;
    wire N__28110;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28086;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28013;
    wire N__28012;
    wire N__28007;
    wire N__28004;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27989;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27955;
    wire N__27954;
    wire N__27953;
    wire N__27950;
    wire N__27943;
    wire N__27938;
    wire N__27937;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27922;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27898;
    wire N__27897;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27885;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27754;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27499;
    wire N__27498;
    wire N__27495;
    wire N__27494;
    wire N__27493;
    wire N__27488;
    wire N__27485;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27467;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27286;
    wire N__27285;
    wire N__27284;
    wire N__27283;
    wire N__27278;
    wire N__27271;
    wire N__27270;
    wire N__27269;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27255;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27194;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27179;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27104;
    wire N__27101;
    wire N__27100;
    wire N__27099;
    wire N__27092;
    wire N__27089;
    wire N__27088;
    wire N__27087;
    wire N__27084;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27019;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26932;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26752;
    wire N__26751;
    wire N__26750;
    wire N__26747;
    wire N__26744;
    wire N__26737;
    wire N__26734;
    wire N__26729;
    wire N__26726;
    wire N__26725;
    wire N__26724;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26146;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26108;
    wire N__26107;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25793;
    wire N__25792;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25673;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire \INVCONTROL.addrstack_addrstack_0_0RCLKN_net ;
    wire \INVDROM.ROMDATA.dintern_0_3RCLKN_net ;
    wire \INVDROM.ROMDATA.dintern_0_2RCLKN_net ;
    wire \INVDROM.ROMDATA.dintern_0_1RCLKN_net ;
    wire VCCG0;
    wire \INVDROM.ROMDATA.dintern_0_0RCLKN_net ;
    wire GNDG0;
    wire clkdivZ0Z_0;
    wire bfn_1_17_0_;
    wire clkdivZ0Z_1;
    wire clkdiv_cry_0;
    wire clkdivZ0Z_2;
    wire clkdiv_cry_1;
    wire clkdivZ0Z_3;
    wire clkdiv_cry_2;
    wire clkdivZ0Z_4;
    wire clkdiv_cry_3;
    wire clkdivZ0Z_5;
    wire clkdiv_cry_4;
    wire clkdivZ0Z_6;
    wire clkdiv_cry_5;
    wire clkdivZ0Z_7;
    wire clkdiv_cry_6;
    wire clkdiv_cry_7;
    wire clkdivZ0Z_8;
    wire bfn_1_18_0_;
    wire clkdivZ0Z_9;
    wire clkdiv_cry_8;
    wire clkdivZ0Z_10;
    wire clkdiv_cry_9;
    wire clkdivZ0Z_11;
    wire clkdiv_cry_10;
    wire clkdivZ0Z_12;
    wire clkdiv_cry_11;
    wire clkdivZ0Z_13;
    wire clkdiv_cry_12;
    wire clkdivZ0Z_14;
    wire clkdiv_cry_13;
    wire clkdivZ0Z_15;
    wire clkdiv_cry_14;
    wire clkdiv_cry_15;
    wire clkdivZ0Z_16;
    wire bfn_1_19_0_;
    wire clkdivZ0Z_17;
    wire clkdiv_cry_16;
    wire clkdivZ0Z_18;
    wire clkdiv_cry_17;
    wire clkdivZ0Z_19;
    wire clkdiv_cry_18;
    wire clkdivZ0Z_20;
    wire clkdiv_cry_19;
    wire clkdivZ0Z_21;
    wire clkdiv_cry_20;
    wire clkdivZ0Z_22;
    wire clkdiv_cry_21;
    wire clkdiv_cry_22;
    wire GPIO3_c;
    wire B_OE_c_i;
    wire B_OE_c;
    wire gpuAddress_11;
    wire \INVCONTROL.gpuAddReg_11C_net ;
    wire gpuAddress_14;
    wire \INVCONTROL.gpuAddReg_14C_net ;
    wire gpuAddress_9;
    wire \INVCONTROL.gpuAddReg_9C_net ;
    wire N_6_0;
    wire RAM_un1_WR_i;
    wire bfn_9_9_0_;
    wire \ALU.status_17_data_tmp_0 ;
    wire \ALU.status_17_data_tmp_1 ;
    wire \ALU.status_17_data_tmp_2 ;
    wire \ALU.status_17_data_tmp_3 ;
    wire \ALU.status_17_data_tmp_4 ;
    wire \ALU.status_17_data_tmp_5 ;
    wire \ALU.status_17_data_tmp_6 ;
    wire \ALU.status_17_data_tmp_7 ;
    wire bfn_9_10_0_;
    wire \ALU.status_17_I_45_c_RNOZ0 ;
    wire bfn_9_11_0_;
    wire \ALU.combOperand2_i_1 ;
    wire \ALU.status_18_cry_0 ;
    wire \ALU.status_18_cry_1 ;
    wire \ALU.status_18_cry_2 ;
    wire \ALU.status_18_cry_3 ;
    wire \ALU.status_18_cry_4 ;
    wire \ALU.status_17_I_27_c_RNOZ0 ;
    wire \ALU.status_18_cry_5 ;
    wire \ALU.combOperand2_i_7 ;
    wire \ALU.status_18_cry_6 ;
    wire \ALU.status_18_cry_7 ;
    wire bfn_9_12_0_;
    wire \ALU.status_18_cry_8 ;
    wire \ALU.status_18_cry_9 ;
    wire \ALU.combOperand2_i_11 ;
    wire \ALU.status_18_cry_10 ;
    wire \ALU.status_18_cry_11 ;
    wire \ALU.status_18_cry_12 ;
    wire \ALU.combOperand2_i_14 ;
    wire \ALU.status_18_cry_13 ;
    wire \ALU.combOperand2_i_15 ;
    wire \ALU.status_18_cry_14 ;
    wire \ALU.status_18_4 ;
    wire bfn_9_13_0_;
    wire \ALU.status_18_cry_10_c_RNOZ0 ;
    wire \ALU.status_18_cry_13_c_RNOZ0 ;
    wire \CONTROL.busState_1_RNIG7366Z0Z_2_cascade_ ;
    wire \CONTROL.busState_1_RNI1JVK1_0Z0Z_2 ;
    wire gpuOut_c_5;
    wire \CONTROL.N_166 ;
    wire D5_in_c;
    wire \CONTROL.N_166_cascade_ ;
    wire romOut_5;
    wire \INVCONTROL.dout_5C_net ;
    wire \ALU.operand2_12_cascade_ ;
    wire \ALU.N_126_cascade_ ;
    wire \ALU.c_RNI670LZ0Z_12_cascade_ ;
    wire \ALU.operand2_7_ns_1_12 ;
    wire \ALU.d_RNI8FCTZ0Z_12 ;
    wire \ALU.operand2_12 ;
    wire \ALU.status_18_cry_12_c_RNOZ0 ;
    wire \ALU.log_1_3cf0_1_10 ;
    wire \ALU.log_1_3cf0_10_cascade_ ;
    wire \ALU.log_1_3cf1_10 ;
    wire \ALU.log_1_3cf1_1_10 ;
    wire \CONTROL.bus_7_a0_2_8_cascade_ ;
    wire \ALU.status_18_cry_8_c_RNOZ0 ;
    wire DROM_ROMDATA_dintern_8ro_cascade_;
    wire DROM_ROMDATA_dintern_8ro;
    wire bus_8;
    wire \DROM.ROMDATA.dintern_0_0_NEW_1 ;
    wire \DROM.ROMDATA.dintern_0_0_OLDZ0Z_1 ;
    wire \INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C_net ;
    wire \DROM.ROMDATA.dintern_0_2_NEW_0 ;
    wire \DROM.ROMDATA.dintern_0_2_OLDZ0Z_0 ;
    wire \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net ;
    wire DROM_ROMDATA_dintern_12ro_cascade_;
    wire \INVCONTROL.aluOperation_3C_net ;
    wire DROM_ROMDATA_dintern_12ro;
    wire bus_12;
    wire \DROM.ROMDATA.dintern_0_3_OLDZ0Z_2 ;
    wire \DROM.ROMDATA.dintern_0_3_NEW_2 ;
    wire \DROM.ROMDATA.dintern_0_3_OLDZ0Z_3 ;
    wire \DROM.ROMDATA.dintern_0_3_NEW_3 ;
    wire bus_10;
    wire gpuAddress_0;
    wire gpuAddress_1;
    wire gpuAddress_10;
    wire gpuAddress_12;
    wire gpuAddress_13;
    wire gpuAddress_15;
    wire \INVCONTROL.gpuAddReg_0C_net ;
    wire CONTROL_romAddReg_7_2;
    wire CONTROL_romAddReg_7_3;
    wire \INVCONTROL.dout_3C_net ;
    wire CONTROL_romAddReg_7_5;
    wire PROM_ROMDATA_dintern_23ro_cascade_;
    wire CONTROL_romAddReg_7_7;
    wire CONTROL_romAddReg_7_6;
    wire \PROM.ROMDATA.m465_bm_cascade_ ;
    wire \PROM.ROMDATA.m471_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m471_ns_cascade_ ;
    wire controlWord_24_cascade_;
    wire CONTROL_romAddReg_7_8;
    wire CONTROL_romAddReg_7_4;
    wire \CONTROL.g0_3_cascade_ ;
    wire \CONTROL.addrstackptr_N_10_mux_0_0_0_cascade_ ;
    wire \CONTROL.addrstackptr_N_7_0_i ;
    wire \CONTROL.N_6_1_cascade_ ;
    wire \CONTROL.N_4_2 ;
    wire \CONTROL.N_4_2_cascade_ ;
    wire \CONTROL.addrstackptr_N_10_mux_0_0_0 ;
    wire \INVCONTROL.addrstackptr_6C_net ;
    wire \CONTROL.tempCounterZ0Z_13 ;
    wire \CONTROL.tempCounterZ0Z_6 ;
    wire \INVCONTROL.tempCounter_13C_net ;
    wire bfn_9_25_0_;
    wire \CONTROL.addrstack_1_cry_0 ;
    wire \CONTROL.addrstack_1_cry_1 ;
    wire \CONTROL.addrstack_1_cry_2 ;
    wire \CONTROL.addrstack_1_cry_3 ;
    wire \CONTROL.addrstack_1_cry_4 ;
    wire \CONTROL.addrstackptrZ0Z_6 ;
    wire \CONTROL.addrstack_1_6 ;
    wire \CONTROL.addrstack_1_cry_5 ;
    wire \CONTROL.addrstack_1_cry_6 ;
    wire \ALU.dout_3_ns_1_5_cascade_ ;
    wire \ALU.dout_6_ns_1_5_cascade_ ;
    wire \ALU.N_1138_cascade_ ;
    wire \ALU.N_1090 ;
    wire aluOut_5_cascade_;
    wire \ALU.status_19_4_cascade_ ;
    wire \ALU.status_17_I_15_c_RNOZ0 ;
    wire \ALU.combOperand2_0_6 ;
    wire \ALU.combOperand2_0_6_cascade_ ;
    wire \ALU.status_19_5_cascade_ ;
    wire \ALU.combOperand2_0_4_cascade_ ;
    wire N_181_cascade_;
    wire \ALU.d_RNIVKK66Z0Z_4 ;
    wire \ALU.d_RNIVKK66Z0Z_4_cascade_ ;
    wire \ALU.combOperand2_0_4 ;
    wire \ALU.status_17_I_33_c_RNOZ0 ;
    wire N_182;
    wire \ALU.combOperand2_0_0_6 ;
    wire \ALU.b_RNI4VJC1Z0Z_12 ;
    wire \ALU.d_RNI4BCTZ0Z_10 ;
    wire \ALU.b_RNI0RJC1Z0Z_10_cascade_ ;
    wire \ALU.operand2_10 ;
    wire \ALU.operand2_10_cascade_ ;
    wire \ALU.status_19_9_cascade_ ;
    wire \ALU.e_RNIBHMNZ0Z_8_cascade_ ;
    wire \ALU.d_RNIIINJZ0Z_8 ;
    wire \ALU.operand2_7_ns_1_8 ;
    wire \ALU.b_RNIE6BVZ0Z_8_cascade_ ;
    wire \ALU.operand2_8 ;
    wire busState_1_RNI05PC2_0;
    wire \ALU.operand2_8_cascade_ ;
    wire \ALU.status_18_cry_3_c_RNOZ0 ;
    wire N_228_0_cascade_;
    wire \INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C_net ;
    wire \DROM.ROMDATA.dintern_0_0_OLDZ0Z_3 ;
    wire \DROM.ROMDATA.dintern_0_0_NEW_3 ;
    wire DROM_ROMDATA_dintern_3ro_cascade_;
    wire DROM_ROMDATA_dintern_1ro;
    wire DROM_ROMDATA_dintern_adflt_cascade_;
    wire \DROM.ROMDATA.dintern_adfltZ0Z_3 ;
    wire \DROM.ROMDATA.dintern_adfltZ0Z_3_cascade_ ;
    wire \DROM.ROMDATA.dintern_adflt_sxZ0 ;
    wire dataRomAddress_13;
    wire dataRomAddress_14;
    wire dataRomAddress_15;
    wire \INVCONTROL.romAddReg_13C_net ;
    wire \INVCONTROL.aluOperation_ne_0C_net ;
    wire \DROM.ROMDATA.dintern_0_3_OLDZ0Z_1 ;
    wire \DROM.ROMDATA.dintern_0_3_NEW_1 ;
    wire DROM_ROMDATA_dintern_13ro_cascade_;
    wire \CONTROL.bus_7_a0_2_8 ;
    wire DROM_ROMDATA_dintern_13ro;
    wire bus_13;
    wire DROM_ROMDATA_dintern_10ro;
    wire \DROM.ROMDATA.dintern_0_1_NEW_1 ;
    wire \DROM.ROMDATA.dintern_0_1_OLDZ0Z_1 ;
    wire \DROM.ROMDATA.dintern_0_1_NEW_2 ;
    wire \DROM.ROMDATA.dintern_0_1_OLDZ0Z_2 ;
    wire \DROM.ROMDATA.dintern_0_2_NEW_1 ;
    wire \DROM.ROMDATA.dintern_0_2_OLDZ0Z_1 ;
    wire \DROM.ROMDATA.dintern_0_2_NEW_2 ;
    wire \DROM.ROMDATA.dintern_0_2_OLDZ0Z_2 ;
    wire \DROM.ROMDATA.dintern_0_2_NEW_3 ;
    wire \DROM.ROMDATA.dintern_0_2_OLDZ0Z_3 ;
    wire \DROM.ROMDATA.dintern_0_3_NEW_0 ;
    wire \DROM.ROMDATA.dintern_0_3_OLDZ0Z_0 ;
    wire \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ;
    wire DROM_ROMDATA_dintern_6ro;
    wire \CONTROL.N_199_cascade_ ;
    wire gpuOut_c_6;
    wire D6_in_c;
    wire \CONTROL.N_167_cascade_ ;
    wire N_183;
    wire \INVCONTROL.dout_6C_net ;
    wire \CONTROL.addrstackptr_N_8_mux_1_0_cascade_ ;
    wire \CONTROL.addrstackptr_N_6_0_1_i ;
    wire \CONTROL.g0_3_i_2_cascade_ ;
    wire \CONTROL.N_4_0 ;
    wire \CONTROL.addrstack_1_5 ;
    wire \CONTROL.N_4_0_cascade_ ;
    wire \CONTROL.addrstackptr_N_8_mux_1_0 ;
    wire \CONTROL.addrstackptrZ0Z_5 ;
    wire \INVCONTROL.addrstackptr_5C_net ;
    wire \CONTROL.g0_3_iZ0Z_1 ;
    wire \CONTROL.g0_3_i_a7Z0Z_2 ;
    wire \CONTROL.g0_0_2 ;
    wire \CONTROL.addrstack_12 ;
    wire \CONTROL.addrstack_11 ;
    wire \CONTROL.addrstack_7 ;
    wire \CONTROL.addrstack_14 ;
    wire \CONTROL.tempCounterZ0Z_11 ;
    wire \CONTROL.tempCounterZ0Z_15 ;
    wire \CONTROL.tempCounterZ0Z_14 ;
    wire \INVCONTROL.tempCounter_11C_net ;
    wire \CONTROL.addrstack_8 ;
    wire \CONTROL.addrstack_9 ;
    wire \ALU.status_17_I_9_c_RNOZ0 ;
    wire \ALU.addsub_cry_3_c_RNIGCKVJZ0Z5_cascade_ ;
    wire \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9_cascade_ ;
    wire \ALU.e_RNI26JMZ0Z_4_cascade_ ;
    wire \ALU.operand2_7_ns_1_4_cascade_ ;
    wire \ALU.operand2_4 ;
    wire \ALU.c_RNI6IVQZ0Z_4 ;
    wire \ALU.dout_6_ns_1_4_cascade_ ;
    wire \ALU.aZ0Z_4 ;
    wire \ALU.dout_3_ns_1_4_cascade_ ;
    wire \ALU.N_1089_cascade_ ;
    wire \ALU.N_1137 ;
    wire aluOut_4_cascade_;
    wire \ALU.d_RNIBJM75Z0Z_4 ;
    wire \ALU.status_19_8_cascade_ ;
    wire \ALU.operand2_7_ns_1_6_cascade_ ;
    wire \ALU.operand2_6 ;
    wire \ALU.b_RNI9JSPZ0Z_6 ;
    wire \ALU.e_RNI6AJMZ0Z_6 ;
    wire \ALU.c_RNIAMVQZ0Z_6 ;
    wire \ALU.d_RNIDV8EZ0Z_6 ;
    wire \ALU.c_RNI230LZ0Z_10 ;
    wire \ALU.a_RNIUI741Z0Z_10_cascade_ ;
    wire \ALU.operand2_7_ns_1_10 ;
    wire \ALU.dout_6_ns_1_8_cascade_ ;
    wire ALU_N_1141_cascade_;
    wire \CONTROL.bus_0_sx_8_cascade_ ;
    wire CONTROL_bus_0_8;
    wire \ALU.dout_3_ns_1_8_cascade_ ;
    wire \ALU.c_RNIFT2SZ0Z_8 ;
    wire dataRomAddress_10;
    wire dataRomAddress_12;
    wire \PROM.ROMDATA.dintern_adfltZ0Z_4_cascade_ ;
    wire \PROM.ROMDATA.dintern_12dflt_0Z0Z_1_cascade_ ;
    wire \PROM.ROMDATA.dintern_adfltZ0Z_4 ;
    wire dataRomAddress_11;
    wire \INVCONTROL.romAddReg_10C_net ;
    wire \CONTROL.busState_1_e_1_0_cascade_ ;
    wire \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0_cascade_ ;
    wire N_29;
    wire \CONTROL.N_352 ;
    wire \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0 ;
    wire \INVCONTROL.busState_1_0C_net ;
    wire \DROM.ROMDATA.dintern_0_1_OLDZ0Z_3 ;
    wire \DROM.ROMDATA.dintern_0_1_NEW_3 ;
    wire \DROM.ROMDATA.dintern_0_1_OLDZ0Z_0 ;
    wire \DROM.ROMDATA.dintern_0_1_NEW_0 ;
    wire DROM_ROMDATA_dintern_4ro;
    wire controlWord_29;
    wire controlWord_29_cascade_;
    wire controlWord_28;
    wire controlWord_28_cascade_;
    wire \INVCONTROL.ramAddReg_13C_net ;
    wire A12_c;
    wire A13_c;
    wire \RAM.un1_WR_105_0Z0Z_10 ;
    wire bfn_11_21_0_;
    wire \CONTROL.programCounter_1_cry_0 ;
    wire \CONTROL.programCounter_1_cry_1 ;
    wire \CONTROL.programCounter_1_axb_3 ;
    wire \CONTROL.programCounter_1_cry_2 ;
    wire \CONTROL.programCounter_1_cry_3 ;
    wire \CONTROL.programCounter_1_cry_4 ;
    wire \CONTROL.programCounter_1_cry_5 ;
    wire \CONTROL.programCounter_1_cry_6 ;
    wire \CONTROL.programCounter_1_cry_7 ;
    wire bfn_11_22_0_;
    wire \CONTROL.programCounter_1_cry_8 ;
    wire \CONTROL.programCounter_1_cry_9 ;
    wire \CONTROL.programCounter_1_cry_10 ;
    wire \CONTROL.programCounter_1_cry_11 ;
    wire \CONTROL.programCounter_1_cry_12 ;
    wire \CONTROL.programCounter_1_cry_13 ;
    wire \CONTROL.programCounter_1_cry_14 ;
    wire \CONTROL.programCounter_1_13 ;
    wire \CONTROL.programCounter_1_reto_13 ;
    wire \CONTROL.dout_reto_13 ;
    wire \CONTROL.N_428_cascade_ ;
    wire progRomAddress_13;
    wire \CONTROL.addrstack_reto_14 ;
    wire progRomAddress_14;
    wire \CONTROL.addrstack_13 ;
    wire \CONTROL.addrstack_reto_13 ;
    wire progRomAddress_10;
    wire \CONTROL.addrstack_reto_12 ;
    wire progRomAddress_12;
    wire \CONTROL.addrstack_10 ;
    wire \CONTROL.addrstack_reto_10 ;
    wire \CONTROL.programCounter_1_reto_8 ;
    wire N_423_cascade_;
    wire \CONTROL.programCounter_1_axb_8 ;
    wire \CONTROL.programCounter10 ;
    wire \CONTROL.programCounter_1_reto_9 ;
    wire \CONTROL.addrstack_reto_9 ;
    wire \CONTROL.N_424_cascade_ ;
    wire progRomAddress_9;
    wire CONTROL_addrstack_reto_8;
    wire N_423;
    wire progRomAddress_9_cascade_;
    wire \PROM.ROMDATA.dintern_adfltZ0Z_3 ;
    wire \CONTROL.tempCounterZ0Z_10 ;
    wire \CONTROL.programCounter_1_9 ;
    wire \CONTROL.tempCounterZ0Z_9 ;
    wire \INVCONTROL.tempCounter_10C_net ;
    wire \INVCONTROL.addrstackptr_0C_net ;
    wire \ALU.rshift_3_ns_1_2 ;
    wire \ALU.status_17_I_1_c_RNOZ0 ;
    wire \ALU.N_834_cascade_ ;
    wire busState_1_RNIDU0U1_2;
    wire \ALU.status_19_2_cascade_ ;
    wire romOut_4;
    wire \CONTROL.busState_1_RNI7U266Z0Z_2 ;
    wire bfn_12_11_0_;
    wire \ALU.mult_3_c3 ;
    wire \ALU.d_RNITK2D51Z0Z_2 ;
    wire \ALU.mult_3_c4 ;
    wire \ALU.d_RNIJBM6GZ0Z_3 ;
    wire \ALU.d_RNIKG0L11Z0Z_2 ;
    wire \ALU.mult_3_c5 ;
    wire \ALU.d_RNI9DAEHZ0Z_3 ;
    wire \ALU.d_RNI07V431Z0Z_2 ;
    wire \ALU.mult_3_c6 ;
    wire \ALU.d_RNIJ0U031Z0Z_2 ;
    wire \ALU.d_RNIV1LMHZ0Z_3 ;
    wire \ALU.mult_3_c7 ;
    wire \ALU.d_RNIS69AHZ0Z_3 ;
    wire \ALU.d_RNI12A911Z0Z_2 ;
    wire \ALU.mult_3_c8 ;
    wire \ALU.d_RNINIF011Z0Z_2 ;
    wire \ALU.mult_3_c9 ;
    wire \ALU.mult_3_c10 ;
    wire \ALU.d_RNIINE1HZ0Z_3 ;
    wire bfn_12_12_0_;
    wire \ALU.d_RNIMCVI41Z0Z_2 ;
    wire \ALU.d_RNITCCHHZ0Z_3 ;
    wire \ALU.mult_3_c11 ;
    wire \ALU.d_RNI18J1JZ0Z_3 ;
    wire \ALU.mult_3_c12 ;
    wire \ALU.mult_3_c13 ;
    wire \ALU.mult_3_c14 ;
    wire \ALU.d_RNI2IA441Z0Z_2 ;
    wire \ALU.d_RNI7SQI21Z0Z_2 ;
    wire \ALU.d_RNID31VFZ0Z_3 ;
    wire \ALU.d_RNIBRFE41Z0Z_2 ;
    wire \ALU.d_RNI9IN2HZ0Z_3 ;
    wire \ALU.a_RNI2N741Z0Z_12 ;
    wire \ALU.d_RNIJRM75Z0Z_5 ;
    wire DROM_ROMDATA_dintern_5ro;
    wire \ALU.d_RNIC0VE6Z0Z_5 ;
    wire \ALU.d_RNI693UNZ0Z_3 ;
    wire \ALU.mult_95_c_RNOZ0Z_0 ;
    wire \ALU.dout_6_ns_1_11_cascade_ ;
    wire \ALU.N_1144 ;
    wire \ALU.N_1096_cascade_ ;
    wire DROM_ROMDATA_dintern_11ro;
    wire aluOut_11_cascade_;
    wire \ALU.operand2_7_ns_1_11_cascade_ ;
    wire \ALU.b_RNI2TJC1Z0Z_11 ;
    wire \ALU.operand2_11_cascade_ ;
    wire \ALU.d_RNIMR627Z0Z_11_cascade_ ;
    wire \ALU.a_RNIV5PUZ0Z_11 ;
    wire \ALU.c_RNI3MHFZ0Z_11 ;
    wire \ALU.dout_3_ns_1_11 ;
    wire \ALU.dout_3_ns_1_10_cascade_ ;
    wire \ALU.dout_6_ns_1_10_cascade_ ;
    wire \ALU.N_1143_cascade_ ;
    wire \ALU.N_1095 ;
    wire aluOut_10_cascade_;
    wire \CONTROL.bus_0_10 ;
    wire ALU_N_1141;
    wire ALU_N_1093;
    wire \INVCONTROL.dout_7C_net ;
    wire gpuOut_c_7;
    wire N_168;
    wire N_168_cascade_;
    wire D7_in_c;
    wire \CONTROL.bus_7_ns_1_7_cascade_ ;
    wire PROM_ROMDATA_dintern_23ro;
    wire \CONTROL.bus_7_a1_1_8_cascade_ ;
    wire \CONTROL.bus_sx_8 ;
    wire gpuAddress_2;
    wire gpuAddress_3;
    wire gpuAddress_4;
    wire gpuAddress_5;
    wire gpuAddress_6;
    wire gpuAddress_7;
    wire gpuAddress_8;
    wire \INVCONTROL.gpuAddReg_2C_net ;
    wire \CONTROL.un1_busState119_1_i_0_1_cascade_ ;
    wire \CONTROL.gpuWrite_RNOZ0Z_2_cascade_ ;
    wire \CONTROL.busState96_cascade_ ;
    wire \CONTROL.busState96 ;
    wire \CONTROL.N_66_0 ;
    wire \CONTROL.gpuWrite_RNOZ0Z_0 ;
    wire gpuWrite;
    wire \INVCONTROL.gpuWriteC_net ;
    wire controlWord_21;
    wire \RAM.un1_WR_105_0Z0Z_3_cascade_ ;
    wire A5_c;
    wire \RAM.un1_WR_105_0Z0Z_11 ;
    wire controlWord_23;
    wire A7_c;
    wire controlWord_18;
    wire controlWord_18_cascade_;
    wire A2_c;
    wire \INVCONTROL.ramAddReg_5C_net ;
    wire \CONTROL.g0_3_i_1_0_cascade_ ;
    wire \CONTROL.N_4_1_cascade_ ;
    wire \INVCONTROL.addrstackptr_4C_net ;
    wire \CONTROL.N_81_0 ;
    wire \CONTROL.g0_3_i_a7_2_0 ;
    wire \CONTROL.N_429 ;
    wire \CONTROL.dout_reto_8 ;
    wire progRomAddress_15;
    wire \CONTROL.programCounter_1_11 ;
    wire \CONTROL.addrstack_1_4 ;
    wire \CONTROL.N_4_1 ;
    wire \CONTROL.un1_addrstackptr_c4_0 ;
    wire \CONTROL.addrstackptr_8_4 ;
    wire \CONTROL.programCounter_1_14 ;
    wire \CONTROL.programCounter_1_reto_14 ;
    wire \CONTROL.programCounter_1_reto_11 ;
    wire \CONTROL.dout_reto_11 ;
    wire \PROM.ROMDATA.m470_am ;
    wire \CONTROL.dout_reto_14 ;
    wire \CONTROL.programCounter_1_10 ;
    wire \CONTROL.programCounter11_reto_rep1 ;
    wire \CONTROL.programCounter_1_reto_10 ;
    wire \CONTROL.N_425 ;
    wire \CONTROL.programCounter_1_axb_1 ;
    wire \CONTROL.addrstackptr_8_1 ;
    wire \CONTROL.addrstackptr_RNI19JNL91Z0Z_0 ;
    wire \CONTROL.dout_reto_9 ;
    wire \ALU.d_RNILJMRC1Z0Z_8_cascade_ ;
    wire bfn_13_9_0_;
    wire \ALU.mult_7_c7 ;
    wire \ALU.d_RNITLGILZ0Z_7 ;
    wire \ALU.mult_7_c8 ;
    wire \ALU.d_RNIUFQIGZ0Z_7 ;
    wire \ALU.d_RNI8JFO21Z0Z_6 ;
    wire \ALU.mult_7_c9 ;
    wire \ALU.d_RNIKHEQHZ0Z_7 ;
    wire \ALU.d_RNIK9E841Z0Z_6 ;
    wire \ALU.mult_7_c10 ;
    wire \ALU.d_RNI73D441Z0Z_6 ;
    wire \ALU.mult_7_c11 ;
    wire \ALU.d_RNI7BDMHZ0Z_7 ;
    wire \ALU.mult_7_c12 ;
    wire \ALU.d_RNIBLU321Z0Z_6 ;
    wire \ALU.mult_7_c13 ;
    wire \ALU.mult_7_c14 ;
    wire bfn_13_10_0_;
    wire \ALU.d_RNIHNHG61Z0Z_6 ;
    wire \ALU.d_RNI4LU7E1Z0Z_6 ;
    wire \ALU.d_RNIA6P2IZ0Z_7 ;
    wire bfn_13_11_0_;
    wire \ALU.mult_1_c1 ;
    wire \ALU.d_RNIFBJI61Z0Z_0 ;
    wire \ALU.mult_1_c2 ;
    wire \ALU.d_RNIIOGRGZ0Z_1 ;
    wire \ALU.d_RNI67HQ21Z0Z_0 ;
    wire \ALU.mult_1_c3 ;
    wire \ALU.d_RNI8Q43IZ0Z_1 ;
    wire \ALU.d_RNIITFA41Z0Z_0 ;
    wire \ALU.mult_1_c4 ;
    wire \ALU.d_RNI5NE641Z0Z_0 ;
    wire \ALU.d_RNIUEFBIZ0Z_1 ;
    wire \ALU.mult_1_c5 ;
    wire \ALU.d_RNIRJ3VHZ0Z_1 ;
    wire \ALU.mult_1_c6 ;
    wire \ALU.d_RNI990621Z0Z_0 ;
    wire \ALU.mult_1_c7 ;
    wire \ALU.mult_1_c8 ;
    wire \ALU.d_RNIH49MHZ0Z_1 ;
    wire bfn_13_12_0_;
    wire \ALU.d_RNISP66IZ0Z_1 ;
    wire \ALU.mult_1_c9 ;
    wire \ALU.d_RNI0LDMJZ0Z_1 ;
    wire \ALU.d_RNIK8R951Z0Z_0 ;
    wire \ALU.mult_1_c10 ;
    wire \ALU.mult_1_c11 ;
    wire \ALU.d_RNI9UI0KZ0Z_1 ;
    wire \ALU.mult_1_c12 ;
    wire \ALU.mult_1_c13 ;
    wire \ALU.mult_3_c14_THRU_CO ;
    wire \ALU.d_RNI3D2O61Z0Z_2 ;
    wire \ALU.mult_1_c14 ;
    wire \ALU.d_RNI83GO51Z0Z_0 ;
    wire \ALU.d_RNIPIBO31Z0Z_0 ;
    wire \ALU.d_RNIIHC6LZ0Z_3 ;
    wire \ALU.d_RNITH0K51Z0Z_0 ;
    wire \ALU.d_RNI0H41KZ0Z_1 ;
    wire \ALU.d_RNIETL861Z0Z_0 ;
    wire \ALU.d_RNI8FM541Z0Z_0 ;
    wire \ALU.d_RNIGIF4D1Z0Z_2 ;
    wire CONTROL_addrstack_reto_11;
    wire N_426;
    wire progRomAddress_11;
    wire \ALU.d_RNILJMRC1_0Z0Z_8 ;
    wire \ALU.combOperand2_1Z0Z_0_cascade_ ;
    wire dintern_adflt_3_x;
    wire DROM_ROMDATA_dintern_0ro_cascade_;
    wire \CONTROL.bus_6_a0_sx_0 ;
    wire \ALU.mult_5_c_RNOZ0Z_0 ;
    wire \DROM.ROMDATA.dintern_0_0_NEW_0 ;
    wire \DROM.ROMDATA.dintern_0_0_OLDZ0Z_0 ;
    wire \INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C_net ;
    wire \INVCONTROL.dout_14C_net ;
    wire gpuOut_c_14;
    wire \CONTROL.ctrlOut_14 ;
    wire D14_in_c;
    wire \CONTROL.N_175_cascade_ ;
    wire N_191_cascade_;
    wire \CONTROL.busState_1_RNIRA1I6Z0Z_2_cascade_ ;
    wire \ALU.d_RNI8VHNHZ0Z_1 ;
    wire \ALU.dout_3_ns_1_12_cascade_ ;
    wire \ALU.dout_6_ns_1_12_cascade_ ;
    wire \ALU.N_1097 ;
    wire \ALU.N_1145_cascade_ ;
    wire aluOut_12_cascade_;
    wire \CONTROL.bus_0_12 ;
    wire gpuOut_c_11;
    wire D11_in_c;
    wire \CONTROL.N_172_cascade_ ;
    wire N_188;
    wire N_204;
    wire N_188_cascade_;
    wire \CONTROL.ctrlOut_11 ;
    wire \INVCONTROL.dout_11C_net ;
    wire gpuOut_c_12;
    wire D12_in_c;
    wire \CONTROL.N_173_cascade_ ;
    wire \CONTROL.N_189 ;
    wire \CONTROL.un1_busState14_1_i_o2_0_cascade_ ;
    wire \CONTROL.un1_busState12_2_i_a2_0_1_tz_0_cascade_ ;
    wire \CONTROL.N_244_cascade_ ;
    wire \INVCONTROL.aluReadBusC_net ;
    wire \CONTROL.un1_busState14_1_i_o2_0 ;
    wire \CONTROL.aluReadBus_r_1 ;
    wire \CONTROL.un1_busState14_1_i_a2_1_iZ0Z_1 ;
    wire \CONTROL.N_244 ;
    wire \CONTROL.N_58 ;
    wire \CONTROL.N_89 ;
    wire \CONTROL.N_89_cascade_ ;
    wire \CONTROL.aluReadBus_1_sqmuxa_0_a2_0Z0Z_0_cascade_ ;
    wire \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_0 ;
    wire gpuOut_c_10;
    wire D10_in_c;
    wire \CONTROL.N_171_cascade_ ;
    wire \CONTROL.N_187 ;
    wire \INVCONTROL.dout_10C_net ;
    wire gpuOut_c_0;
    wire D0_in_c;
    wire \CONTROL.N_161_cascade_ ;
    wire \PROM.ROMDATA.m520 ;
    wire gpuOut_c_15;
    wire N_176;
    wire D15_in_c;
    wire N_176_cascade_;
    wire \PROM.ROMDATA.m471_ns ;
    wire \INVCONTROL.dout_15C_net ;
    wire gpuOut_c_8;
    wire \CONTROL.ctrlOut_8 ;
    wire A0_c;
    wire A1_c;
    wire controlWord_26;
    wire controlWord_27;
    wire A10_c;
    wire A11_c;
    wire \RAM.un1_WR_105_0Z0Z_9 ;
    wire controlWord_25;
    wire A9_c;
    wire controlWord_24;
    wire A8_c;
    wire \INVCONTROL.ramAddReg_0C_net ;
    wire \CONTROL.g1_0 ;
    wire \CONTROL.addrstack_1_1 ;
    wire \CONTROL.g1_0_cascade_ ;
    wire \INVCONTROL.addrstackptr_1C_net ;
    wire \CONTROL.g0_1_i_a6Z0Z_4_cascade_ ;
    wire \CONTROL.N_9 ;
    wire \CONTROL.g0_0_1 ;
    wire \CONTROL.N_366 ;
    wire \CONTROL.g0_1_i_3 ;
    wire \CONTROL.addrstack_15 ;
    wire \CONTROL.addrstack_reto_15 ;
    wire controlWord_30;
    wire \INVCONTROL.ramAddReg_14C_net ;
    wire \ALU.mult_173_c_RNOZ0Z_0 ;
    wire bfn_14_8_0_;
    wire \ALU.mult_5_c5 ;
    wire \ALU.d_RNIFGNR61Z0Z_4 ;
    wire \ALU.mult_5_c6 ;
    wire \ALU.d_RNICP0UGZ0Z_5 ;
    wire \ALU.d_RNI6CL331Z0Z_4 ;
    wire \ALU.mult_5_c7 ;
    wire \ALU.d_RNI2RK5IZ0Z_5 ;
    wire \ALU.mult_5_c8 ;
    wire \ALU.d_RNIOFVDIZ0Z_5 ;
    wire \ALU.d_RNI5SIF41Z0Z_4 ;
    wire \ALU.mult_5_c9 ;
    wire \ALU.d_RNILKJ1IZ0Z_5 ;
    wire \ALU.d_RNIJTUN21Z0Z_4 ;
    wire \ALU.mult_5_c10 ;
    wire \ALU.d_RNI6HBMGZ0Z_5 ;
    wire \ALU.d_RNI9E4F21Z0Z_4 ;
    wire \ALU.mult_5_c11 ;
    wire \ALU.mult_5_c12 ;
    wire \ALU.d_RNIB5POHZ0Z_5 ;
    wire \ALU.d_RNIPNF141Z0Z_4 ;
    wire bfn_14_9_0_;
    wire \ALU.d_RNI88K161Z0Z_4 ;
    wire \ALU.d_RNIMQM8IZ0Z_5 ;
    wire \ALU.mult_5_c13 ;
    wire \ALU.mult_7_c14_THRU_CO ;
    wire \ALU.d_RNIKDVI51Z0Z_4 ;
    wire \ALU.d_RNIRU9M31Z0Z_6 ;
    wire \ALU.mult_5_c14 ;
    wire bus_0_12;
    wire \ALU.mult_239_c_RNOZ0Z_0 ;
    wire \ALU.mult_239_c_RNOZ0 ;
    wire \ALU.mult_1_2 ;
    wire bfn_14_10_0_;
    wire \ALU.mult_1_3 ;
    wire \ALU.mult_17_c2 ;
    wire \ALU.mult_3_4 ;
    wire \ALU.mult_1_4 ;
    wire \ALU.mult_17_c3 ;
    wire \ALU.mult_1_5 ;
    wire \ALU.mult_3_5 ;
    wire \ALU.mult_17_c4 ;
    wire \ALU.mult_1_6 ;
    wire \ALU.mult_3_6 ;
    wire \ALU.mult_17_c5 ;
    wire \ALU.mult_1_7 ;
    wire \ALU.mult_3_7 ;
    wire \ALU.mult_17_c6 ;
    wire \ALU.mult_1_8 ;
    wire \ALU.mult_3_8 ;
    wire \ALU.mult_17_c7 ;
    wire \ALU.mult_1_9 ;
    wire \ALU.mult_3_9 ;
    wire \ALU.mult_17_c8 ;
    wire \ALU.mult_17_c9 ;
    wire \ALU.mult_3_10 ;
    wire \ALU.mult_1_10 ;
    wire bfn_14_11_0_;
    wire \ALU.mult_1_11 ;
    wire \ALU.mult_3_11 ;
    wire \ALU.mult_17_c10 ;
    wire \ALU.mult_1_12 ;
    wire \ALU.mult_3_12 ;
    wire \ALU.mult_17_c11 ;
    wire \ALU.mult_1_13 ;
    wire \ALU.mult_3_13 ;
    wire \ALU.mult_17_c12 ;
    wire \ALU.mult_1_14 ;
    wire \ALU.mult_3_14 ;
    wire \ALU.mult_17_c13 ;
    wire \ALU.mult_227_c_RNIBPRVZ0Z92 ;
    wire \ALU.mult_83_c_RNIKEU6BZ0Z2 ;
    wire \ALU.mult_17_c14 ;
    wire \ALU.d_RNIHU6RLZ0Z_1 ;
    wire \ALU.d_RNI2E4JE1Z0Z_4 ;
    wire \ALU.N_860 ;
    wire \ALU.mult_5_c_RNOZ0 ;
    wire \ALU.d_RNI290AE1Z0Z_0 ;
    wire \ALU.d_RNI5MTIOZ0Z_1 ;
    wire busState_1_RNICT0U1_2_cascade_;
    wire busState_1_RNICT0U1_2;
    wire N_227_0_cascade_;
    wire \ALU.status_18_cry_2_c_RNOZ0 ;
    wire DROM_ROMDATA_dintern_2ro;
    wire \DROM.ROMDATA.dintern_0_0_NEW_2 ;
    wire \DROM.ROMDATA.dintern_0_0_OLDZ0Z_2 ;
    wire \INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C_net ;
    wire \DROM.ROMDATA.dintern_0_0_sr_enZ0 ;
    wire \ALU.eZ0Z_4 ;
    wire \ALU.eZ0Z_10 ;
    wire \ALU.eZ0Z_11 ;
    wire CONSTANT_ONE_NET;
    wire \ALU.dout_6_ns_1_6_cascade_ ;
    wire \ALU.eZ0Z_6 ;
    wire \ALU.dout_3_ns_1_6_cascade_ ;
    wire \ALU.N_1091_cascade_ ;
    wire \ALU.N_1139 ;
    wire aluOut_6_cascade_;
    wire \ALU.d_RNIR3N75Z0Z_6 ;
    wire \ALU.dout_6_ns_1_1_cascade_ ;
    wire ALU_N_1134_cascade_;
    wire \CONTROL.operand1_ne_RNIBQE03Z0Z_0 ;
    wire busState_1_RNI9P5V3_2;
    wire \ALU.dout_3_ns_1_1_cascade_ ;
    wire ALU_N_1086_cascade_;
    wire ALU_N_1134;
    wire \INVCONTROL.operand1_ne_1C_net ;
    wire \ALU.d_RNIHD7AOZ0Z_7 ;
    wire \CONTROL.operand1_ne_RNIHKCU2Z0Z_0_cascade_ ;
    wire operand1_ne_RNIDN8E7_0;
    wire \ALU.dout_6_ns_1_0 ;
    wire aluOperand1_2_rep1;
    wire \ALU.dout_3_ns_1_0_cascade_ ;
    wire ALU_N_1085_cascade_;
    wire \CONTROL.operand1_ne_RNIHKCU2_0Z0Z_0 ;
    wire ALU_N_1133;
    wire ALU_N_1085;
    wire \ALU.operand2_3_ns_1_2_cascade_ ;
    wire \ALU.N_1199_cascade_ ;
    wire \ALU.N_1199 ;
    wire \ALU.c_RNIJ1JO4_0Z0Z_2_cascade_ ;
    wire \ALU.c_RNIJ1JO4Z0Z_2 ;
    wire \ALU.d_RNIARKGBZ0Z_2 ;
    wire \ALU.operand2_6_ns_1_2 ;
    wire \ALU.N_1247 ;
    wire gpuOut_c_13;
    wire D13_in_c;
    wire \CONTROL.N_174_cascade_ ;
    wire \CONTROL.N_169 ;
    wire D8_in_c;
    wire \CONTROL.N_185 ;
    wire \INVCONTROL.busState_1_2C_net ;
    wire D4_in_c;
    wire \CONTROL.busState_1_RNIU83C1_0Z0Z_2 ;
    wire D2_in_c;
    wire N_228_0;
    wire \CONTROL.busState_1_RNILAEH1Z0Z_2 ;
    wire gpuOut_c_1;
    wire N_162;
    wire D1_in_c;
    wire N_162_cascade_;
    wire \INVCONTROL.busState_1_1C_net ;
    wire \CONTROL.N_180 ;
    wire gpuOut_c_3;
    wire N_164;
    wire D3_in_c;
    wire N_164_cascade_;
    wire controlWord_16;
    wire CONTROL_romAddReg_7_0;
    wire controlWord_17;
    wire controlWord_17_cascade_;
    wire CONTROL_romAddReg_7_1;
    wire \INVCONTROL.dout_1C_net ;
    wire \CONTROL.N_430 ;
    wire \CONTROL.un1_busState98_1_1_0Z0Z_0 ;
    wire \CONTROL.programCounter_1_15 ;
    wire \CONTROL.programCounter_1_reto_15 ;
    wire \CONTROL.ctrlOut_15 ;
    wire \CONTROL.dout_reto_15 ;
    wire \PROM.ROMDATA.m465_am ;
    wire \CONTROL.ctrlOut_7 ;
    wire \CONTROL.tempCounterZ0Z_0 ;
    wire \CONTROL.tempCounterZ0Z_5 ;
    wire \CONTROL.tempCounterZ0Z_3 ;
    wire \CONTROL.programCounter_1_8 ;
    wire \CONTROL.tempCounterZ0Z_8 ;
    wire \INVCONTROL.tempCounter_0C_net ;
    wire \CONTROL.tempCounterZ0Z_4 ;
    wire \CONTROL.tempCounterZ0Z_1 ;
    wire \CONTROL.tempCounterZ0Z_7 ;
    wire \CONTROL.tempCounterZ0Z_12 ;
    wire \CONTROL.tempCounterZ0Z_2 ;
    wire \INVCONTROL.tempCounter_4C_net ;
    wire \CONTROL.addrstack_1_i ;
    wire \ALU.d_RNII2KJ41Z0Z_4 ;
    wire bus_4;
    wire \ALU.mult_173_c_RNOZ0 ;
    wire \ALU.mult_5_6 ;
    wire bfn_15_9_0_;
    wire \ALU.mult_7_7 ;
    wire \ALU.mult_5_7 ;
    wire \ALU.mult_19_c6 ;
    wire \ALU.mult_7_8 ;
    wire \ALU.mult_5_8 ;
    wire \ALU.mult_19_c7 ;
    wire \ALU.mult_7_9 ;
    wire \ALU.mult_5_9 ;
    wire \ALU.mult_19_c8 ;
    wire \ALU.mult_7_10 ;
    wire \ALU.mult_5_10 ;
    wire \ALU.mult_19_c9 ;
    wire \ALU.mult_7_11 ;
    wire \ALU.mult_5_11 ;
    wire \ALU.mult_19_c10 ;
    wire \ALU.mult_5_12 ;
    wire \ALU.mult_7_12 ;
    wire \ALU.mult_19_c11 ;
    wire \ALU.mult_5_13 ;
    wire \ALU.mult_7_13 ;
    wire \ALU.mult_19_c12 ;
    wire \ALU.mult_19_c13 ;
    wire \ALU.mult_5_14 ;
    wire \ALU.mult_7_14 ;
    wire bfn_15_10_0_;
    wire \ALU.mult_19_c14 ;
    wire \ALU.mult_19_c14_THRU_CO ;
    wire \ALU.mult_3_2 ;
    wire \ALU.mult_486_c_RNIPJD0IZ0Z5_cascade_ ;
    wire \ALU.combOperand2_0_5 ;
    wire \ALU.d_RNICGRJGZ0Z_1 ;
    wire \ALU.addsub_cry_4_c_RNI2RZ0Z6596 ;
    wire \ALU.d_RNIBVMTLZ0Z_5 ;
    wire \ALU.d_RNIVMDLOZ0Z_5 ;
    wire \ALU.mult_3_3 ;
    wire busState_1_RNIBS0U1_2;
    wire operand1_ne_RNIR8FK7_0;
    wire \ALU.status_19_0_cascade_ ;
    wire \ALU.mult_95_c_RNOZ0 ;
    wire \ALU.mult_3 ;
    wire \ALU.addsub_cry_2_c_RNIUFTGNZ0Z3_cascade_ ;
    wire \ALU.mult_388_c_RNIBULDPZ0Z3 ;
    wire \ALU.mult_388_c_RNIEAAJHZ0Z7_cascade_ ;
    wire bus_3;
    wire \ALU.mult_388_c_RNIEAAJHZ0Z7 ;
    wire \ALU.mult_388_c_RNIPGN6QZ0Z7_cascade_ ;
    wire \ALU.a_15_d_sZ0Z_5 ;
    wire \ALU.mult_2 ;
    wire \ALU.log_1_2 ;
    wire \ALU.a_15_d_sZ0Z_3 ;
    wire \ALU.addsub_cry_1_c_RNI8FKPLZ0Z3_cascade_ ;
    wire \ALU.mult_5_c_RNI6ET5DZ0Z3 ;
    wire \ALU.addsub_cry_1_c_RNIJP8KZ0Z37_cascade_ ;
    wire \ALU.addsub_cry_1_c_RNIJP8KZ0Z37 ;
    wire \ALU.addsub_cry_1_c_RNIICPECZ0Z7_cascade_ ;
    wire \ALU.dout_3_ns_1_9_cascade_ ;
    wire \ALU.dout_6_ns_1_9_cascade_ ;
    wire \ALU.N_1094 ;
    wire \ALU.N_1142_cascade_ ;
    wire aluOut_9_cascade_;
    wire h_2;
    wire \ALU.dout_6_ns_1_2_cascade_ ;
    wire \ALU.aZ0Z_2 ;
    wire \ALU.eZ0Z_2 ;
    wire \ALU.dout_3_ns_1_2_cascade_ ;
    wire \ALU.N_1087_cascade_ ;
    wire \ALU.N_1135 ;
    wire ALU_N_1086;
    wire \CONTROL.operand1_ne_RNIBQE03_0Z0Z_0 ;
    wire \PROM.ROMDATA.m238_am_1_cascade_ ;
    wire \PROM.ROMDATA.m238_am_cascade_ ;
    wire \PROM.ROMDATA.m244_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m244_ns_1 ;
    wire \INVCONTROL.operand1_fast_ne_1C_net ;
    wire \ALU.dout_6_ns_1_3_cascade_ ;
    wire \ALU.dout_3_ns_1_3_cascade_ ;
    wire \ALU.N_1136 ;
    wire \ALU.N_1088_cascade_ ;
    wire aluOut_3_cascade_;
    wire busState_1_RNIH16V3_2;
    wire \ALU.dout_3_ns_1_13_cascade_ ;
    wire aluOperand1_2_rep2;
    wire \ALU.dout_6_ns_1_13_cascade_ ;
    wire \ALU.N_1098 ;
    wire \ALU.N_1146_cascade_ ;
    wire \CONTROL.N_190 ;
    wire \CONTROL.bus_7_a1_1_8 ;
    wire aluOut_13_cascade_;
    wire \CONTROL.bus_0_13 ;
    wire \ALU.c_RNIJMOB4_0Z0Z_1_cascade_ ;
    wire \ALU.d_RNID42JAZ0Z_1 ;
    wire \ALU.operand2_6_ns_1_1 ;
    wire \ALU.N_1246 ;
    wire \ALU.operand2_3_ns_1_1_cascade_ ;
    wire \ALU.N_1198 ;
    wire \ALU.combOperand2_d_bmZ0Z_1 ;
    wire \ALU.N_1198_cascade_ ;
    wire \ALU.c_RNIJMOB4Z0Z_1 ;
    wire \CONTROL.g0_3_i_a7_2_1 ;
    wire \CONTROL.N_5_cascade_ ;
    wire \CONTROL.addrstackptr_8_3 ;
    wire gpuOut_c_2;
    wire \CONTROL.N_163 ;
    wire \CONTROL.g0_3_i_2_1 ;
    wire \CONTROL.un1_addrstackptr_c3_0 ;
    wire \CONTROL.addrstack_1_3 ;
    wire \CONTROL.N_5 ;
    wire \CONTROL.addrstackptrZ0Z_3 ;
    wire \INVCONTROL.addrstackptr_3C_net ;
    wire \INVCONTROL.aluOperation_ne_1C_net ;
    wire \CONTROL.N_83_0_cascade_ ;
    wire \CONTROL.m28_0_120_i_i_4 ;
    wire \CONTROL.N_75_0 ;
    wire \CONTROL.N_75_0_cascade_ ;
    wire \CONTROL.m38_i_2 ;
    wire \CONTROL.N_339 ;
    wire \CONTROL.N_219_cascade_ ;
    wire \CONTROL.m28_0_120_i_i_a2_0_0_cascade_ ;
    wire \CONTROL.busState_1_RNO_1Z0Z_1_cascade_ ;
    wire \CONTROL.busState_1_RNO_0Z0Z_1 ;
    wire \CONTROL.g0_3_i_1_1 ;
    wire \CONTROL.N_350_1 ;
    wire \CONTROL.N_345 ;
    wire \CONTROL.N_346 ;
    wire \CONTROL.N_255 ;
    wire \CONTROL.N_345_cascade_ ;
    wire ramWrite;
    wire \INVCONTROL.ramWriteC_net ;
    wire \CONTROL.un1_busState114_1_0Z0Z_0 ;
    wire \CONTROL.ctrlOut_10 ;
    wire \CONTROL.dout_reto_10 ;
    wire \PROM.ROMDATA.m1_cascade_ ;
    wire \PROM.ROMDATA.m2_cascade_ ;
    wire \ALU.mult_7_6 ;
    wire \ALU.status_18_cry_0_c_RNOZ0 ;
    wire \ALU.mult_5_4 ;
    wire \ALU.mult_17_4 ;
    wire \ALU.mult_391_c_RNIEC73TZ0Z4 ;
    wire bfn_16_9_0_;
    wire \ALU.mult_17_5 ;
    wire \ALU.mult_5 ;
    wire \ALU.mult_25_c4 ;
    wire \ALU.mult_173_c_RNIO8AOZ0Z16 ;
    wire \ALU.mult_17_6 ;
    wire \ALU.mult_25_c5 ;
    wire \ALU.mult_19_7 ;
    wire \ALU.mult_17_7 ;
    wire \ALU.mult_25_c6 ;
    wire \ALU.mult_17_8 ;
    wire \ALU.mult_19_8 ;
    wire \ALU.mult_25_c7 ;
    wire \ALU.mult_17_9 ;
    wire \ALU.mult_19_9 ;
    wire \ALU.mult_25_c8 ;
    wire \ALU.mult_19_10 ;
    wire \ALU.mult_17_10 ;
    wire \ALU.mult_25_c9 ;
    wire \ALU.mult_17_11 ;
    wire \ALU.mult_19_11 ;
    wire \ALU.mult_25_c10 ;
    wire \ALU.mult_25_c11 ;
    wire \ALU.mult_17_12 ;
    wire \ALU.mult_19_12 ;
    wire bfn_16_10_0_;
    wire \ALU.mult_17_13 ;
    wire \ALU.mult_19_13 ;
    wire \ALU.mult_25_c12 ;
    wire \ALU.mult_17_14 ;
    wire \ALU.mult_19_14 ;
    wire \ALU.mult_25_c13 ;
    wire \ALU.mult_424_c_RNIUVTALZ0Z4 ;
    wire \ALU.mult_25_c14 ;
    wire \ALU.d_RNIUT8OG4Z0Z_0 ;
    wire \ALU.lshift_3_ns_1_14 ;
    wire \ALU.N_646_cascade_ ;
    wire \ALU.lshift_15_ns_1_14_cascade_ ;
    wire g_2;
    wire g_4;
    wire g_6;
    wire g_10;
    wire g_11;
    wire f_2;
    wire f_10;
    wire f_11;
    wire CONSTANT_ZERO_NET;
    wire \ALU.cZ0Z_2 ;
    wire \ALU.cZ0Z_4 ;
    wire \ALU.cZ0Z_6 ;
    wire \ALU.cZ0Z_10 ;
    wire \ALU.cZ0Z_11 ;
    wire \ALU.dZ0Z_2 ;
    wire \ALU.dZ0Z_6 ;
    wire \ALU.dZ0Z_10 ;
    wire \ALU.dZ0Z_11 ;
    wire \ALU.d_RNI6DCTZ0Z_11 ;
    wire \INVCONTROL.operand2_fast_ne_2C_net ;
    wire \ALU.N_920 ;
    wire \ALU.operand2_3_ns_1_15 ;
    wire \ALU.dout_3_ns_1_15_cascade_ ;
    wire aluOperand1_fast_2;
    wire aluOperand1_fast_1;
    wire \CONTROL.increment28lto5_1_1_3 ;
    wire \CONTROL.increment28lto5_1_1_1_cascade_ ;
    wire \CONTROL.g0_3_i_a7Z0Z_3 ;
    wire \PROM.ROMDATA.m221cf1_cascade_ ;
    wire \PROM.ROMDATA.m221cf1 ;
    wire \INVCONTROL.operand1_ne_0C_net ;
    wire \CONTROL.un1_busState98_1_0_0_0 ;
    wire \PROM.ROMDATA.m217 ;
    wire \PROM.ROMDATA.m221cf0 ;
    wire \CONTROL.increment28lto5_1_1_0 ;
    wire \CONTROL.N_101_0 ;
    wire \CONTROL.N_320_cascade_ ;
    wire \CONTROL.un1_busState103_0_0_cascade_ ;
    wire \INVCONTROL.aluParams_1_0C_net ;
    wire \CONTROL.N_95_0 ;
    wire \CONTROL.N_318 ;
    wire \CONTROL.N_340_cascade_ ;
    wire \INVCONTROL.aluParams_1_ne_1C_net ;
    wire \CONTROL.un1_busState103_0_0 ;
    wire \CONTROL.un1_busState114_2_0_0_xZ0Z0_cascade_ ;
    wire \CONTROL.un1_busState114_2_0_0_xZ0Z1 ;
    wire \CONTROL.un1_busState114_2_0_0_0_cascade_ ;
    wire \CONTROL.aluReadBus_1_sqmuxa_0_a2_2Z0Z_0 ;
    wire \CONTROL.N_83_0 ;
    wire \CONTROL.N_48_0_cascade_ ;
    wire \INVCONTROL.aluOperation_4C_net ;
    wire \CONTROL.un1_controlWord_14_i_0 ;
    wire \CONTROL.N_87_0 ;
    wire \CONTROL.un1_busState97_1_0_1_0 ;
    wire \CONTROL.dout_reto_7 ;
    wire \CONTROL.addrstack_reto_7 ;
    wire \CONTROL.N_422_cascade_ ;
    wire progRomAddress_7_cascade_;
    wire \INVCONTROL.dout_2C_net ;
    wire \CONTROL.N_420_cascade_ ;
    wire \CONTROL.programCounter_1_axb_5 ;
    wire \CONTROL.programCounter_1_axb_0 ;
    wire \CONTROL.N_105_i ;
    wire \CONTROL.N_427 ;
    wire PROM_ROMDATA_dintern_5ro_cascade_;
    wire \CONTROL.N_80_0 ;
    wire \CONTROL.g0_1_i_3Z0Z_1 ;
    wire \CONTROL.N_384_0 ;
    wire \CONTROL.N_209_cascade_ ;
    wire \CONTROL.un1_busState114_1_0_0_0 ;
    wire \CONTROL.N_349_cascade_ ;
    wire \CONTROL.N_246 ;
    wire \CONTROL.m38_i_1 ;
    wire \CONTROL.N_348 ;
    wire \CONTROL.programCounter_1_12 ;
    wire \CONTROL.programCounter_1_reto_12 ;
    wire controlWord_1_cascade_;
    wire \PROM.ROMDATA.m506_cascade_ ;
    wire \PROM.ROMDATA.N_571_mux ;
    wire N_177;
    wire \ALU.d_RNI64MA6Z0Z_0_cascade_ ;
    wire \ALU.log_1_3_ns_1_1_0_cascade_ ;
    wire \ALU.log_1_3_ns_1_0_cascade_ ;
    wire \ALU.log_1_0_cascade_ ;
    wire \ALU.status_8_5_0_cascade_ ;
    wire \ALU.mult_365_c_RNOZ0 ;
    wire bfn_17_9_0_;
    wire \ALU.c_RNIF6GEF1Z0Z_12 ;
    wire \ALU.c_RNINUT6PZ0Z_13 ;
    wire \ALU.mult_13_c13 ;
    wire \ALU.c_RNIS83N71Z0Z_12 ;
    wire \ALU.mult_13_c14 ;
    wire \ALU.d_RNIL4PC21Z0Z_6 ;
    wire \ALU.mult_5_5 ;
    wire bfn_17_10_0_;
    wire \ALU.mult_9_9 ;
    wire \ALU.mult_25_9 ;
    wire \ALU.mult_29_c8 ;
    wire \ALU.mult_29_c9 ;
    wire \ALU.mult_25_11 ;
    wire \ALU.mult_29_c10 ;
    wire \ALU.mult_29_c11 ;
    wire \ALU.mult_25_13 ;
    wire \ALU.mult_29_c12 ;
    wire \ALU.mult_25_14 ;
    wire \ALU.mult_29_c13 ;
    wire \ALU.mult_516_c_RNI98SKDCZ0 ;
    wire \ALU.mult_29_c14 ;
    wire bus_0_10;
    wire \ALU.mult_10 ;
    wire \ALU.mult_549_c_RNIB6TIDGZ0_cascade_ ;
    wire \ALU.a_15_am_1_10 ;
    wire \ALU.mult_549_c_RNIE7260OZ0_cascade_ ;
    wire \ALU.aZ0Z_10 ;
    wire \ALU.a_15_m3_sZ0Z_13_cascade_ ;
    wire \ALU.a32Z0Z_0_cascade_ ;
    wire \ALU.aZ0Z_1 ;
    wire \ALU.d_RNICUA7B5Z0Z_0_cascade_ ;
    wire \ALU.d_RNIL3JT71Z0Z_0 ;
    wire \ALU.N_556 ;
    wire \ALU.N_556_cascade_ ;
    wire \ALU.d_RNI3MGBH1Z0Z_1 ;
    wire \ALU.status_17_I_39_c_RNOZ0 ;
    wire \ALU.mult_365_c_RNOZ0Z_0 ;
    wire \ALU.N_572 ;
    wire bus_11;
    wire \ALU.mult_11 ;
    wire \ALU.mult_552_c_RNI70R9DAZ0_cascade_ ;
    wire \ALU.rshift_11 ;
    wire \ALU.a_15_am_rn_0_11 ;
    wire \ALU.mult_552_c_RNI70R9DAZ0 ;
    wire \ALU.mult_552_c_RNIOT7VLFZ0_cascade_ ;
    wire \ALU.aZ0Z_11 ;
    wire \ALU.a_15_am_snZ0Z_11 ;
    wire h_1;
    wire \ALU.mult_6 ;
    wire \ALU.mult_489_c_RNIGEUL1AZ0_cascade_ ;
    wire \ALU.mult_489_c_RNIGEUL1AZ0 ;
    wire \ALU.mult_489_c_RNIPGBQMCZ0Z_0_cascade_ ;
    wire \ALU.mult_489_c_RNIPGBQMCZ0 ;
    wire \ALU.mult_489_c_RNI1J3GCUZ0_cascade_ ;
    wire h_6;
    wire \ALU.a_15_m2_d_d_ns_1_0_0_cascade_ ;
    wire bus_0;
    wire \ALU.lshift62 ;
    wire \ALU.d_RNI4D6E01Z0Z_0_cascade_ ;
    wire \ALU.d_RNIQQ9O83Z0Z_0_cascade_ ;
    wire \ALU.d_RNI4HL061Z0Z_0 ;
    wire \ALU.d_RNINUGCF4Z0Z_0_cascade_ ;
    wire \ALU.aZ0Z_0 ;
    wire h_0;
    wire \ALU.e_RNI933SZ0Z_0 ;
    wire \ALU.c_RNIDFF01Z0Z_0_cascade_ ;
    wire \ALU.d_RNI0G5DZ0Z_0 ;
    wire \ALU.b_RNIS3POZ0Z_0_cascade_ ;
    wire \ALU.operand2_7_ns_1_0 ;
    wire \ALU.operand2_0 ;
    wire \ALU.dZ0Z_3 ;
    wire \ALU.operand2_6_ns_1_3_cascade_ ;
    wire \ALU.aZ0Z_3 ;
    wire \ALU.eZ0Z_3 ;
    wire \ALU.cZ0Z_3 ;
    wire g_3;
    wire \ALU.operand2_3_ns_1_3_cascade_ ;
    wire \ALU.N_1200_cascade_ ;
    wire \ALU.N_1248 ;
    wire \ALU.d_RNIGMEO4Z0Z_3_cascade_ ;
    wire \ALU.combOperand2_d_bmZ0Z_3 ;
    wire \ALU.d_RNI2CUG6Z0Z_3 ;
    wire gpuOut_c_4;
    wire \CONTROL.N_165 ;
    wire h_9;
    wire \ALU.e_RNICGJMZ0Z_9 ;
    wire \ALU.d_RNIKKNJZ0Z_9 ;
    wire \ALU.operand2_7_ns_1_9_cascade_ ;
    wire \ALU.b_RNIG8BVZ0Z_9 ;
    wire \ALU.operand2_9_cascade_ ;
    wire \ALU.status_RNO_2Z0Z_0 ;
    wire \ALU.status_e_1_0 ;
    wire \CONTROL.increment28lto5_1Z0Z_1_cascade_ ;
    wire PROM_ROMDATA_dintern_8ro;
    wire \CONTROL.increment28lto5_1_1_2_cascade_ ;
    wire PROM_ROMDATA_dintern_7ro;
    wire \CONTROL.increment28lto5_1Z0Z_2 ;
    wire \INVCONTROL.aluOperation_ne_5C_net ;
    wire \CONTROL.N_48_0 ;
    wire controlWord_6_cascade_;
    wire \CONTROL.N_140_0 ;
    wire \CONTROL.un1_busState96_1_i_i_a2_1Z0Z_1_cascade_ ;
    wire \CONTROL.un1_busState96_1_i_i_a2_0Z0Z_1 ;
    wire \CONTROL.un1_busState96_1_i_iZ0Z_0_cascade_ ;
    wire controlWord_5_cascade_;
    wire \CONTROL.N_134_0 ;
    wire \CONTROL.N_327 ;
    wire \CONTROL.N_133_0_1 ;
    wire PROM_ROMDATA_dintern_3ro_cascade_;
    wire \CONTROL.g0_3_i_2_0 ;
    wire \CONTROL.g0_2_i_a7Z0Z_3 ;
    wire \CONTROL.g0_2_i_a7Z0Z_2 ;
    wire \CONTROL.g0_2_i_2_cascade_ ;
    wire \CONTROL.addrstack_1_2 ;
    wire \CONTROL.addrstackptrZ0Z_1 ;
    wire \CONTROL.N_5_0_cascade_ ;
    wire \CONTROL.g0_12_1_cascade_ ;
    wire \CONTROL.addrstackptr_8_2 ;
    wire controlWord_4_cascade_;
    wire \CONTROL.N_5_0 ;
    wire \CONTROL.g0_12_1 ;
    wire \INVCONTROL.addrstackptr_2C_net ;
    wire \CONTROL.N_360 ;
    wire \CONTROL.N_362 ;
    wire \CONTROL.m28_0_120_i_i_0 ;
    wire \CONTROL.N_321 ;
    wire \CONTROL.N_338 ;
    wire PROM_ROMDATA_dintern_0ro;
    wire PROM_ROMDATA_dintern_0ro_cascade_;
    wire \CONTROL.un1_busState_0_sqmuxa_i_a2_0 ;
    wire \CONTROL.N_304_0 ;
    wire \PROM.ROMDATA.m433_ns ;
    wire \PROM.ROMDATA.m294_bm_cascade_ ;
    wire \PROM.ROMDATA.m31_cascade_ ;
    wire \CONTROL.ctrlOut_12 ;
    wire \CONTROL.dout_reto_12 ;
    wire \PROM.ROMDATA.m391_cascade_ ;
    wire \PROM.ROMDATA.m433_bm ;
    wire \PROM.ROMDATA.m382_ns ;
    wire busState_1_RNIAR0U1_2;
    wire N_225_0_cascade_;
    wire \ALU.mult_13_15 ;
    wire \ALU.mult_15_14_cascade_ ;
    wire \ALU.mult_13_14 ;
    wire \ALU.lshift_3_ns_1_15_cascade_ ;
    wire \ALU.d_RNI64MA6Z0Z_0 ;
    wire N_225_0;
    wire \ALU.mult_25_12 ;
    wire \ALU.mult_13_12_cascade_ ;
    wire \ALU.mult_467_c_RNICRDK6BZ0 ;
    wire \ALU.mult_13_12 ;
    wire bfn_18_10_0_;
    wire \ALU.mult_13_13 ;
    wire \ALU.mult_27_13 ;
    wire \ALU.mult_27_c12 ;
    wire \ALU.mult_365_c_RNI8ALOZ0Z96 ;
    wire \ALU.mult_27_14 ;
    wire \ALU.mult_27_c13 ;
    wire \ALU.mult_27_c14 ;
    wire \ALU.mult_27_c14_THRU_CO ;
    wire \ALU.mult_9 ;
    wire \ALU.mult_13 ;
    wire \ALU.N_642 ;
    wire \ALU.d_RNIULN025Z0Z_2_cascade_ ;
    wire \ALU.d_RNIULN025_0Z0Z_2 ;
    wire \ALU.lshift_10_cascade_ ;
    wire \ALU.c_RNIO0KOKEZ0Z_10_cascade_ ;
    wire \ALU.bZ0Z_10 ;
    wire \ALU.N_1025 ;
    wire \ALU.N_864 ;
    wire \ALU.N_965_cascade_ ;
    wire \ALU.d_RNIFHCRU4Z0Z_2 ;
    wire \ALU.mult_15_15 ;
    wire \ALU.c_RNINT9PO2Z0Z_10 ;
    wire \ALU.c_RNI890LZ0Z_13 ;
    wire \ALU.a_RNI4P741Z0Z_13_cascade_ ;
    wire \ALU.d_RNIAHCTZ0Z_13 ;
    wire \ALU.operand2_7_ns_1_13_cascade_ ;
    wire \ALU.b_RNI61KC1Z0Z_13 ;
    wire \ALU.operand2_13 ;
    wire bus_0_13;
    wire \ALU.operand2_13_cascade_ ;
    wire \ALU.d_RNI02EVNBZ0Z_4 ;
    wire \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ;
    wire \ALU.addsub_cry_1_c_RNIICPECZ0Z7 ;
    wire \ALU.bZ0Z_2 ;
    wire \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9 ;
    wire \ALU.addsub_cry_4_c_RNI5L6IQAZ0 ;
    wire \ALU.bZ0Z_6 ;
    wire \ALU.bZ0Z_3 ;
    wire \ALU.bZ0Z_11 ;
    wire \ALU.bZ0Z_12 ;
    wire \CONTROL.gZ0Z3 ;
    wire \ALU.lshift_15_0_sx_1 ;
    wire bus_14;
    wire \ALU.lshift_15_0_1_cascade_ ;
    wire \ALU.a_15_m0_sx_14 ;
    wire \ALU.lshift_15_0_1 ;
    wire \ALU.mult_1_cascade_ ;
    wire \ALU.a_15_m3_d_ns_1_1 ;
    wire \ALU.d_RNIJOQE21Z0Z_0 ;
    wire g_5;
    wire \ALU.cZ0Z_5 ;
    wire \ALU.eZ0Z_5 ;
    wire \ALU.aZ0Z_5 ;
    wire \ALU.c_RNI8KVQZ0Z_5 ;
    wire \ALU.e_RNI48JMZ0Z_5_cascade_ ;
    wire \ALU.operand2_7_ns_1_5_cascade_ ;
    wire \ALU.operand2_5 ;
    wire f_5;
    wire \ALU.bZ0Z_5 ;
    wire \ALU.b_RNI7HSPZ0Z_5 ;
    wire h_5;
    wire \ALU.dZ0Z_5 ;
    wire \ALU.d_RNIBT8EZ0Z_5 ;
    wire \INVCONTROL.operand2_2_rep1_neC_net ;
    wire \PROM.ROMDATA.m407_cascade_ ;
    wire \PROM.ROMDATA.m488_ns_cascade_ ;
    wire \INVCONTROL.operand2_fast_ne_1C_net ;
    wire \CONTROL.aluReadBus_1_sqmuxa ;
    wire \ALU.un14_log_a0_2Z0Z_15 ;
    wire \ALU.d_RNIN8NU4Z0Z_9 ;
    wire \ALU.combOperand2_0_0_9 ;
    wire DROM_ROMDATA_dintern_9ro;
    wire gpuOut_c_9;
    wire D9_in_c;
    wire \CONTROL.N_170_cascade_ ;
    wire N_186;
    wire \CONTROL.N_202 ;
    wire N_186_cascade_;
    wire bus_9;
    wire \CONTROL.ctrlOut_9 ;
    wire \INVCONTROL.dout_9C_net ;
    wire \PROM.ROMDATA.m284 ;
    wire \PROM.ROMDATA.dintern_12dfltZ0Z_0 ;
    wire \PROM.ROMDATA.m284_cascade_ ;
    wire controlWord_12_cascade_;
    wire \CONTROL.increment28lto5_0 ;
    wire \PROM.ROMDATA.m273 ;
    wire \PROM.ROMDATA.m273_cascade_ ;
    wire PROM_ROMDATA_dintern_11ro_cascade_;
    wire \CONTROL.increment28lto5_0_xZ0Z1 ;
    wire \CONTROL.increment28lto5_0_xZ0Z0 ;
    wire PROM_ROMDATA_dintern_11ro;
    wire aluStatus_4;
    wire controlWord_12;
    wire \CONTROL.g0_1_i_a6Z0Z_0 ;
    wire \CONTROL.g0_1_i_a6Z0Z_1 ;
    wire \CONTROL.g0_3_i_a7Z0Z_0 ;
    wire \PROM.ROMDATA.m271_1 ;
    wire \PROM.ROMDATA.m271_1_cascade_ ;
    wire \PROM.ROMDATA.m258_ns ;
    wire \PROM.ROMDATA.m258_ns_cascade_ ;
    wire PROM_ROMDATA_dintern_9ro_cascade_;
    wire \CONTROL.increment28lto5_1Z0Z_0 ;
    wire \PROM.ROMDATA.N_566_mux ;
    wire \PROM.ROMDATA.m470_bm ;
    wire \CONTROL.N_215 ;
    wire \CONTROL.N_86_0_cascade_ ;
    wire controlWord_1;
    wire \CONTROL.N_135 ;
    wire \CONTROL.N_74_0 ;
    wire \CONTROL.N_249 ;
    wire controlWord_5;
    wire \CONTROL.N_74_0_cascade_ ;
    wire controlWord_6;
    wire \CONTROL.un1_busState96_1_i_i_232_1_cascade_ ;
    wire \CONTROL.programCounter_ret_36_RNINU4NARZ0Z_7 ;
    wire \PROM.ROMDATA.m23_cascade_ ;
    wire PROM_ROMDATA_dintern_31_0__N_556_mux;
    wire \PROM.ROMDATA.m294_am ;
    wire \PROM.ROMDATA.m31 ;
    wire m125_e_cascade_;
    wire \PROM.ROMDATA.N_557_mux ;
    wire \PROM.ROMDATA.m77 ;
    wire m93_ns;
    wire m93_ns_cascade_;
    wire \CONTROL.addrstack_5 ;
    wire \CONTROL.addrstack_reto_5 ;
    wire \CONTROL.programCounter_1_5 ;
    wire \CONTROL.programCounter_1_reto_5 ;
    wire \CONTROL.un1_programCounter9_reto_rep1 ;
    wire \CONTROL.g0_2Z0Z_1 ;
    wire \CONTROL.N_133_0_0 ;
    wire \CONTROL.N_114_i ;
    wire \CONTROL.g1_1_4 ;
    wire \CONTROL.un1_busState114_2_0_0 ;
    wire \CONTROL.g1_1_cascade_ ;
    wire \CONTROL.addrstackptr_N_7_i ;
    wire \CONTROL.g1_0_0 ;
    wire \CONTROL.g0_i_m2_1 ;
    wire \CONTROL.addrstack_1_7 ;
    wire \CONTROL.g0_4Z0Z_2 ;
    wire \CONTROL.g0_i_m2_1_cascade_ ;
    wire \CONTROL.g1_1 ;
    wire \CONTROL.addrstackptrZ0Z_7 ;
    wire \INVCONTROL.increment_0C_net ;
    wire PROM_ROMDATA_dintern_5ro;
    wire \CONTROL.g0_2_iZ0Z_1 ;
    wire \PROM.ROMDATA.m381_am ;
    wire \PROM.ROMDATA.m375_am ;
    wire \PROM.ROMDATA.m382_ns_1 ;
    wire \ALU.rshift_3_ns_1_0 ;
    wire \ALU.N_858_cascade_ ;
    wire \ALU.rshift_15_ns_1_0_cascade_ ;
    wire \ALU.rshift_3_ns_1_4_cascade_ ;
    wire \ALU.N_862 ;
    wire \ALU.N_862_cascade_ ;
    wire \ALU.N_922_cascade_ ;
    wire \ALU.d_RNIR6J013Z0Z_2 ;
    wire \ALU.d_RNI1AHUF8Z0Z_2 ;
    wire \ALU.mult_25_10 ;
    wire \ALU.mult_11_10 ;
    wire \ALU.mult_293_c_RNIOCJMDZ0Z9 ;
    wire bfn_19_9_0_;
    wire \ALU.mult_11_11 ;
    wire \ALU.mult_21_11 ;
    wire \ALU.mult_21_c10 ;
    wire \ALU.mult_21_12 ;
    wire \ALU.mult_21_c11 ;
    wire \ALU.mult_21_13 ;
    wire \ALU.mult_21_c12 ;
    wire \ALU.mult_21_14 ;
    wire \ALU.mult_21_c13 ;
    wire \ALU.mult_23_15 ;
    wire \ALU.mult_21_c14 ;
    wire \ALU.mult_476_c_RNIFLP0OZ0Z7 ;
    wire \ALU.N_836 ;
    wire \ALU.mult_293_c_RNOZ0 ;
    wire bfn_19_10_0_;
    wire \ALU.d_RNI34ECOZ0Z_9 ;
    wire \ALU.d_RNI0PI3E1Z0Z_8 ;
    wire \ALU.mult_9_10 ;
    wire \ALU.mult_9_c9 ;
    wire \ALU.d_RNIFCNKLZ0Z_9 ;
    wire \ALU.d_RNIDR5C61Z0Z_8 ;
    wire \ALU.mult_9_11 ;
    wire \ALU.mult_9_c10 ;
    wire \ALU.d_RNIG61LGZ0Z_9 ;
    wire \ALU.mult_9_12 ;
    wire \ALU.mult_9_c11 ;
    wire \ALU.d_RNI68LSHZ0Z_9 ;
    wire \ALU.mult_9_13 ;
    wire \ALU.mult_9_c12 ;
    wire \ALU.d_RNISSV4IZ0Z_9 ;
    wire \ALU.d_RNI371041Z0Z_8 ;
    wire \ALU.mult_9_14 ;
    wire \ALU.mult_9_c13 ;
    wire \ALU.c_RNI0QV651Z0Z_10 ;
    wire \ALU.mult_9_c14 ;
    wire \ALU.mult_323_c_RNIAA0BZ0Z82 ;
    wire \ALU.d_RNIGD2441Z0Z_8 ;
    wire \ALU.N_639_cascade_ ;
    wire \ALU.d_RNIC6EBM2Z0Z_2 ;
    wire \ALU.d_RNIFVCT15Z0Z_8_cascade_ ;
    wire \ALU.lshift_11 ;
    wire \ALU.N_851 ;
    wire \ALU.N_851_cascade_ ;
    wire \ALU.c_RNINT9PO2_0Z0Z_10 ;
    wire \ALU.N_978 ;
    wire \ALU.N_978_cascade_ ;
    wire \ALU.addsub_axb_1_1 ;
    wire \ALU.N_1026 ;
    wire \ALU.mult_293_c_RNOZ0Z_0 ;
    wire \ALU.N_1011 ;
    wire \ALU.N_852_cascade_ ;
    wire \ALU.N_966 ;
    wire \ALU.N_766_cascade_ ;
    wire \ALU.N_634 ;
    wire \ALU.N_634_cascade_ ;
    wire \ALU.N_811_cascade_ ;
    wire \ALU.d_RNIK8M6K5Z0Z_6 ;
    wire \ALU.a_15_sZ0Z_11 ;
    wire \ALU.d_RNIK8M6K5Z0Z_6_cascade_ ;
    wire \ALU.mult_489_c_RNI1J3GCUZ0 ;
    wire \ALU.aZ0Z_6 ;
    wire \ALU.N_766 ;
    wire \ALU.N_606_cascade_ ;
    wire \ALU.N_606 ;
    wire \ALU.N_638 ;
    wire \ALU.a_15_m0_amZ0Z_2 ;
    wire \ALU.a_15_m1_9_cascade_ ;
    wire \ALU.aZ0Z_9 ;
    wire N_227_0;
    wire N_179;
    wire bus_2;
    wire \ALU.bZ0Z_4 ;
    wire \ALU.b_RNI5FSPZ0Z_4 ;
    wire \ALU.c_RNIHV2SZ0Z_9 ;
    wire h_4;
    wire \ALU.dZ0Z_4 ;
    wire \ALU.d_RNI9R8EZ0Z_4 ;
    wire aluOperand2_2;
    wire \ALU.N_1252_cascade_ ;
    wire \ALU.N_1204 ;
    wire \ALU.d_RNIO5IF4Z0Z_7_cascade_ ;
    wire \ALU.combOperand2_d_bmZ0Z_7 ;
    wire \ALU.d_RNIM3JB6Z0Z_7_cascade_ ;
    wire \ALU.dout_3_ns_1_7_cascade_ ;
    wire \ALU.operand2_6_ns_1_7 ;
    wire aluOperand2_2_rep1;
    wire \ALU.operand2_3_ns_1_7 ;
    wire aluOperand1_1_rep1;
    wire h_7;
    wire \ALU.dout_6_ns_1_7_cascade_ ;
    wire \ALU.N_1140_cascade_ ;
    wire \ALU.N_1092 ;
    wire DROM_ROMDATA_dintern_7ro;
    wire aluOut_7_cascade_;
    wire N_200;
    wire \PROM.ROMDATA.m267_cascade_ ;
    wire \PROM.ROMDATA.m442 ;
    wire \PROM.ROMDATA.m282 ;
    wire \PROM.ROMDATA.dintern_29dfltZ0Z_1 ;
    wire \PROM.ROMDATA.m282_cascade_ ;
    wire \CONTROL.ctrlOut_13 ;
    wire \INVCONTROL.dout_13C_net ;
    wire \CONTROL.N_35 ;
    wire \PROM.ROMDATA.m444_am ;
    wire \PROM.ROMDATA.m444_bm_cascade_ ;
    wire \PROM.ROMDATA.m289 ;
    wire \PROM.ROMDATA.m418_ns_1 ;
    wire PROM_ROMDATA_dintern_19ro;
    wire PROM_ROMDATA_dintern_19ro_cascade_;
    wire controlWord_19;
    wire f_3;
    wire controlWord_19_cascade_;
    wire controlWord_20;
    wire f_4;
    wire A14_c;
    wire A4_c;
    wire A3_c;
    wire \RAM.un1_WR_105_0Z0Z_7 ;
    wire controlWord_31;
    wire A15_c;
    wire \INVCONTROL.ramAddReg_3C_net ;
    wire \PROM.ROMDATA.m266 ;
    wire \PROM.ROMDATA.m157_cascade_ ;
    wire \PROM.ROMDATA.m265_cascade_ ;
    wire \PROM.ROMDATA.m268 ;
    wire \PROM.ROMDATA.m270_bm ;
    wire \CONTROL.aluOperation_12_i_0_6 ;
    wire controlWord_3;
    wire \CONTROL.N_219 ;
    wire controlWord_2;
    wire \INVCONTROL.aluOperation_6C_net ;
    wire \PROM.ROMDATA.N_544_mux ;
    wire \PROM.ROMDATA.m258_bm ;
    wire \CONTROL.programCounter_1_1 ;
    wire \CONTROL.programCounter_ret_19_RNIT3IGZ0Z_5 ;
    wire \CONTROL.programCounter_ret_1_RNI4MHFZ0Z_5 ;
    wire \CONTROL.un1_programCounter9_reto ;
    wire progRomAddress_5_cascade_;
    wire \PROM.ROMDATA.m243_1_cascade_ ;
    wire \PROM.ROMDATA.m244_ns_1_1 ;
    wire \CONTROL.ctrlOut_0 ;
    wire \PROM.ROMDATA.m243_1 ;
    wire \PROM.ROMDATA.m260_1 ;
    wire N_417_cascade_;
    wire \CONTROL.programCounter_1_2 ;
    wire \CONTROL.programCounter_ret_1_RNI6OHFZ0Z_6 ;
    wire \CONTROL.ctrlOut_3 ;
    wire \CONTROL.programCounter_1_4 ;
    wire \PROM.ROMDATA.m215_ns_1_N_2L1_cascade_ ;
    wire \PROM.ROMDATA.m215_ns_1 ;
    wire \CONTROL.g0_3_i_a7_0_0 ;
    wire \CONTROL.addrstack_2 ;
    wire \PROM.ROMDATA.m36 ;
    wire \PROM.ROMDATA.N_526_mux_cascade_ ;
    wire \PROM.ROMDATA.m238_bm ;
    wire aluStatus_i_3;
    wire PROM_ROMDATA_dintern_10ro;
    wire \CONTROL.g0_5Z0Z_0 ;
    wire \PROM.ROMDATA.m258_am ;
    wire PROM_ROMDATA_dintern_31_0__N_555_mux;
    wire \CONTROL.ctrlOut_5 ;
    wire \CONTROL.dout_reto_5 ;
    wire \CONTROL.programCounter_ret_19_RNIV5IGZ0Z_6 ;
    wire \CONTROL.addrstack_6 ;
    wire \CONTROL.addrstack_reto_6 ;
    wire \PROM.ROMDATA.m48 ;
    wire \CONTROL.ctrlOut_6 ;
    wire \CONTROL.dout_reto_6 ;
    wire \PROM.ROMDATA.m7 ;
    wire \PROM.ROMDATA.m392_bm_cascade_ ;
    wire \PROM.ROMDATA.m392_ns_cascade_ ;
    wire \PROM.ROMDATA.m134 ;
    wire \PROM.ROMDATA.m396_bm ;
    wire \PROM.ROMDATA.m396_am_cascade_ ;
    wire \PROM.ROMDATA.m396_ns_cascade_ ;
    wire \PROM.ROMDATA.m401_ns_1 ;
    wire \PROM.ROMDATA.m401_ns ;
    wire \ALU.N_607 ;
    wire \ALU.N_767 ;
    wire \ALU.N_607_cascade_ ;
    wire \ALU.lshift_3_ns_1_11 ;
    wire \ALU.d_RNI4N3K21Z0Z_8 ;
    wire \ALU.d_RNIH8D821Z0Z_8 ;
    wire \ALU.mult_335_c_RNOZ0 ;
    wire bfn_20_10_0_;
    wire \ALU.c_RNIBQSTOZ0Z_11 ;
    wire \ALU.c_RNIG5G6F1Z0Z_10 ;
    wire \ALU.mult_11_12 ;
    wire \ALU.mult_11_c11 ;
    wire \ALU.c_RNIN266MZ0Z_11 ;
    wire \ALU.c_RNIT73F71Z0Z_10 ;
    wire \ALU.mult_11_13 ;
    wire \ALU.mult_11_c12 ;
    wire \ALU.c_RNIK31N31Z0Z_10 ;
    wire \ALU.mult_11_14 ;
    wire \ALU.mult_11_c13 ;
    wire \ALU.mult_11_c14 ;
    wire \ALU.mult_11_c14_THRU_CO ;
    wire \ALU.c_RNIOSF6HZ0Z_11 ;
    wire \ALU.mult_335_c_RNOZ0Z_0 ;
    wire \ALU.N_835_cascade_ ;
    wire \ALU.N_852 ;
    wire \ALU.rshift_7_ns_1_7_cascade_ ;
    wire \ALU.N_925_cascade_ ;
    wire \ALU.N_833 ;
    wire \ALU.N_837 ;
    wire \ALU.rshift_7_ns_1_3_cascade_ ;
    wire \ALU.N_921 ;
    wire bus_7;
    wire \ALU.N_1030 ;
    wire \ALU.c_RNI08R632Z0Z_15 ;
    wire \ALU.eZ0Z_1 ;
    wire \ALU.eZ0Z_0 ;
    wire \ALU.eZ0Z_7 ;
    wire \ALU.eZ0Z_8 ;
    wire \ALU.eZ0Z_15 ;
    wire \ALU.eZ0Z_9 ;
    wire \ALU.N_647 ;
    wire \ALU.N_643 ;
    wire \ALU.N_707 ;
    wire \ALU.addsub_cry_14_c_RNI134CV5Z0Z_0_cascade_ ;
    wire \ALU.addsub_cry_14_c_RNIKS9S5HZ0_cascade_ ;
    wire \ALU.c_RNIE4B6N4Z0Z_15 ;
    wire \ALU.a_15_1_15_cascade_ ;
    wire \ALU.aZ0Z_15 ;
    wire \ALU.N_812 ;
    wire \ALU.N_812_cascade_ ;
    wire \ALU.addsub_cry_14_c_RNI134CVZ0Z5 ;
    wire \ALU.N_635 ;
    wire \ALU.N_639 ;
    wire \ALU.cZ0Z_1 ;
    wire \ALU.cZ0Z_0 ;
    wire \ALU.cZ0Z_7 ;
    wire \ALU.cZ0Z_8 ;
    wire \ALU.cZ0Z_15 ;
    wire \ALU.cZ0Z_9 ;
    wire \ALU.log_1_7_cascade_ ;
    wire \ALU.mult_7 ;
    wire \ALU.mult_492_c_RNIQ5BZ0Z457_cascade_ ;
    wire \ALU.lshift_7 ;
    wire \ALU.mult_492_c_RNIGN2JECZ0_cascade_ ;
    wire \ALU.aZ0Z_7 ;
    wire \ALU.d_RNIO75BGZ0Z_7 ;
    wire aluOperand2_2_rep2;
    wire \ALU.c_RNI9SHFZ0Z_14 ;
    wire \ALU.a_RNI5CPUZ0Z_14_cascade_ ;
    wire aluOperand2_1;
    wire \ALU.d_RNICJCTZ0Z_14 ;
    wire \ALU.operand2_7_ns_1_14_cascade_ ;
    wire \ALU.b_RNI83KC1Z0Z_14 ;
    wire N_191;
    wire \ALU.operand2_14_cascade_ ;
    wire \ALU.d_RNINISC7Z0Z_14 ;
    wire \ALU.dout_3_ns_1_14_cascade_ ;
    wire aluOperand1_2;
    wire \ALU.dout_6_ns_1_14_cascade_ ;
    wire aluOperand1_1;
    wire \ALU.N_1099 ;
    wire \ALU.N_1147_cascade_ ;
    wire DROM_ROMDATA_dintern_14ro;
    wire aluOut_14_cascade_;
    wire N_207;
    wire \CONTROL.un1_busState114_2_0_o2_0_0 ;
    wire \CONTROL.N_361_1 ;
    wire \CONTROL.un1_busState114_2_0_0_0 ;
    wire \INVCONTROL.increment_1C_net ;
    wire \PROM.ROMDATA.m422_am ;
    wire \PROM.ROMDATA.m422_bm_cascade_ ;
    wire \PROM.ROMDATA.m381_bm ;
    wire \PROM.ROMDATA.m298_am ;
    wire \CONTROL.programCounter_1_axb_4 ;
    wire \PROM.ROMDATA.N_543_mux_2_cascade_ ;
    wire \PROM.ROMDATA.N_559_mux ;
    wire \PROM.ROMDATA.m392_am ;
    wire \PROM.ROMDATA.m163_cascade_ ;
    wire \PROM.ROMDATA.m176_x ;
    wire \PROM.ROMDATA.N_543_mux_2 ;
    wire \PROM.ROMDATA.N_569_mux ;
    wire \PROM.ROMDATA.m109_am_1_cascade_ ;
    wire \CONTROL.addrstack_0 ;
    wire N_415;
    wire N_419;
    wire \CONTROL.addrstackZ0Z_1 ;
    wire \CONTROL.dout_reto_3 ;
    wire \CONTROL.programCounter_ret_1_RNILA8IZ0Z_3_cascade_ ;
    wire \CONTROL.programCounter_ret_19_RNIEO8JZ0Z_3 ;
    wire \CONTROL.programCounter_1_reto_0 ;
    wire \CONTROL.addrstack_3 ;
    wire \PROM.ROMDATA.m30 ;
    wire \PROM.ROMDATA.m35_1 ;
    wire \PROM.ROMDATA.m35 ;
    wire \CONTROL.programCounter_1_reto_2 ;
    wire \PROM.ROMDATA.m215_ns_1_1_1_cascade_ ;
    wire \PROM.ROMDATA.m215_ns_1_1 ;
    wire \PROM.ROMDATA.m256 ;
    wire \PROM.ROMDATA.m38 ;
    wire \PROM.ROMDATA.m251 ;
    wire \PROM.ROMDATA.m253 ;
    wire \CONTROL.programCounter_1_6 ;
    wire \CONTROL.programCounter_1_reto_6 ;
    wire \PROM.ROMDATA.m51 ;
    wire \PROM.ROMDATA.m433_am ;
    wire \PROM.ROMDATA.m399_am_cascade_ ;
    wire \PROM.ROMDATA.m399_bm ;
    wire \PROM.ROMDATA.m399_ns ;
    wire \PROM.ROMDATA.m461_ns_1 ;
    wire \CONTROL.addrstack_4 ;
    wire \PROM.ROMDATA.m22 ;
    wire \PROM.ROMDATA.m451_bm_cascade_ ;
    wire \PROM.ROMDATA.m451_am ;
    wire \PROM.ROMDATA.m451_ns ;
    wire \PROM.ROMDATA.m375_bm ;
    wire \PROM.ROMDATA.m376 ;
    wire \PROM.ROMDATA.N_256_i ;
    wire \PROM.ROMDATA.m389_bm ;
    wire \PROM.ROMDATA.m389_am_cascade_ ;
    wire \PROM.ROMDATA.m389_ns ;
    wire \ALU.lshift_3_ns_1_13_cascade_ ;
    wire \ALU.N_645_cascade_ ;
    wire \ALU.N_806_1 ;
    wire \ALU.a_15_m1_am_1_13_cascade_ ;
    wire \ALU.N_611_cascade_ ;
    wire \ALU.N_609 ;
    wire \ALU.N_641 ;
    wire \ALU.N_641_cascade_ ;
    wire \ALU.N_637 ;
    wire \ALU.d_RNITG2137Z0Z_0 ;
    wire \ALU.N_765 ;
    wire \ALU.a_15_m1_am_1_9 ;
    wire \ALU.a_15_m3_d_d_0_ns_1_3 ;
    wire \ALU.d_RNILTVJG3Z0Z_3 ;
    wire \ALU.mult_555_c_RNIJF56AMZ0_cascade_ ;
    wire \ALU.aZ0Z_12 ;
    wire \ALU.N_612 ;
    wire \ALU.N_614 ;
    wire \ALU.lshift_7_ns_1_12_cascade_ ;
    wire \ALU.N_704_cascade_ ;
    wire \ALU.d_RNIGNBT49Z0Z_8 ;
    wire \ALU.d_RNIGNBT49Z0Z_8_cascade_ ;
    wire \ALU.N_18_0 ;
    wire h_8;
    wire \ALU.mult_12 ;
    wire \ALU.mult_555_c_RNI5VJUOIZ0 ;
    wire \ALU.mult_546_c_RNIG1E6IZ0Z8 ;
    wire aluStatus_0;
    wire \ALU.status_14_12_0_cascade_ ;
    wire \ALU.status_RNO_1Z0Z_0 ;
    wire \ALU.bZ0Z_1 ;
    wire \ALU.bZ0Z_0 ;
    wire \ALU.bZ0Z_7 ;
    wire \ALU.bZ0Z_8 ;
    wire \ALU.bZ0Z_9 ;
    wire \ALU.mult_9_8 ;
    wire \ALU.mult_25_8 ;
    wire \ALU.mult_495_c_RNIKOB51JZ0_cascade_ ;
    wire \ALU.aZ0Z_8 ;
    wire \ALU.lshift_15_ns_1_8 ;
    wire \ALU.N_610 ;
    wire \ALU.N_608 ;
    wire \ALU.N_640 ;
    wire \ALU.addsub_cry_7_c_RNIDLTNZ0Z71_cascade_ ;
    wire \ALU.lshift_8 ;
    wire \ALU.N_636 ;
    wire \ALU.N_794_1 ;
    wire \ALU.N_809 ;
    wire f_1;
    wire f_0;
    wire f_7;
    wire f_8;
    wire f_9;
    wire g_1;
    wire g_0;
    wire g_7;
    wire g_8;
    wire g_15;
    wire \ALU.c_RNID85GQ_0Z0Z_15_cascade_ ;
    wire \ALU.c_RNI9DCRE2Z0Z_15 ;
    wire DROM_ROMDATA_dintern_adflt;
    wire DROM_ROMDATA_dintern_15ro;
    wire busState_1;
    wire N_208_cascade_;
    wire \ALU.status_19_14_cascade_ ;
    wire N_208;
    wire busState_0;
    wire \CONTROL.bus_7_ns_1_15 ;
    wire busState_2;
    wire bus_15;
    wire \ALU.a_15_m2_d_d_sZ0Z_0 ;
    wire bus_15_cascade_;
    wire \ALU.c_RNIJI6SHZ0Z_15 ;
    wire \ALU.c_RNID85GQZ0Z_15 ;
    wire \PROM.ROMDATA.m248_ns_cascade_ ;
    wire \PROM.ROMDATA.m249 ;
    wire \PROM.ROMDATA.m359 ;
    wire \PROM.ROMDATA.m150_cascade_ ;
    wire \PROM.ROMDATA.m228_am_cascade_ ;
    wire \PROM.ROMDATA.m25 ;
    wire \PROM.ROMDATA.m280 ;
    wire \PROM.ROMDATA.m438 ;
    wire \PROM.ROMDATA.m173 ;
    wire \PROM.ROMDATA.m23 ;
    wire PROM_ROMDATA_dintern_31_0__g1;
    wire \PROM.ROMDATA.m169_cascade_ ;
    wire \PROM.ROMDATA.m270_am ;
    wire \PROM.ROMDATA.m13_cascade_ ;
    wire \PROM.ROMDATA.m188 ;
    wire \PROM.ROMDATA.m13 ;
    wire \PROM.ROMDATA.m263 ;
    wire \CONTROL.ctrlOut_1 ;
    wire \CONTROL.dout_reto_0 ;
    wire CONTROL_addrstack_reto_0;
    wire \PROM.ROMDATA.m248_ns_1 ;
    wire \CONTROL.incrementZ0Z_0 ;
    wire \CONTROL.incrementZ0Z_1 ;
    wire \PROM.ROMDATA.m284_1 ;
    wire \CONTROL.programCounter_ret_19_RNI8I8JZ0Z_0 ;
    wire \CONTROL.programCounter_ret_1_RNIF48IZ0Z_0 ;
    wire progRomAddress_0_cascade_;
    wire \PROM.ROMDATA.m72_cascade_ ;
    wire \PROM.ROMDATA.m74 ;
    wire \PROM.ROMDATA.m80_am_cascade_ ;
    wire \PROM.ROMDATA.m93_ns_1 ;
    wire \CONTROL.programCounter_ret_1_RNIJ88IZ0Z_2 ;
    wire \CONTROL.programCounter_ret_19_RNICM8JZ0Z_2 ;
    wire progRomAddress_2_cascade_;
    wire \PROM.ROMDATA.m195_am ;
    wire \PROM.ROMDATA.m196_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m179 ;
    wire \PROM.ROMDATA.m185_am ;
    wire \PROM.ROMDATA.m191_cascade_ ;
    wire \PROM.ROMDATA.m193 ;
    wire \PROM.ROMDATA.m195_bm ;
    wire \CONTROL.programCounter_1_3 ;
    wire \CONTROL.programCounter_1_reto_3 ;
    wire \PROM.ROMDATA.m92_am ;
    wire \PROM.ROMDATA.m62_cascade_ ;
    wire \PROM.ROMDATA.m53_am ;
    wire \PROM.ROMDATA.m53_bm ;
    wire \PROM.ROMDATA.m64_bm ;
    wire \PROM.ROMDATA.m65_ns_1_cascade_ ;
    wire m65_ns;
    wire \PROM.ROMDATA.m58_cascade_ ;
    wire \PROM.ROMDATA.m64_am ;
    wire \PROM.ROMDATA.m45 ;
    wire \ALU.log_1_7 ;
    wire \ALU.log_1_5 ;
    wire \ALU.log_1_11 ;
    wire \ALU.log_1_10 ;
    wire \ALU.N_22_0 ;
    wire \ALU.N_20_0 ;
    wire \ALU.status_8_10_0_cascade_ ;
    wire \ALU.status_8_13_0 ;
    wire \ALU.status_8_3_1_0 ;
    wire \ALU.log_1_15_cascade_ ;
    wire \ALU.status_8_13_1_0 ;
    wire \ALU.c_RNIV5AOKZ0Z_13_cascade_ ;
    wire \ALU.c_RNIO5N04A_0Z0Z_13_cascade_ ;
    wire \ALU.bZ0Z_13 ;
    wire \ALU.c_RNIV5AOKZ0Z_13 ;
    wire \ALU.d_RNIRFBHE9Z0Z_0 ;
    wire \ALU.log_1_4 ;
    wire \ALU.N_16_0_cascade_ ;
    wire \ALU.status_8_8_0 ;
    wire \ALU.log_1_9 ;
    wire \ALU.d_RNI7KS2IZ0Z_9 ;
    wire \ALU.eZ0Z_12 ;
    wire \ALU.eZ0Z_13 ;
    wire \ALU.eZ0Z_14 ;
    wire g_12;
    wire g_13;
    wire g_14;
    wire \ALU.a_15_ns_1_1 ;
    wire \ALU.dZ0Z_1 ;
    wire \ALU.d_RNINUGCF4Z0Z_0 ;
    wire \ALU.rshift_0 ;
    wire \ALU.dZ0Z_0 ;
    wire \ALU.a_15_m0_7 ;
    wire \ALU.mult_492_c_RNIGN2JECZ0 ;
    wire \ALU.dZ0Z_7 ;
    wire \ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ;
    wire \ALU.a_15_m3_sZ0Z_13 ;
    wire \ALU.mult_495_c_RNIKOB51JZ0 ;
    wire \ALU.dZ0Z_8 ;
    wire \ALU.mult_15 ;
    wire \ALU.a_15_1_15 ;
    wire \ALU.a_15_m1_9 ;
    wire \ALU.mult_546_c_RNIJOT4JZ0Z8 ;
    wire \ALU.dZ0Z_9 ;
    wire \ALU.N_835 ;
    wire \ALU.d_RNIPFFDD1_0Z0Z_6_cascade_ ;
    wire \ALU.N_863_cascade_ ;
    wire \ALU.d_RNIN3H0DZ0Z_3 ;
    wire \ALU.d_RNIGPBNB6Z0Z_2_cascade_ ;
    wire \ALU.a_15_m0_5 ;
    wire bus_5;
    wire \ALU.c_RNINGV0T2Z0Z_15 ;
    wire \ALU.d_RNIPFFDD1Z0Z_6 ;
    wire \ALU.status_14_0_0_cascade_ ;
    wire \ALU.status_14_5_0 ;
    wire \ALU.status_14_7_0_cascade_ ;
    wire \ALU.status_14_13_0 ;
    wire \ALU.N_979 ;
    wire \ALU.N_979_cascade_ ;
    wire \ALU.combOperand2_a0_0Z0Z_6 ;
    wire \ALU.status_RNO_22Z0Z_0 ;
    wire \ALU.status_14_6_0 ;
    wire \ALU.status_17_I_21_c_RNOZ0 ;
    wire \ALU.status_e_0_RNO_0Z0Z_2_cascade_ ;
    wire \ALU.N_570_cascade_ ;
    wire \ALU.status_e_0_RNO_1Z0Z_2 ;
    wire aluStatus_2;
    wire PROM_ROMDATA_dintern_9ro;
    wire \CONTROL.g3Z0Z_0 ;
    wire \ALU.bZ0Z_15 ;
    wire aluOperand2_fast_2;
    wire f_15;
    wire aluOperand2_fast_1;
    wire \ALU.operand2_6_ns_1_15_cascade_ ;
    wire aluOperand2_1_rep1;
    wire \ALU.dZ0Z_15 ;
    wire \ALU.dout_6_ns_1_15 ;
    wire aluOperand1_1_rep2;
    wire h_15;
    wire \ALU.N_1100 ;
    wire \ALU.N_1148_cascade_ ;
    wire aluOperand1_0;
    wire \ALU.N_1260 ;
    wire \ALU.N_1212 ;
    wire aluOperand2_0;
    wire \ALU.combOperand2_d_bmZ0Z_15 ;
    wire \ALU.c_RNI8VV95Z0Z_15_cascade_ ;
    wire \ALU.c_RNIJTKD7Z0Z_15 ;
    wire \PROM.ROMDATA.m320_bm_cascade_ ;
    wire \PROM.ROMDATA.m410_am ;
    wire \PROM.ROMDATA.m413_am_cascade_ ;
    wire \CONTROL.ctrlOut_2 ;
    wire \CONTROL.dout_reto_2 ;
    wire \CONTROL.N_136_0 ;
    wire \CONTROL.N_86_0 ;
    wire \CONTROL.N_98_0 ;
    wire controlWord_4;
    wire \PROM.ROMDATA.m320_am ;
    wire \PROM.ROMDATA.m150 ;
    wire \PROM.ROMDATA.N_558_mux ;
    wire \PROM.ROMDATA.m49_cascade_ ;
    wire \PROM.ROMDATA.m229_1 ;
    wire \PROM.ROMDATA.m228_bm_cascade_ ;
    wire \PROM.ROMDATA.m229 ;
    wire \PROM.ROMDATA.m437_ns ;
    wire \PROM.ROMDATA.m312_bm ;
    wire \PROM.ROMDATA.m312_am ;
    wire \PROM.ROMDATA.m437_ns_1 ;
    wire \PROM.ROMDATA.m11_bm ;
    wire \PROM.ROMDATA.m18_bm_cascade_ ;
    wire \PROM.ROMDATA.m11_am ;
    wire \PROM.ROMDATA.m19_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m18_am ;
    wire \PROM.ROMDATA.m19_ns ;
    wire \PROM.ROMDATA.m33 ;
    wire \CONTROL.dout_reto_1 ;
    wire \CONTROL.programCounter_1_reto_1 ;
    wire \CONTROL.programCounter_ret_1_RNIH68IZ0Z_1_cascade_ ;
    wire \CONTROL.programCounter_ret_19_RNIAK8JZ0Z_1 ;
    wire progRomAddress_1_cascade_;
    wire \PROM.ROMDATA.m55 ;
    wire \CONTROL.programCounter_1_reto_4 ;
    wire CONTROL_addrstack_reto_4;
    wire \CONTROL.programCounter11_reto_fast ;
    wire \CONTROL.un1_programCounter9_reto_fast ;
    wire \CONTROL.programCounter_ret_1_RNINC8IZ0Z_4_cascade_ ;
    wire \CONTROL.programCounter_ret_19_RNIGQ8JZ0Z_4 ;
    wire \PROM.ROMDATA.m143 ;
    wire progRomAddress_4_cascade_;
    wire \PROM.ROMDATA.m145 ;
    wire \PROM.ROMDATA.m90 ;
    wire \PROM.ROMDATA.m92_bm ;
    wire \PROM.ROMDATA.m183_cascade_ ;
    wire \PROM.ROMDATA.m185_bm ;
    wire \PROM.ROMDATA.N_525_mux_cascade_ ;
    wire \PROM.ROMDATA.i4_mux ;
    wire \PROM.ROMDATA.m103 ;
    wire \PROM.ROMDATA.m226 ;
    wire \PROM.ROMDATA.m92_am_1 ;
    wire \PROM.ROMDATA.m158 ;
    wire \PROM.ROMDATA.m158_cascade_ ;
    wire \PROM.ROMDATA.m196_ns ;
    wire PROM_ROMDATA_dintern_6ro;
    wire \CONTROL.ctrlOut_4 ;
    wire \CONTROL.dout_reto_4 ;
    wire \ALU.aluOut_i_0 ;
    wire bfn_23_7_0_;
    wire \ALU.aluOut_i_1 ;
    wire \ALU.status_19_cry_0 ;
    wire \ALU.aluOut_i_2 ;
    wire \ALU.status_19_cry_1 ;
    wire \ALU.aluOut_i_3 ;
    wire \ALU.status_19_cry_2 ;
    wire \ALU.status_19_3 ;
    wire \ALU.aluOut_i_4 ;
    wire \ALU.status_19_cry_3 ;
    wire \ALU.status_19_4 ;
    wire \ALU.aluOut_i_5 ;
    wire \ALU.status_19_cry_4 ;
    wire \ALU.status_19_5 ;
    wire \ALU.aluOut_i_6 ;
    wire \ALU.status_19_cry_5 ;
    wire \ALU.status_19_6 ;
    wire \ALU.aluOut_i_7 ;
    wire \ALU.status_19_cry_6 ;
    wire \ALU.status_19_cry_7 ;
    wire \ALU.status_19_7 ;
    wire \ALU.aluOut_i_8 ;
    wire bfn_23_8_0_;
    wire \ALU.status_19_8 ;
    wire \ALU.aluOut_i_9 ;
    wire \ALU.status_19_cry_8 ;
    wire \ALU.status_19_9 ;
    wire \ALU.aluOut_i_10 ;
    wire \ALU.status_19_cry_9 ;
    wire \ALU.status_19_10 ;
    wire \ALU.aluOut_i_11 ;
    wire \ALU.status_19_cry_10 ;
    wire \ALU.N_126 ;
    wire \ALU.aluOut_i_12 ;
    wire \ALU.status_19_cry_11 ;
    wire \ALU.N_125 ;
    wire \ALU.aluOut_i_13 ;
    wire \ALU.status_19_cry_12 ;
    wire \ALU.status_19_13 ;
    wire \ALU.aluOut_i_14 ;
    wire \ALU.status_19_cry_13 ;
    wire \ALU.aluOut_i_15 ;
    wire \ALU.status_19_cry_14 ;
    wire \ALU.status_19Z0Z_5 ;
    wire bfn_23_9_0_;
    wire aluStatus_5;
    wire \ALU.un1_a41_0 ;
    wire \ALU.aZ0Z32 ;
    wire \ALU.N_866 ;
    wire \ALU.N_967 ;
    wire \ALU.log_1_3 ;
    wire \ALU.lshift62_2 ;
    wire \ALU.mult_558_c_RNIB3E8DCZ0 ;
    wire \ALU.a_15_d_ns_1_13_cascade_ ;
    wire \ALU.mult_558_c_RNIB75F9GZ0_cascade_ ;
    wire \ALU.aZ0Z_13 ;
    wire \ALU.d_RNIJ7J1M5_0Z0Z_2 ;
    wire \ALU.a_15_m3_d_sZ0Z_8 ;
    wire bus_0_8;
    wire \ALU.a_15_m3_d_sZ0Z_8_cascade_ ;
    wire \ALU.d_RNI12L8C5Z0Z_2 ;
    wire \ALU.d_RNIJ7J1M5Z0Z_2 ;
    wire f_12;
    wire f_13;
    wire f_14;
    wire \ALU.log_1_14 ;
    wire \ALU.a_15_m0_14 ;
    wire \ALU.addsub_cry_13_c_RNIBVHEA1Z0Z_0_cascade_ ;
    wire \ALU.addsub_cry_13_c_RNIBVHEAZ0Z1 ;
    wire \ALU.addsub_cry_13_c_RNIJMTGAZ0Z5_cascade_ ;
    wire \ALU.mult_14 ;
    wire \ALU.a_15_ns_rn_0_14_cascade_ ;
    wire \ALU.aZ0Z_14 ;
    wire \ALU.a_15_sZ0Z_3 ;
    wire \ALU.a_15_m2_sZ0Z_15 ;
    wire \ALU.a_15_sm0 ;
    wire aluOperation_1;
    wire \ALU.a_15_ns_1_7 ;
    wire \ALU.mult_388_c_RNIPGN6QZ0Z7 ;
    wire \ALU.rshift_3 ;
    wire \ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ;
    wire h_3;
    wire \ALU.a_15_sZ0Z_13 ;
    wire \ALU.c_RNIO0KOKEZ0Z_10 ;
    wire \ALU.mult_549_c_RNIE7260OZ0 ;
    wire h_10;
    wire \ALU.c_RNIBN2FN8Z0Z_11 ;
    wire \ALU.mult_552_c_RNIOT7VLFZ0Z_0 ;
    wire \ALU.mult_552_c_RNIOT7VLFZ0 ;
    wire h_11;
    wire h_12;
    wire h_13;
    wire h_14;
    wire \CONTROL.addrstack_1 ;
    wire \CONTROL.addrstackptrZ0Z_4 ;
    wire \CONTROL.addrstackptrZ0Z_2 ;
    wire \CONTROL.g1_1_3 ;
    wire bfn_23_14_0_;
    wire aluOut_0;
    wire \ALU.d_RNI27KBDZ0Z_0 ;
    wire \ALU.addsub_0 ;
    wire \ALU.addsub_cry_0_c_THRU_CO ;
    wire \ALU.d_RNIIEOKOZ0Z_1 ;
    wire \ALU.addsub_1 ;
    wire \ALU.addsub_cry_0 ;
    wire \ALU.d_RNIN178LZ0Z_2 ;
    wire \ALU.addsub_2 ;
    wire \ALU.addsub_cry_1 ;
    wire aluOut_3;
    wire \ALU.d_RNI04H8GZ0Z_3 ;
    wire \ALU.addsub_3 ;
    wire \ALU.addsub_cry_2 ;
    wire aluOut_4;
    wire \ALU.d_RNI7BF7IZ0Z_4 ;
    wire \ALU.addsub_4 ;
    wire \ALU.addsub_cry_3 ;
    wire aluOut_5;
    wire \ALU.d_RNI58QFIZ0Z_5 ;
    wire \ALU.addsub_5 ;
    wire \ALU.addsub_cry_4 ;
    wire aluOut_6;
    wire \ALU.d_RNIALE3IZ0Z_6 ;
    wire \ALU.addsub_6 ;
    wire \ALU.addsub_cry_5 ;
    wire \ALU.addsub_cry_6 ;
    wire aluOut_7;
    wire \ALU.d_RNI500DGZ0Z_7 ;
    wire \ALU.addsub_7 ;
    wire bfn_23_15_0_;
    wire aluOut_8;
    wire \ALU.d_RNIAJ1KHZ0Z_8 ;
    wire \ALU.addsub_8 ;
    wire \ALU.addsub_cry_7 ;
    wire \ALU.addsub_cry_8 ;
    wire \ALU.c_RNI1QK5KZ0Z_10 ;
    wire aluOut_10;
    wire \ALU.addsub_10 ;
    wire \ALU.addsub_cry_9 ;
    wire aluOut_11;
    wire \ALU.c_RNIRRB4IZ0Z_11 ;
    wire \ALU.addsub_11 ;
    wire \ALU.addsub_cry_10 ;
    wire \ALU.c_RNITVOEKZ0Z_12 ;
    wire aluOut_12;
    wire \ALU.addsub_12 ;
    wire \ALU.addsub_cry_11 ;
    wire \ALU.c_RNIVHVMKZ0Z_13 ;
    wire aluOut_13;
    wire \ALU.addsub_13 ;
    wire \ALU.addsub_cry_12 ;
    wire \ALU.c_RNIDDGOIZ0Z_14 ;
    wire aluOut_14;
    wire \ALU.addsub_14 ;
    wire \ALU.addsub_cry_13 ;
    wire \ALU.addsub_cry_14 ;
    wire \ALU.c_RNI0NMSHZ0Z_15 ;
    wire aluOut_15;
    wire \ALU.addsub_15 ;
    wire bfn_23_16_0_;
    wire aluStatus_1;
    wire \ALU.addsub_cry_15 ;
    wire \ALU.N_545 ;
    wire bus_6;
    wire \ALU.c_RNIPBAG72Z0Z_14 ;
    wire aluParams_0;
    wire \ALU.combOperand2_0_9 ;
    wire aluOut_9;
    wire \ALU.d_RNI70I1IZ0Z_9 ;
    wire \ALU.N_980 ;
    wire \ALU.N_1029 ;
    wire \PROM.ROMDATA.m500_ns_1 ;
    wire \PROM.ROMDATA.m500_ns ;
    wire \PROM.ROMDATA.m498_bm ;
    wire \PROM.ROMDATA.m498_am_cascade_ ;
    wire \PROM.ROMDATA.m498_ns ;
    wire \PROM.ROMDATA.m317_am ;
    wire \PROM.ROMDATA.m317_bm_cascade_ ;
    wire \PROM.ROMDATA.m312_ns ;
    wire \PROM.ROMDATA.m317_ns_cascade_ ;
    wire \PROM.ROMDATA.m325_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m320_ns ;
    wire \PROM.ROMDATA.m325_ns ;
    wire PROM_ROMDATA_dintern_14ro_cascade_;
    wire \PROM.ROMDATA.m494_ns ;
    wire \PROM.ROMDATA.m414_ns_1 ;
    wire \PROM.ROMDATA.m413_bm ;
    wire \PROM.ROMDATA.m414_ns ;
    wire \PROM.ROMDATA.m304 ;
    wire PROM_ROMDATA_dintern_13ro_cascade_;
    wire \INVCONTROL.results_1C_net ;
    wire \PROM.ROMDATA.m198 ;
    wire \PROM.ROMDATA.m16 ;
    wire \CONTROL.N_45_0 ;
    wire PROM_ROMDATA_dintern_15ro_cascade_;
    wire \INVCONTROL.results_2C_net ;
    wire \PROM.ROMDATA.m139 ;
    wire \PROM.ROMDATA.N_564_mux ;
    wire \PROM.ROMDATA.m298_bm ;
    wire \PROM.ROMDATA.N_72_i ;
    wire \PROM.ROMDATA.N_565_mux ;
    wire \PROM.ROMDATA.m287_cascade_ ;
    wire \PROM.ROMDATA.m410_bm ;
    wire \PROM.ROMDATA.m66 ;
    wire \PROM.ROMDATA.m163 ;
    wire \PROM.ROMDATA.m490 ;
    wire \PROM.ROMDATA.m149 ;
    wire \PROM.ROMDATA.m118 ;
    wire \PROM.ROMDATA.m117 ;
    wire \PROM.ROMDATA.m157 ;
    wire \PROM.ROMDATA.m456_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m456_ns ;
    wire N_418;
    wire CONTROL_addrstack_reto_3;
    wire \PROM.ROMDATA.m166_e ;
    wire \PROM.ROMDATA.m104_ns_1 ;
    wire \PROM.ROMDATA.m107 ;
    wire \PROM.ROMDATA.m104_ns_cascade_ ;
    wire \PROM.ROMDATA.m109_am ;
    wire \PROM.ROMDATA.m109_bm_cascade_ ;
    wire \PROM.ROMDATA.m121_ns ;
    wire \PROM.ROMDATA.m114 ;
    wire \PROM.ROMDATA.m111 ;
    wire \PROM.ROMDATA.m120_am_cascade_ ;
    wire \PROM.ROMDATA.m120_bm ;
    wire \PROM.ROMDATA.m121_ns_1 ;
    wire \PROM.ROMDATA.m140 ;
    wire \PROM.ROMDATA.m138_cascade_ ;
    wire \PROM.ROMDATA.m80_bm_1_cascade_ ;
    wire \PROM.ROMDATA.m80_bm ;
    wire N_417;
    wire CONTROL_addrstack_reto_2;
    wire CONTROL_programCounter11_reto_rep2;
    wire \PROM.ROMDATA.m135 ;
    wire \PROM.ROMDATA.m132 ;
    wire \PROM.ROMDATA.m83 ;
    wire \PROM.ROMDATA.m83_cascade_ ;
    wire \PROM.ROMDATA.m133 ;
    wire \PROM.ROMDATA.m161 ;
    wire \PROM.ROMDATA.m15 ;
    wire \PROM.ROMDATA.m171_ns_cascade_ ;
    wire \PROM.ROMDATA.m162 ;
    wire \PROM.ROMDATA.m172 ;
    wire \PROM.ROMDATA.m20 ;
    wire \PROM.ROMDATA.m156 ;
    wire \PROM.ROMDATA.m171_bm ;
    wire \PROM.ROMDATA.m383_cascade_ ;
    wire \PROM.ROMDATA.m427_bm ;
    wire \PROM.ROMDATA.m427_am_cascade_ ;
    wire \PROM.ROMDATA.m427_ns ;
    wire \PROM.ROMDATA.m492_am ;
    wire \PROM.ROMDATA.m492_bm ;
    wire \PROM.ROMDATA.m494_ns_1 ;
    wire \PROM.ROMDATA.m88 ;
    wire \PROM.ROMDATA.m514_ns_1 ;
    wire \PROM.ROMDATA.m181_cascade_ ;
    wire \PROM.ROMDATA.m514_ns ;
    wire \PROM.ROMDATA.N_525_mux ;
    wire \PROM.ROMDATA.m164 ;
    wire \PROM.ROMDATA.m171_am ;
    wire \ALU.dZ0Z_12 ;
    wire \ALU.dZ0Z_13 ;
    wire \ALU.dZ0Z_14 ;
    wire \ALU.c_RNIBRG4Q9Z0Z_12 ;
    wire \ALU.c_RNIBRG4Q9_0Z0Z_12 ;
    wire \ALU.mult_555_c_RNIJF56AMZ0 ;
    wire \ALU.cZ0Z_12 ;
    wire \ALU.c_RNIO5N04A_0Z0Z_13 ;
    wire \ALU.c_RNIO5N04AZ0Z_13 ;
    wire \ALU.mult_558_c_RNIB75F9GZ0 ;
    wire \ALU.cZ0Z_13 ;
    wire \ALU.cZ0Z_14 ;
    wire aluOperation_0;
    wire \ALU.a_15_d_sZ0Z_10 ;
    wire \ALU.addsub_9 ;
    wire \ALU.a_15_d_ns_sx_9 ;
    wire \ALU.status_19 ;
    wire aluOut_2;
    wire \ALU.status_19_0 ;
    wire aluOut_1;
    wire \ALU.d_RNIMGKJC1_0Z0Z_2 ;
    wire \ALU.d_RNIMGKJC1Z0Z_2_cascade_ ;
    wire \ALU.N_831 ;
    wire \ALU.N_863 ;
    wire \ALU.N_859_cascade_ ;
    wire \ALU.rshift_15_ns_1_1_cascade_ ;
    wire \ALU.a_15_m2_sZ0Z_1 ;
    wire \ALU.rshift_1_cascade_ ;
    wire bus_1;
    wire \ALU.c_RNI98D92DZ0Z_15 ;
    wire \ALU.status_19_1 ;
    wire \ALU.N_968 ;
    wire \ALU.status_19_2 ;
    wire \ALU.N_867 ;
    wire \ALU.c_RNICBIG85Z0Z_15 ;
    wire \ALU.a_15_ns_snZ0Z_14 ;
    wire \ALU.lshift_14 ;
    wire \ALU.a_15_ns_rn_0_14 ;
    wire \ALU.bZ0Z_14 ;
    wire \ALU.un1_a41_8_0 ;
    wire \ALU.un1_a41_4_0 ;
    wire \ALU.un1_operation_5_0 ;
    wire aluOperation_5;
    wire \ALU.un1_operation_10_0_cascade_ ;
    wire \ALU.un1_a41_7_0_2 ;
    wire \ALU.un1_operation_13Z0Z_2_cascade_ ;
    wire \ALU.un1_a41_4_0_2 ;
    wire \ALU.un1_a41_4_0_2_cascade_ ;
    wire \ALU.un1_a41_6_0 ;
    wire aluOperation_2;
    wire aluOperation_4;
    wire aluOperation_3;
    wire \ALU.a32Z0Z_0 ;
    wire \ALU.un1_operationZ0Z_7 ;
    wire \ALU.un1_a41_2_0 ;
    wire \PROM.ROMDATA.m160 ;
    wire aluOperation_6;
    wire aluResults_0;
    wire \ALU.un1_a41_3_0_1_cascade_ ;
    wire \ALU.un1_a41_5_0 ;
    wire \ALU.un1_a41_7_0 ;
    wire \ALU.un1_operation_13Z0Z_2 ;
    wire \ALU.un1_operation_10_0 ;
    wire aluReadBus;
    wire \ALU.un1_operation_13_0_cascade_ ;
    wire \ALU.un1_a41_9_0 ;
    wire \ALU.un1_a41_3_0_1 ;
    wire \ALU.un1_operation_13_0 ;
    wire \ALU.un1_a41_3_0 ;
    wire aluResults_2;
    wire aluResults_1;
    wire \ALU.un1_a41_2Z0Z_1 ;
    wire controlWord_22;
    wire \CONTROL.un1_busState101_3_0_0_0 ;
    wire f_6;
    wire \CONTROL.un1_busState101_3_0Z0Z_1 ;
    wire A6_c;
    wire \INVCONTROL.ramAddReg_6C_net ;
    wire \CONTROL.N_60 ;
    wire \PROM.ROMDATA.m281_cascade_ ;
    wire \PROM.ROMDATA.m60 ;
    wire \CONTROL.programCounter_1_7 ;
    wire \CONTROL.programCounter_1_reto_7 ;
    wire CLK_c_g;
    wire \PROM.ROMDATA.m181 ;
    wire \PROM.ROMDATA.m480_bm ;
    wire \PROM.ROMDATA.m480_am_cascade_ ;
    wire \PROM.ROMDATA.N_551_mux ;
    wire progRomAddress_7;
    wire \PROM.ROMDATA.m480_ns_cascade_ ;
    wire PROM_ROMDATA_dintern_25ro;
    wire g_9;
    wire PROM_ROMDATA_dintern_adflt;
    wire PROM_ROMDATA_dintern_25ro_cascade_;
    wire PROM_ROMDATA_dintern_3ro;
    wire CONTROL_romAddReg_7_9;
    wire \PROM.ROMDATA.m446_bm ;
    wire \PROM.ROMDATA.m447_ns_1 ;
    wire \PROM.ROMDATA.m446_am ;
    wire \PROM.ROMDATA.m447_ns ;
    wire \PROM.ROMDATA.m488_ns_1 ;
    wire m125_e;
    wire \PROM.ROMDATA.N_570_mux ;
    wire \PROM.ROMDATA.m2 ;
    wire \PROM.ROMDATA.m493_am ;
    wire CONTROL_addrstack_reto_1;
    wire CONTROL_programCounter11_reto;
    wire N_416;
    wire \PROM.ROMDATA.m1 ;
    wire \PROM.ROMDATA.m493_bm ;
    wire \PROM.ROMDATA.m361_am ;
    wire \PROM.ROMDATA.m211_ns_N_2L1 ;
    wire \PROM.ROMDATA.m211_ns_cascade_ ;
    wire \PROM.ROMDATA.m221cf0_1 ;
    wire \PROM.ROMDATA.m211_ns ;
    wire \PROM.ROMDATA.m221cf1_1 ;
    wire \PROM.ROMDATA.m369 ;
    wire \PROM.ROMDATA.m373 ;
    wire \PROM.ROMDATA.m298_ns ;
    wire \PROM.ROMDATA.m303_ns ;
    wire \PROM.ROMDATA.m262 ;
    wire \PROM.ROMDATA.m422_ns ;
    wire \PROM.ROMDATA.m424 ;
    wire \PROM.ROMDATA.m361_bm ;
    wire \PROM.ROMDATA.m127 ;
    wire \PROM.ROMDATA.m128 ;
    wire \PROM.ROMDATA.m137_am_cascade_ ;
    wire \PROM.ROMDATA.m137_bm ;
    wire \PROM.ROMDATA.m147_am ;
    wire \PROM.ROMDATA.m147_bm ;
    wire \PROM.ROMDATA.m148_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m148_ns ;
    wire \PROM.ROMDATA.m292 ;
    wire \PROM.ROMDATA.m299 ;
    wire \PROM.ROMDATA.m301 ;
    wire \PROM.ROMDATA.m357_bm ;
    wire \PROM.ROMDATA.m357_am_cascade_ ;
    wire \PROM.ROMDATA.m178 ;
    wire \PROM.ROMDATA.m287 ;
    wire \PROM.ROMDATA.m294_ns ;
    wire \PROM.ROMDATA.m290_cascade_ ;
    wire \PROM.ROMDATA.m303_ns_1 ;
    wire \PROM.ROMDATA.m361_ns ;
    wire \PROM.ROMDATA.m357_ns ;
    wire \PROM.ROMDATA.m363_ns ;
    wire \PROM.ROMDATA.m353_am_cascade_ ;
    wire \PROM.ROMDATA.m353_bm ;
    wire \PROM.ROMDATA.m353_ns_cascade_ ;
    wire \PROM.ROMDATA.m363_ns_1 ;
    wire \PROM.ROMDATA.m347 ;
    wire \PROM.ROMDATA.m112 ;
    wire \PROM.ROMDATA.m349_am ;
    wire \PROM.ROMDATA.m349_bm_cascade_ ;
    wire \PROM.ROMDATA.m349_ns ;
    wire \PROM.ROMDATA.m331_bm_cascade_ ;
    wire \PROM.ROMDATA.m323_bm ;
    wire \PROM.ROMDATA.m323_am_cascade_ ;
    wire \PROM.ROMDATA.m323_ns ;
    wire aluParams_1;
    wire \ALU.un14_log_0_0_15 ;
    wire \ALU.status_19_14 ;
    wire \ALU.N_586 ;
    wire \PROM.ROMDATA.m331_am ;
    wire \PROM.ROMDATA.m331_ns ;
    wire progRomAddress_5;
    wire progRomAddress_6;
    wire \PROM.ROMDATA.m343_ns_1_cascade_ ;
    wire \PROM.ROMDATA.m343_ns ;
    wire \PROM.ROMDATA.m4 ;
    wire \PROM.ROMDATA.N_28_i ;
    wire \PROM.ROMDATA.m183 ;
    wire \PROM.ROMDATA.m334_ns_1_cascade_ ;
    wire \PROM.ROMDATA.i3_mux_0 ;
    wire progRomAddress_1;
    wire progRomAddress_2;
    wire progRomAddress_0;
    wire \PROM.ROMDATA.m338_bm ;
    wire \PROM.ROMDATA.m338_am_cascade_ ;
    wire \PROM.ROMDATA.m338_ns ;
    wire \PROM.ROMDATA.m246 ;
    wire progRomAddress_4;
    wire \PROM.ROMDATA.m341_ns_1 ;
    wire progRomAddress_3;
    wire \PROM.ROMDATA.m341_ns ;
    wire _gnd_net_;

    defparam \DROM.ROMDATA.dintern_0_0_physical .WRITE_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_0_physical .READ_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_F=256'b0001000100010001000000000000000100010001000100010000000000000001000100000000000100000001000000010000000000010000000000010001000000010001000000010001000100010001000100010001000000010000000000010001000100010000000000000001000000000001000000010001000100010001;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_E=256'b0001000100010000000000000000000100010001000100000001000100010001000100010001000000010001000100010001000100010001000000010001000000010001000100010000000000000000000000000000000000010001000100010001000000010001000000010000000000010001000100010001000100010001;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_D=256'b0000000000000000000100000000000000000000000000010001000100010001000000000000000100010001000100010000000100000000000100010001000100010001000000010000000100000001000100010001000000000001000000010000000100000001000100010001000100000001000000010000000100000001;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_C=256'b0001000100010001000100010001000000000000000000010001000100010001000000000000000100000000000000010001000100010000000100000001000000000001000000010001000100010001000100010001000000000001000000010001000100010000000000010001000000000001000000010001000100010000;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_B=256'b0000000000010001000000010000000100000000010001010000000101000100010100000001010001100000000000010011000000010000001100000001010000110000010100000000010001000101000100000001000000000101000000000100000000000000000101000001010000000100000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_A=256'b0001010000010000010001000100000000010001000101010000000100000001000001010001010100010101000100010100000100000101000100010101000100000000000100010000000101000101000100000000000100010101010001010100010101000001010100010001010001010000010001010000000101000001;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_9=256'b0100010101010101000101010101010100000001000000000100000101010001000101000001010001000101000000010000000000000001010001000001010001000001000001010001000001000101010000000100000000010001000100010000010000010100000101010101000100000000000001010101000100010000;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_8=256'b0000000000010001000001010100010001010100010001000100010001000000000000000000000001000000000001000000000101000100000001010000010001000001010001000100010001000000000100000000000000000000000000000100010101000100010101010101010000000001000000000000000100000001;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_7=256'b0010001000110010001000110010001100100010001000100001000100010010000000000010001100000000001000010001001100010000001000000010001000000000000000100000000000010001001000000010001000010001000000000000000100010011001100010011001100000010000100000000001100100000;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_6=256'b0011001000100001001000010010000100110011001100010011000000010000000100110011000100010000001100000011001100010001000000000011000100100010001000000010001000010001001000100010000000100011001100010010000000000000001000100010000000100010001000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_5=256'b0011001100110001000100010011000100110011001100110001000100110001001000000010000100110011001100010001001100010001000000000010000100010001001100010011001100010001001000100010000100010001001100010011001100010001001000100000000100010001001100010011001100110001;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_4=256'b0010001000000001000100010011000100110011000100010010001000000001000100010011000100110011001100010010001000100001001100110011000100110011001100010000000000000001001100110011001100010001000100110000000000100001001100110001000100110011001100110010001000000011;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_3=256'b0001000100010001000100010001000100000000000000010011001100010011000100010001000101100010000000010101000100110001011100110011001101100010001000010011000100110001001100110001000100000010000000110011001100110001000100110001000100000010001000010011000100110001;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_2=256'b0011001100010001001000100010001100010001001100010011001100010001000000000010000100010001001100010011001100010001001000100000000100010001001100010011001100110011001000100000000100010011001100010011000100110001000000000000000100010001001100010001000100010011;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_1=256'b0000000000000001000100010001000100010001000100010000000000100001000100010001001100010001001100010010001000100011000100010001001100010001000100110010000000000001000100110001000100010001001100010000000000000011000100010001001100110011001100110000000000100011;
    defparam \DROM.ROMDATA.dintern_0_0_physical .INIT_0=256'b0001001100010011001100010001001100000000001000110011001100010001000100010011001100100000001000110001001100010001001100010011001100100010001000110011001100010001001100110011001100000010001000110011000100010001000100110011001100100010001000110001000100010001;
    SB_RAM40_4K \DROM.ROMDATA.dintern_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,\DROM.ROMDATA.dintern_0_0_NEW_3 ,dangling_wire_2,dangling_wire_3,dangling_wire_4,\DROM.ROMDATA.dintern_0_0_NEW_2 ,dangling_wire_5,dangling_wire_6,dangling_wire_7,\DROM.ROMDATA.dintern_0_0_NEW_1 ,dangling_wire_8,dangling_wire_9,dangling_wire_10,\DROM.ROMDATA.dintern_0_0_NEW_0 ,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__71657,N__26564,N__26639,N__26606,N__26369,N__26537,N__26399,N__26432,N__33233,N__33293}),
            .WADDR({dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23}),
            .MASK({dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39}),
            .WDATA({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55}),
            .RCLKE(N__28122),
            .RCLK(\INVDROM.ROMDATA.dintern_0_0RCLKN_net ),
            .RE(N__32495),
            .WCLKE(N__35927),
            .WCLK(GNDG0),
            .WE());
    defparam \DROM.ROMDATA.dintern_0_1_physical .WRITE_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_1_physical .READ_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000010010001000000001000000100000000100100010000000000010000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000001;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_E=256'b0000000000000000000000000000000100000000000000000000000000000001000000000000000000100010001000010000000000100001001000100010000000100010001000010010001000000001001000000000000100000000000000010000000000000001000000000000000000000000000000010000000000000000;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_D=256'b0000000000000001000000000000000000000000000000010000000000000001000000000000000100100010001000110010000000000010001000100010001100100010001000110010001000100001001000100000000000000000000000000000000000000000000000000000000100000000000000010000000000000001;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_C=256'b0000000000000001000000000000000000000000000000010000000000000001000000000000000100100010001000110010000000000010001000100010001000000010001000110010001000100001001000100000000100000000000000000000000000000001000000000000000100000000000000010000000000000000;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_B=256'b0000000000000000000000000000000100000100010001000000010001000000000001000100000000000110011000110010011001000100000001100110001000100100011001100010011001100011001000100110000000000100010001000000010001000100000001000100000000000100010001010000000001000000;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_A=256'b0000010001000000000001000100000000000100010000000000000001000001000001000100000100100110011001110010010001000011001001100110011100000110011001100010011001100100001000100100000100000100010000010000010001000001000001000100000100000100010000000000010001000101;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_9=256'b0000010001000001000001000100010100000000010000000000000001000000000001000100000000100110011000010000010001100101001001100110000100100110011000010010011001000101000000000100000000000000010000010000010001000000000001000100010000000100010000010000010001000001;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_8=256'b0000000001000000000001000100010000000100010000010000010001000000000000000100000100100110001000000000000001100100011001100010000001100010011000000010011001000000000000000100000000000000010000010100010001000100010001000100010000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_7=256'b0000000000000010000000000000001000000000000000100000000000000000000000000000000100000000000000010000000000000000000000000000001000000000000000100000000000000000000000000000001000000000000000010000000000000011000000000000001000000000000000010000000000000010;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_6=256'b0000000000000010000000000000001000000000000000110000000000100000000000000000000100000000000000100000000000000001000000000000001000000000000000100000000000000010000000000000001000000000000000010000000000000010000000000000000000000000000000100000000000000010;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_5=256'b0000000000000001000000000000001100000000000000110000000000000001000000000000000100000000010000110100010001000011000000000100000101000100010000010100010000000011010001000010001101000000000000110100000000000001010000000000000100000000000000110000000000100011;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_4=256'b0000000000000001000000000000001101000100000000010100010000000011010001000000000101000000000001110100010001000111010000000000010101000100010001110100010001000011010001000100001101000100010000110100010000000011010001000000000101000100000000110000000000000011;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_3=256'b0000000000100001000000000000001101000100000000010100010000000011010001000000000101000100000000110100010001000101010001000000001101000100010001110100010001100101010001000100010100000100010000010000010001000011010001000000000101000100000000110000000000000011;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_2=256'b0000000000000001000000000000001100000000000000110100000000000001010000000000001101000000000001110100010001000101010000000000010101000100010001110100010001000011010001000100001101000100000000110100010000000011010000000000000100000000000000010000000000000001;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_1=256'b0000000000000011000000000000001100000000000000110000000000000001000000000000000100000000010000010100010001000011000000000100001101000100010000110100010000000001010000000000000100000000000000010000000000000011000000000000001100000000000000110000000000000011;
    defparam \DROM.ROMDATA.dintern_0_1_physical .INIT_0=256'b0000000000000011000000000000001100000000000000010000000000000011000000000000000100000100010000110100010001000001000001000100001101000100010000110100010000000001010000000000001100000000000000010000000000000011000000000000000100000000000000110000000000000011;
    SB_RAM40_4K \DROM.ROMDATA.dintern_0_1_physical  (
            .RDATA({dangling_wire_56,dangling_wire_57,\DROM.ROMDATA.dintern_0_1_NEW_3 ,dangling_wire_58,dangling_wire_59,dangling_wire_60,\DROM.ROMDATA.dintern_0_1_NEW_2 ,dangling_wire_61,dangling_wire_62,dangling_wire_63,\DROM.ROMDATA.dintern_0_1_NEW_1 ,dangling_wire_64,dangling_wire_65,dangling_wire_66,\DROM.ROMDATA.dintern_0_1_NEW_0 ,dangling_wire_67}),
            .RADDR({dangling_wire_68,N__71651,N__26558,N__26633,N__26600,N__26363,N__26531,N__26393,N__26426,N__33227,N__33287}),
            .WADDR({dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79}),
            .MASK({dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .WDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111}),
            .RCLKE(N__28112),
            .RCLK(\INVDROM.ROMDATA.dintern_0_1RCLKN_net ),
            .RE(N__32513),
            .WCLKE(N__35928),
            .WCLK(GNDG0),
            .WE());
    defparam \DROM.ROMDATA.dintern_0_2_physical .WRITE_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_2_physical .READ_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000010001000100010001000100010000000100010001000100010001000100010000000100010001000100010001000000010001000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000001000100010001000100010001000100010001000100000000000100010000000100010001000000010001000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000010001000100010000000100010001000100010000000000010001000100010001000000010001000000000001000100000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000010000000000000001000100000000000100010001000000010001000100010001000100000000000100010001000100010000000100010001000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000010001000000000001000100010000000100010001000100000001000100010000000100010000000000010001000100010001000000010001000100000001000100000000000000010000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000010000000000000001000100000000000100010001000100000001000100010000000100000001000100000001000000010000000100010001000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000100010001000100010001000100010001000100010001000100000000000100000001000100010000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001000100010001000100010000000100110001000100010001000100110010000100110000000100010001000000010001000100000001000100000010001000100010000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000010000000000000001000100000001000100010001000100010001000100010001000100010001000100010001000100010001000100000001000100010000000000010001000000000000000100000000000000010000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000100000001000100010001000100010001000100010001000000010001000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000010000000000000001000100000000000100010000000100010001000100010001000100010001000100010001000100000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000100000000000000010001000000010001000100000001000100010001000100010001000100010001000100010001000100010000000000000000000000000001000000000000000100000000000000010000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000100010000000100010001000000010001000100010001000100010001000100010001000100010001000100000000000100010000000000010001000000010001000000000001000100000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_2_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000010001000100010001000100000001000100010001000100010001000100000000000100010000000100010001000100010001000000010001000000000000000000000000000000000000000000;
    SB_RAM40_4K \DROM.ROMDATA.dintern_0_2_physical  (
            .RDATA({dangling_wire_112,dangling_wire_113,\DROM.ROMDATA.dintern_0_2_NEW_3 ,dangling_wire_114,dangling_wire_115,dangling_wire_116,\DROM.ROMDATA.dintern_0_2_NEW_2 ,dangling_wire_117,dangling_wire_118,dangling_wire_119,\DROM.ROMDATA.dintern_0_2_NEW_1 ,dangling_wire_120,dangling_wire_121,dangling_wire_122,\DROM.ROMDATA.dintern_0_2_NEW_0 ,dangling_wire_123}),
            .RADDR({dangling_wire_124,N__71645,N__26552,N__26627,N__26594,N__26357,N__26525,N__26387,N__26420,N__33221,N__33281}),
            .WADDR({dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .MASK({dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151}),
            .WDATA({dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167}),
            .RCLKE(N__28123),
            .RCLK(\INVDROM.ROMDATA.dintern_0_2RCLKN_net ),
            .RE(N__32514),
            .WCLKE(N__35929),
            .WCLK(GNDG0),
            .WE());
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001000100010001000000010001000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .WRITE_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_3_physical .READ_MODE=2;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001000100000001000100000000000100010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001000100000001000100000001000000000000000100000000000100010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000001000100000000000100010001000100010001000100010000000000010001000000000000000000000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000001000100010000000100010001000000000001000100000000000000010000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000001000100000000000100010000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000010000000000010001000000000001000100000001000100000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100001000000000000000000000010001100110000000100010001000100010011000000000001000000000010001000100010000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000001000100000000000100010001000000000000000100000000000000010000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000001000100000000000100010000000000010001000000000000000100000000000000010000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000100010000000000010001000000000001000100000000000000010000000000000001000000000000000000000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000;
    defparam \DROM.ROMDATA.dintern_0_3_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000100000000000100010000000000000001000000000001000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \DROM.ROMDATA.dintern_0_3_physical  (
            .RDATA({dangling_wire_168,dangling_wire_169,\DROM.ROMDATA.dintern_0_3_NEW_3 ,dangling_wire_170,dangling_wire_171,dangling_wire_172,\DROM.ROMDATA.dintern_0_3_NEW_2 ,dangling_wire_173,dangling_wire_174,dangling_wire_175,\DROM.ROMDATA.dintern_0_3_NEW_1 ,dangling_wire_176,dangling_wire_177,dangling_wire_178,\DROM.ROMDATA.dintern_0_3_NEW_0 ,dangling_wire_179}),
            .RADDR({dangling_wire_180,N__71639,N__26546,N__26621,N__26588,N__26351,N__26519,N__26381,N__26414,N__33215,N__33275}),
            .WADDR({dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191}),
            .MASK({dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207}),
            .WDATA({dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223}),
            .RCLKE(N__28124),
            .RCLK(\INVDROM.ROMDATA.dintern_0_3RCLKN_net ),
            .RE(N__32530),
            .WCLKE(N__35930),
            .WCLK(GNDG0),
            .WE());
    defparam \CONTROL.addrstack_addrstack_0_0_physical .WRITE_MODE=0;
    defparam \CONTROL.addrstack_addrstack_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \CONTROL.addrstack_addrstack_0_0_physical  (
            .RDATA({\CONTROL.addrstack_15 ,\CONTROL.addrstack_14 ,\CONTROL.addrstack_13 ,\CONTROL.addrstack_12 ,\CONTROL.addrstack_11 ,\CONTROL.addrstack_10 ,\CONTROL.addrstack_9 ,\CONTROL.addrstack_8 ,\CONTROL.addrstack_7 ,\CONTROL.addrstack_6 ,\CONTROL.addrstack_5 ,\CONTROL.addrstack_4 ,\CONTROL.addrstack_3 ,\CONTROL.addrstack_2 ,\CONTROL.addrstackZ0Z_1 ,\CONTROL.addrstack_0 }),
            .RADDR({dangling_wire_224,dangling_wire_225,dangling_wire_226,N__41885,N__26690,N__27554,N__29663,N__34619,N__38369,N__29777,N__29765}),
            .WADDR({dangling_wire_227,dangling_wire_228,dangling_wire_229,N__42322,N__26724,N__27528,N__29700,N__34795,N__38461,N__31524,N__33797}),
            .MASK({dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245}),
            .WDATA({N__27725,N__27713,N__26657,N__33509,N__27737,N__28505,N__28481,N__33569,N__33524,N__26651,N__33620,N__33554,N__33605,N__33497,N__33539,N__33635}),
            .RCLKE(),
            .RCLK(\INVCONTROL.addrstack_addrstack_0_0RCLKN_net ),
            .RE(N__32544),
            .WCLKE(N__28367),
            .WCLK(N__73292),
            .WE(N__32563));
    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__80916),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__80918),
            .DIN(N__80917),
            .DOUT(N__80916),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__80918),
            .PADOUT(N__80917),
            .PADIN(N__80916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_15_iopad (
            .OE(N__80907),
            .DIN(N__80906),
            .DOUT(N__80905),
            .PACKAGEPIN(BUFFER_ADDRESS[15]));
    defparam BUFFER_ADDRESS_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_15_preio (
            .PADOEN(N__80907),
            .PADOUT(N__80906),
            .PADIN(N__80905),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26453),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D3_obuft_iopad (
            .OE(N__80898),
            .DIN(N__80897),
            .DOUT(N__80896),
            .PACKAGEPIN(D3));
    defparam D3_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D3_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D3_obuft_preio (
            .PADOEN(N__80898),
            .PADOUT(N__80897),
            .PADIN(N__80896),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35113),
            .DIN0(),
            .DOUT0(N__34244),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_12_iopad (
            .OE(N__80889),
            .DIN(N__80888),
            .DOUT(N__80887),
            .PACKAGEPIN(BUFFER_DATA_IN[12]));
    defparam BUFFER_DATA_IN_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_12_preio (
            .PADOEN(N__80889),
            .PADOUT(N__80888),
            .PADIN(N__80887),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_4_iopad (
            .OE(N__80880),
            .DIN(N__80879),
            .DOUT(N__80878),
            .PACKAGEPIN(BUFFER_ADDRESS[4]));
    defparam BUFFER_ADDRESS_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_4_preio (
            .PADOEN(N__80880),
            .PADOUT(N__80879),
            .PADIN(N__80878),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29312),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D10_obuft_iopad (
            .OE(N__80871),
            .DIN(N__80870),
            .DOUT(N__80869),
            .PACKAGEPIN(D10));
    defparam D10_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D10_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D10_obuft_preio (
            .PADOEN(N__80871),
            .PADOUT(N__80870),
            .PADIN(N__80869),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35050),
            .DIN0(),
            .DOUT0(N__26228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D7_obuft_iopad (
            .OE(N__80862),
            .DIN(N__80861),
            .DOUT(N__80860),
            .PACKAGEPIN(D7));
    defparam D7_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D7_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D7_obuft_preio (
            .PADOEN(N__80862),
            .PADOUT(N__80861),
            .PADIN(N__80860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35102),
            .DIN0(),
            .DOUT0(N__46043),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_2_iopad (
            .OE(N__80853),
            .DIN(N__80852),
            .DOUT(N__80851),
            .PACKAGEPIN(BUFFER_DATA_IN[2]));
    defparam BUFFER_DATA_IN_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_2_preio (
            .PADOEN(N__80853),
            .PADOUT(N__80852),
            .PADIN(N__80851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_CE_obuf_iopad (
            .OE(N__80844),
            .DIN(N__80843),
            .DOUT(N__80842),
            .PACKAGEPIN(B_CE));
    defparam B_CE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam B_CE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO B_CE_obuf_preio (
            .PADOEN(N__80844),
            .PADOUT(N__80843),
            .PADIN(N__80842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32493),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D0_obuft_iopad (
            .OE(N__80835),
            .DIN(N__80834),
            .DOUT(N__80833),
            .PACKAGEPIN(D0));
    defparam D0_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D0_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D0_obuft_preio (
            .PADOEN(N__80835),
            .PADOUT(N__80834),
            .PADIN(N__80833),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35117),
            .DIN0(),
            .DOUT0(N__37688),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_8_iopad (
            .OE(N__80826),
            .DIN(N__80825),
            .DOUT(N__80824),
            .PACKAGEPIN(BUFFER_DATA_OUT[8]));
    defparam BUFFER_DATA_OUT_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_8_preio (
            .PADOEN(N__80826),
            .PADOUT(N__80825),
            .PADIN(N__80824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26131),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D9_in_ibuf_iopad (
            .OE(N__80817),
            .DIN(N__80816),
            .DOUT(N__80815),
            .PACKAGEPIN(D9_in));
    defparam D9_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D9_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D9_in_ibuf_preio (
            .PADOEN(N__80817),
            .PADOUT(N__80816),
            .PADIN(N__80815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D9_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_13_iopad (
            .OE(N__80808),
            .DIN(N__80807),
            .DOUT(N__80806),
            .PACKAGEPIN(BUFFER_DATA_OUT[13]));
    defparam BUFFER_DATA_OUT_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_13_preio (
            .PADOEN(N__80808),
            .PADOUT(N__80807),
            .PADIN(N__80806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27235),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_8_iopad (
            .OE(N__80799),
            .DIN(N__80798),
            .DOUT(N__80797),
            .PACKAGEPIN(BUFFER_DATA_IN[8]));
    defparam BUFFER_DATA_IN_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_8_preio (
            .PADOEN(N__80799),
            .PADOUT(N__80798),
            .PADIN(N__80797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_8_iopad (
            .OE(N__80790),
            .DIN(N__80789),
            .DOUT(N__80788),
            .PACKAGEPIN(BUFFER_ADDRESS[8]));
    defparam BUFFER_ADDRESS_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_8_preio (
            .PADOEN(N__80790),
            .PADOUT(N__80789),
            .PADIN(N__80788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29234),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_12_iopad (
            .OE(N__80781),
            .DIN(N__80780),
            .DOUT(N__80779),
            .PACKAGEPIN(BUFFER_ADDRESS[12]));
    defparam BUFFER_ADDRESS_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_12_preio (
            .PADOEN(N__80781),
            .PADOUT(N__80780),
            .PADIN(N__80779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26492),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D6_obuft_iopad (
            .OE(N__80772),
            .DIN(N__80771),
            .DOUT(N__80770),
            .PACKAGEPIN(D6));
    defparam D6_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D6_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D6_obuft_preio (
            .PADOEN(N__80772),
            .PADOUT(N__80771),
            .PADIN(N__80770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35071),
            .DIN0(),
            .DOUT0(N__63380),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D10_in_ibuf_iopad (
            .OE(N__80763),
            .DIN(N__80762),
            .DOUT(N__80761),
            .PACKAGEPIN(D10_in));
    defparam D10_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D10_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D10_in_ibuf_preio (
            .PADOEN(N__80763),
            .PADOUT(N__80762),
            .PADIN(N__80761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D10_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D2_obuft_iopad (
            .OE(N__80754),
            .DIN(N__80753),
            .DOUT(N__80752),
            .PACKAGEPIN(D2));
    defparam D2_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D2_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D2_obuft_preio (
            .PADOEN(N__80754),
            .PADOUT(N__80753),
            .PADIN(N__80752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35099),
            .DIN0(),
            .DOUT0(N__43481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D4_in_ibuf_iopad (
            .OE(N__80745),
            .DIN(N__80744),
            .DOUT(N__80743),
            .PACKAGEPIN(D4_in));
    defparam D4_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D4_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D4_in_ibuf_preio (
            .PADOEN(N__80745),
            .PADOUT(N__80744),
            .PADIN(N__80743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D4_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_13_iopad (
            .OE(N__80736),
            .DIN(N__80735),
            .DOUT(N__80734),
            .PACKAGEPIN(BUFFER_DATA_IN[13]));
    defparam BUFFER_DATA_IN_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_13_preio (
            .PADOEN(N__80736),
            .PADOUT(N__80735),
            .PADIN(N__80734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_5_iopad (
            .OE(N__80727),
            .DIN(N__80726),
            .DOUT(N__80725),
            .PACKAGEPIN(BUFFER_DATA_OUT[5]));
    defparam BUFFER_DATA_OUT_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_5_preio (
            .PADOEN(N__80727),
            .PADOUT(N__80726),
            .PADIN(N__80725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__52531),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_7_iopad (
            .OE(N__80718),
            .DIN(N__80717),
            .DOUT(N__80716),
            .PACKAGEPIN(BUFFER_DATA_IN[7]));
    defparam BUFFER_DATA_IN_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_7_preio (
            .PADOEN(N__80718),
            .PADOUT(N__80717),
            .PADIN(N__80716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A4_obuf_iopad (
            .OE(N__80709),
            .DIN(N__80708),
            .DOUT(N__80707),
            .PACKAGEPIN(A4));
    defparam A4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A4_obuf_preio (
            .PADOEN(N__80709),
            .PADOUT(N__80708),
            .PADIN(N__80707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44072),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_7_iopad (
            .OE(N__80700),
            .DIN(N__80699),
            .DOUT(N__80698),
            .PACKAGEPIN(BUFFER_ADDRESS[7]));
    defparam BUFFER_ADDRESS_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_7_preio (
            .PADOEN(N__80700),
            .PADOUT(N__80699),
            .PADIN(N__80698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29252),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D0_in_ibuf_iopad (
            .OE(N__80691),
            .DIN(N__80690),
            .DOUT(N__80689),
            .PACKAGEPIN(D0_in));
    defparam D0_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D0_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D0_in_ibuf_preio (
            .PADOEN(N__80691),
            .PADOUT(N__80690),
            .PADIN(N__80689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D0_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A10_obuf_iopad (
            .OE(N__80682),
            .DIN(N__80681),
            .DOUT(N__80680),
            .PACKAGEPIN(A10));
    defparam A10_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A10_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A10_obuf_preio (
            .PADOEN(N__80682),
            .PADOUT(N__80681),
            .PADIN(N__80680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31202),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_9_iopad (
            .OE(N__80673),
            .DIN(N__80672),
            .DOUT(N__80671),
            .PACKAGEPIN(BUFFER_DATA_OUT[9]));
    defparam BUFFER_DATA_OUT_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_9_preio (
            .PADOEN(N__80673),
            .PADOUT(N__80672),
            .PADIN(N__80671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__40385),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_12_iopad (
            .OE(N__80664),
            .DIN(N__80663),
            .DOUT(N__80662),
            .PACKAGEPIN(BUFFER_DATA_OUT[12]));
    defparam BUFFER_DATA_OUT_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_12_preio (
            .PADOEN(N__80664),
            .PADOUT(N__80663),
            .PADIN(N__80662),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26320),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D3_in_ibuf_iopad (
            .OE(N__80655),
            .DIN(N__80654),
            .DOUT(N__80653),
            .PACKAGEPIN(D3_in));
    defparam D3_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D3_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D3_in_ibuf_preio (
            .PADOEN(N__80655),
            .PADOUT(N__80654),
            .PADIN(N__80653),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D3_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UB_obuf_iopad (
            .OE(N__80646),
            .DIN(N__80645),
            .DOUT(N__80644),
            .PACKAGEPIN(UB));
    defparam UB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UB_obuf_preio (
            .PADOEN(N__80646),
            .PADOUT(N__80645),
            .PADIN(N__80644),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25684),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_LB_obuf_iopad (
            .OE(N__80637),
            .DIN(N__80636),
            .DOUT(N__80635),
            .PACKAGEPIN(B_LB));
    defparam B_LB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam B_LB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO B_LB_obuf_preio (
            .PADOEN(N__80637),
            .PADOUT(N__80636),
            .PADIN(N__80635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25791),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D15_obuft_iopad (
            .OE(N__80628),
            .DIN(N__80627),
            .DOUT(N__80626),
            .PACKAGEPIN(D15));
    defparam D15_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D15_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D15_obuft_preio (
            .PADOEN(N__80628),
            .PADOUT(N__80627),
            .PADIN(N__80626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35025),
            .DIN0(),
            .DOUT0(N__49219),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_13_iopad (
            .OE(N__80619),
            .DIN(N__80618),
            .DOUT(N__80617),
            .PACKAGEPIN(BUFFER_ADDRESS[13]));
    defparam BUFFER_ADDRESS_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_13_preio (
            .PADOEN(N__80619),
            .PADOUT(N__80618),
            .PADIN(N__80617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26474),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D14_in_ibuf_iopad (
            .OE(N__80610),
            .DIN(N__80609),
            .DOUT(N__80608),
            .PACKAGEPIN(D14_in));
    defparam D14_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D14_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D14_in_ibuf_preio (
            .PADOEN(N__80610),
            .PADOUT(N__80609),
            .PADIN(N__80608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D14_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A6_obuf_iopad (
            .OE(N__80601),
            .DIN(N__80600),
            .DOUT(N__80599),
            .PACKAGEPIN(A6));
    defparam A6_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A6_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A6_obuf_preio (
            .PADOEN(N__80601),
            .PADOUT(N__80600),
            .PADIN(N__80599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__70373),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WR_obuf_iopad (
            .OE(N__80592),
            .DIN(N__80591),
            .DOUT(N__80590),
            .PACKAGEPIN(WR));
    defparam WR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WR_obuf_preio (
            .PADOEN(N__80592),
            .PADOUT(N__80591),
            .PADIN(N__80590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25672),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D13_obuft_iopad (
            .OE(N__80583),
            .DIN(N__80582),
            .DOUT(N__80581),
            .PACKAGEPIN(D13));
    defparam D13_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D13_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D13_obuft_preio (
            .PADOEN(N__80583),
            .PADOUT(N__80582),
            .PADIN(N__80581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35007),
            .DIN0(),
            .DOUT0(N__27242),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_10_iopad (
            .OE(N__80574),
            .DIN(N__80573),
            .DOUT(N__80572),
            .PACKAGEPIN(BUFFER_DATA_IN[10]));
    defparam BUFFER_DATA_IN_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_10_preio (
            .PADOEN(N__80574),
            .PADOUT(N__80573),
            .PADIN(N__80572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D11_in_ibuf_iopad (
            .OE(N__80565),
            .DIN(N__80564),
            .DOUT(N__80563),
            .PACKAGEPIN(D11_in));
    defparam D11_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D11_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D11_in_ibuf_preio (
            .PADOEN(N__80565),
            .PADOUT(N__80564),
            .PADIN(N__80563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D11_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A8_obuf_iopad (
            .OE(N__80556),
            .DIN(N__80555),
            .DOUT(N__80554),
            .PACKAGEPIN(A8));
    defparam A8_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A8_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A8_obuf_preio (
            .PADOEN(N__80556),
            .PADOUT(N__80555),
            .PADIN(N__80554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31058),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_2_iopad (
            .OE(N__80547),
            .DIN(N__80546),
            .DOUT(N__80545),
            .PACKAGEPIN(BUFFER_DATA_OUT[2]));
    defparam BUFFER_DATA_OUT_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_2_preio (
            .PADOEN(N__80547),
            .PADOUT(N__80546),
            .PADIN(N__80545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43474),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_6_iopad (
            .OE(N__80538),
            .DIN(N__80537),
            .DOUT(N__80536),
            .PACKAGEPIN(BUFFER_DATA_IN[6]));
    defparam BUFFER_DATA_IN_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_6_preio (
            .PADOEN(N__80538),
            .PADOUT(N__80537),
            .PADIN(N__80536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_6_iopad (
            .OE(N__80529),
            .DIN(N__80528),
            .DOUT(N__80527),
            .PACKAGEPIN(BUFFER_ADDRESS[6]));
    defparam BUFFER_ADDRESS_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_6_preio (
            .PADOEN(N__80529),
            .PADOUT(N__80528),
            .PADIN(N__80527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29267),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A9_obuf_iopad (
            .OE(N__80520),
            .DIN(N__80519),
            .DOUT(N__80518),
            .PACKAGEPIN(A9));
    defparam A9_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A9_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A9_obuf_preio (
            .PADOEN(N__80520),
            .PADOUT(N__80519),
            .PADIN(N__80518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31112),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LB_obuf_iopad (
            .OE(N__80511),
            .DIN(N__80510),
            .DOUT(N__80509),
            .PACKAGEPIN(LB));
    defparam LB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LB_obuf_preio (
            .PADOEN(N__80511),
            .PADOUT(N__80510),
            .PADIN(N__80509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25688),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D8_obuft_iopad (
            .OE(N__80502),
            .DIN(N__80501),
            .DOUT(N__80500),
            .PACKAGEPIN(D8));
    defparam D8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D8_obuft_preio (
            .PADOEN(N__80502),
            .PADOUT(N__80501),
            .PADIN(N__80500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35100),
            .DIN0(),
            .DOUT0(N__26138),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_11_iopad (
            .OE(N__80493),
            .DIN(N__80492),
            .DOUT(N__80491),
            .PACKAGEPIN(BUFFER_DATA_OUT[11]));
    defparam BUFFER_DATA_OUT_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_11_preio (
            .PADOEN(N__80493),
            .PADOUT(N__80492),
            .PADIN(N__80491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37354),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A7_obuf_iopad (
            .OE(N__80484),
            .DIN(N__80483),
            .DOUT(N__80482),
            .PACKAGEPIN(A7));
    defparam A7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A7_obuf_preio (
            .PADOEN(N__80484),
            .PADOUT(N__80483),
            .PADIN(N__80482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29354),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OE_obuf_iopad (
            .OE(N__80475),
            .DIN(N__80474),
            .DOUT(N__80473),
            .PACKAGEPIN(OE));
    defparam OE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam OE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO OE_obuf_preio (
            .PADOEN(N__80475),
            .PADOUT(N__80474),
            .PADIN(N__80473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25703),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO3_obuf_iopad (
            .OE(N__80466),
            .DIN(N__80465),
            .DOUT(N__80464),
            .PACKAGEPIN(GPIO3));
    defparam GPIO3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO3_obuf_preio (
            .PADOEN(N__80466),
            .PADOUT(N__80465),
            .PADIN(N__80464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25811),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_10_iopad (
            .OE(N__80457),
            .DIN(N__80456),
            .DOUT(N__80455),
            .PACKAGEPIN(BUFFER_ADDRESS[10]));
    defparam BUFFER_ADDRESS_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_10_preio (
            .PADOEN(N__80457),
            .PADOUT(N__80456),
            .PADIN(N__80455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26510),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D2_in_ibuf_iopad (
            .OE(N__80448),
            .DIN(N__80447),
            .DOUT(N__80446),
            .PACKAGEPIN(D2_in));
    defparam D2_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D2_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D2_in_ibuf_preio (
            .PADOEN(N__80448),
            .PADOUT(N__80447),
            .PADIN(N__80446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D2_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_11_iopad (
            .OE(N__80439),
            .DIN(N__80438),
            .DOUT(N__80437),
            .PACKAGEPIN(BUFFER_DATA_IN[11]));
    defparam BUFFER_DATA_IN_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_11_preio (
            .PADOEN(N__80439),
            .PADOUT(N__80438),
            .PADIN(N__80437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A14_obuf_iopad (
            .OE(N__80430),
            .DIN(N__80429),
            .DOUT(N__80428),
            .PACKAGEPIN(A14));
    defparam A14_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A14_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A14_obuf_preio (
            .PADOEN(N__80430),
            .PADOUT(N__80429),
            .PADIN(N__80428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44111),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A5_obuf_iopad (
            .OE(N__80421),
            .DIN(N__80420),
            .DOUT(N__80419),
            .PACKAGEPIN(A5));
    defparam A5_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A5_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A5_obuf_preio (
            .PADOEN(N__80421),
            .PADOUT(N__80420),
            .PADIN(N__80419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29414),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_3_iopad (
            .OE(N__80412),
            .DIN(N__80411),
            .DOUT(N__80410),
            .PACKAGEPIN(BUFFER_DATA_OUT[3]));
    defparam BUFFER_DATA_OUT_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_3_preio (
            .PADOEN(N__80412),
            .PADOUT(N__80411),
            .PADIN(N__80410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_1_iopad (
            .OE(N__80403),
            .DIN(N__80402),
            .DOUT(N__80401),
            .PACKAGEPIN(BUFFER_DATA_IN[1]));
    defparam BUFFER_DATA_IN_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_1_preio (
            .PADOEN(N__80403),
            .PADOUT(N__80402),
            .PADIN(N__80401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D9_obuft_iopad (
            .OE(N__80394),
            .DIN(N__80393),
            .DOUT(N__80392),
            .PACKAGEPIN(D9));
    defparam D9_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D9_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D9_obuft_preio (
            .PADOEN(N__80394),
            .PADOUT(N__80393),
            .PADIN(N__80392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35097),
            .DIN0(),
            .DOUT0(N__40384),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_1_iopad (
            .OE(N__80385),
            .DIN(N__80384),
            .DOUT(N__80383),
            .PACKAGEPIN(BUFFER_ADDRESS[1]));
    defparam BUFFER_ADDRESS_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_1_preio (
            .PADOEN(N__80385),
            .PADOUT(N__80384),
            .PADIN(N__80383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26159),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D11_obuft_iopad (
            .OE(N__80376),
            .DIN(N__80375),
            .DOUT(N__80374),
            .PACKAGEPIN(D11));
    defparam D11_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D11_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D11_obuft_preio (
            .PADOEN(N__80376),
            .PADOUT(N__80375),
            .PADIN(N__80374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35098),
            .DIN0(),
            .DOUT0(N__37358),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D12_in_ibuf_iopad (
            .OE(N__80367),
            .DIN(N__80366),
            .DOUT(N__80365),
            .PACKAGEPIN(D12_in));
    defparam D12_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D12_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D12_in_ibuf_preio (
            .PADOEN(N__80367),
            .PADOUT(N__80366),
            .PADIN(N__80365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D12_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A15_obuf_iopad (
            .OE(N__80358),
            .DIN(N__80357),
            .DOUT(N__80356),
            .PACKAGEPIN(A15));
    defparam A15_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A15_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A15_obuf_preio (
            .PADOEN(N__80358),
            .PADOUT(N__80357),
            .PADIN(N__80356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44978),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A13_obuf_iopad (
            .OE(N__80349),
            .DIN(N__80348),
            .DOUT(N__80347),
            .PACKAGEPIN(A13));
    defparam A13_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A13_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A13_obuf_preio (
            .PADOEN(N__80349),
            .PADOUT(N__80348),
            .PADIN(N__80347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28175),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A1_obuf_iopad (
            .OE(N__80340),
            .DIN(N__80339),
            .DOUT(N__80338),
            .PACKAGEPIN(A1));
    defparam A1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A1_obuf_preio (
            .PADOEN(N__80340),
            .PADOUT(N__80339),
            .PADIN(N__80338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31310),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_10_iopad (
            .OE(N__80331),
            .DIN(N__80330),
            .DOUT(N__80329),
            .PACKAGEPIN(BUFFER_DATA_OUT[10]));
    defparam BUFFER_DATA_OUT_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_10_preio (
            .PADOEN(N__80331),
            .PADOUT(N__80330),
            .PADIN(N__80329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26224),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_UB_obuf_iopad (
            .OE(N__80322),
            .DIN(N__80321),
            .DOUT(N__80320),
            .PACKAGEPIN(B_UB));
    defparam B_UB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam B_UB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO B_UB_obuf_preio (
            .PADOEN(N__80322),
            .PADOUT(N__80321),
            .PADIN(N__80320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25792),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D7_in_ibuf_iopad (
            .OE(N__80313),
            .DIN(N__80312),
            .DOUT(N__80311),
            .PACKAGEPIN(D7_in));
    defparam D7_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D7_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D7_in_ibuf_preio (
            .PADOEN(N__80313),
            .PADOUT(N__80312),
            .PADIN(N__80311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D7_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_WR_obuf_iopad (
            .OE(N__80304),
            .DIN(N__80303),
            .DOUT(N__80302),
            .PACKAGEPIN(B_WR));
    defparam B_WR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam B_WR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO B_WR_obuf_preio (
            .PADOEN(N__80304),
            .PADOUT(N__80303),
            .PADIN(N__80302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25793),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_14_iopad (
            .OE(N__80295),
            .DIN(N__80294),
            .DOUT(N__80293),
            .PACKAGEPIN(BUFFER_DATA_IN[14]));
    defparam BUFFER_DATA_IN_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_14_preio (
            .PADOEN(N__80295),
            .PADOUT(N__80294),
            .PADIN(N__80293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_11_iopad (
            .OE(N__80286),
            .DIN(N__80285),
            .DOUT(N__80284),
            .PACKAGEPIN(BUFFER_ADDRESS[11]));
    defparam BUFFER_ADDRESS_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_11_preio (
            .PADOEN(N__80286),
            .PADOUT(N__80285),
            .PADIN(N__80284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25748),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO11_obuf_iopad (
            .OE(N__80277),
            .DIN(N__80276),
            .DOUT(N__80275),
            .PACKAGEPIN(GPIO11));
    defparam GPIO11_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO11_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO11_obuf_preio (
            .PADOEN(N__80277),
            .PADOUT(N__80276),
            .PADIN(N__80275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_6_iopad (
            .OE(N__80268),
            .DIN(N__80267),
            .DOUT(N__80266),
            .PACKAGEPIN(BUFFER_DATA_OUT[6]));
    defparam BUFFER_DATA_OUT_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_6_preio (
            .PADOEN(N__80268),
            .PADOUT(N__80267),
            .PADIN(N__80266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__63370),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A2_obuf_iopad (
            .OE(N__80259),
            .DIN(N__80258),
            .DOUT(N__80257),
            .PACKAGEPIN(A2));
    defparam A2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A2_obuf_preio (
            .PADOEN(N__80259),
            .PADOUT(N__80258),
            .PADIN(N__80257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29576),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D5_obuft_iopad (
            .OE(N__80250),
            .DIN(N__80249),
            .DOUT(N__80248),
            .PACKAGEPIN(D5));
    defparam D5_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D5_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D5_obuft_preio (
            .PADOEN(N__80250),
            .PADOUT(N__80249),
            .PADIN(N__80248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35052),
            .DIN0(),
            .DOUT0(N__52541),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D4_obuft_iopad (
            .OE(N__80241),
            .DIN(N__80240),
            .DOUT(N__80239),
            .PACKAGEPIN(D4));
    defparam D4_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D4_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D4_obuft_preio (
            .PADOEN(N__80241),
            .PADOUT(N__80240),
            .PADIN(N__80239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35101),
            .DIN0(),
            .DOUT0(N__33764),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A3_obuf_iopad (
            .OE(N__80232),
            .DIN(N__80231),
            .DOUT(N__80230),
            .PACKAGEPIN(A3));
    defparam A3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A3_obuf_preio (
            .PADOEN(N__80232),
            .PADOUT(N__80231),
            .PADIN(N__80230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__44048),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_0_iopad (
            .OE(N__80223),
            .DIN(N__80222),
            .DOUT(N__80221),
            .PACKAGEPIN(BUFFER_DATA_OUT[0]));
    defparam BUFFER_DATA_OUT_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_0_preio (
            .PADOEN(N__80223),
            .PADOUT(N__80222),
            .PADIN(N__80221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37684),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_0_iopad (
            .OE(N__80214),
            .DIN(N__80213),
            .DOUT(N__80212),
            .PACKAGEPIN(BUFFER_DATA_IN[0]));
    defparam BUFFER_DATA_IN_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_0_preio (
            .PADOEN(N__80214),
            .PADOUT(N__80213),
            .PADIN(N__80212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_0_iopad (
            .OE(N__80205),
            .DIN(N__80204),
            .DOUT(N__80203),
            .PACKAGEPIN(BUFFER_ADDRESS[0]));
    defparam BUFFER_ADDRESS_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_0_preio (
            .PADOEN(N__80205),
            .PADOUT(N__80204),
            .PADIN(N__80203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26177),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_15_iopad (
            .OE(N__80196),
            .DIN(N__80195),
            .DOUT(N__80194),
            .PACKAGEPIN(BUFFER_DATA_OUT[15]));
    defparam BUFFER_DATA_OUT_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_15_preio (
            .PADOEN(N__80196),
            .PADOUT(N__80195),
            .PADIN(N__80194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__49232),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A11_obuf_iopad (
            .OE(N__80187),
            .DIN(N__80186),
            .DOUT(N__80185),
            .PACKAGEPIN(A11));
    defparam A11_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A11_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A11_obuf_preio (
            .PADOEN(N__80187),
            .PADOUT(N__80186),
            .PADIN(N__80185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO9_obuf_iopad (
            .OE(N__80178),
            .DIN(N__80177),
            .DOUT(N__80176),
            .PACKAGEPIN(GPIO9));
    defparam GPIO9_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO9_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO9_obuf_preio (
            .PADOEN(N__80178),
            .PADOUT(N__80177),
            .PADIN(N__80176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32573),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D5_in_ibuf_iopad (
            .OE(N__80169),
            .DIN(N__80168),
            .DOUT(N__80167),
            .PACKAGEPIN(D5_in));
    defparam D5_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D5_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D5_in_ibuf_preio (
            .PADOEN(N__80169),
            .PADOUT(N__80168),
            .PADIN(N__80167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D5_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_14_iopad (
            .OE(N__80160),
            .DIN(N__80159),
            .DOUT(N__80158),
            .PACKAGEPIN(BUFFER_ADDRESS[14]));
    defparam BUFFER_ADDRESS_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_14_preio (
            .PADOEN(N__80160),
            .PADOUT(N__80159),
            .PADIN(N__80158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25733),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D15_in_ibuf_iopad (
            .OE(N__80151),
            .DIN(N__80150),
            .DOUT(N__80149),
            .PACKAGEPIN(D15_in));
    defparam D15_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D15_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D15_in_ibuf_preio (
            .PADOEN(N__80151),
            .PADOUT(N__80150),
            .PADIN(N__80149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D15_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D1_in_ibuf_iopad (
            .OE(N__80142),
            .DIN(N__80141),
            .DOUT(N__80140),
            .PACKAGEPIN(D1_in));
    defparam D1_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D1_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D1_in_ibuf_preio (
            .PADOEN(N__80142),
            .PADOUT(N__80141),
            .PADIN(N__80140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D1_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD B_OE_obuf_iopad (
            .OE(N__80133),
            .DIN(N__80132),
            .DOUT(N__80131),
            .PACKAGEPIN(B_OE));
    defparam B_OE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam B_OE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO B_OE_obuf_preio (
            .PADOEN(N__80133),
            .PADOUT(N__80132),
            .PADIN(N__80131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25775),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_15_iopad (
            .OE(N__80124),
            .DIN(N__80123),
            .DOUT(N__80122),
            .PACKAGEPIN(BUFFER_DATA_IN[15]));
    defparam BUFFER_DATA_IN_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_15_preio (
            .PADOEN(N__80124),
            .PADOUT(N__80123),
            .PADIN(N__80122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_7_iopad (
            .OE(N__80115),
            .DIN(N__80114),
            .DOUT(N__80113),
            .PACKAGEPIN(BUFFER_DATA_OUT[7]));
    defparam BUFFER_DATA_OUT_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_7_preio (
            .PADOEN(N__80115),
            .PADOUT(N__80114),
            .PADIN(N__80113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__46039),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_5_iopad (
            .OE(N__80106),
            .DIN(N__80105),
            .DOUT(N__80104),
            .PACKAGEPIN(BUFFER_DATA_IN[5]));
    defparam BUFFER_DATA_IN_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_5_preio (
            .PADOEN(N__80106),
            .PADOUT(N__80105),
            .PADIN(N__80104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D12_obuft_iopad (
            .OE(N__80097),
            .DIN(N__80096),
            .DOUT(N__80095),
            .PACKAGEPIN(D12));
    defparam D12_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D12_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D12_obuft_preio (
            .PADOEN(N__80097),
            .PADOUT(N__80096),
            .PADIN(N__80095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35051),
            .DIN0(),
            .DOUT0(N__26327),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_5_iopad (
            .OE(N__80088),
            .DIN(N__80087),
            .DOUT(N__80086),
            .PACKAGEPIN(BUFFER_ADDRESS[5]));
    defparam BUFFER_ADDRESS_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_5_preio (
            .PADOEN(N__80088),
            .PADOUT(N__80087),
            .PADIN(N__80086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29288),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TX_obuft_iopad (
            .OE(N__80079),
            .DIN(N__80078),
            .DOUT(N__80077),
            .PACKAGEPIN(TX));
    defparam TX_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TX_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TX_obuft_preio (
            .PADOEN(N__80079),
            .PADOUT(N__80078),
            .PADIN(N__80077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D8_in_ibuf_iopad (
            .OE(N__80070),
            .DIN(N__80069),
            .DOUT(N__80068),
            .PACKAGEPIN(D8_in));
    defparam D8_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D8_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D8_in_ibuf_preio (
            .PADOEN(N__80070),
            .PADOUT(N__80069),
            .PADIN(N__80068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D8_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_1_iopad (
            .OE(N__80061),
            .DIN(N__80060),
            .DOUT(N__80059),
            .PACKAGEPIN(BUFFER_DATA_OUT[1]));
    defparam BUFFER_DATA_OUT_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_1_preio (
            .PADOEN(N__80061),
            .PADOUT(N__80060),
            .PADIN(N__80059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__69070),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D6_in_ibuf_iopad (
            .OE(N__80052),
            .DIN(N__80051),
            .DOUT(N__80050),
            .PACKAGEPIN(D6_in));
    defparam D6_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D6_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D6_in_ibuf_preio (
            .PADOEN(N__80052),
            .PADOUT(N__80051),
            .PADIN(N__80050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D6_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_3_iopad (
            .OE(N__80043),
            .DIN(N__80042),
            .DOUT(N__80041),
            .PACKAGEPIN(BUFFER_DATA_IN[3]));
    defparam BUFFER_DATA_IN_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_3_preio (
            .PADOEN(N__80043),
            .PADOUT(N__80042),
            .PADIN(N__80041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D13_in_ibuf_iopad (
            .OE(N__80034),
            .DIN(N__80033),
            .DOUT(N__80032),
            .PACKAGEPIN(D13_in));
    defparam D13_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam D13_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO D13_in_ibuf_preio (
            .PADOEN(N__80034),
            .PADOUT(N__80033),
            .PADIN(N__80032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(D13_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_3_iopad (
            .OE(N__80025),
            .DIN(N__80024),
            .DOUT(N__80023),
            .PACKAGEPIN(BUFFER_ADDRESS[3]));
    defparam BUFFER_ADDRESS_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_3_preio (
            .PADOEN(N__80025),
            .PADOUT(N__80024),
            .PADIN(N__80023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29333),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_14_iopad (
            .OE(N__80016),
            .DIN(N__80015),
            .DOUT(N__80014),
            .PACKAGEPIN(BUFFER_DATA_OUT[14]));
    defparam BUFFER_DATA_OUT_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_14_preio (
            .PADOEN(N__80016),
            .PADOUT(N__80015),
            .PADIN(N__80014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__39752),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_9_iopad (
            .OE(N__80007),
            .DIN(N__80006),
            .DOUT(N__80005),
            .PACKAGEPIN(BUFFER_DATA_IN[9]));
    defparam BUFFER_DATA_IN_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_9_preio (
            .PADOEN(N__80007),
            .PADOUT(N__80006),
            .PADIN(N__80005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_9_iopad (
            .OE(N__79998),
            .DIN(N__79997),
            .DOUT(N__79996),
            .PACKAGEPIN(BUFFER_ADDRESS[9]));
    defparam BUFFER_ADDRESS_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_9_preio (
            .PADOEN(N__79998),
            .PADOUT(N__79997),
            .PADIN(N__79996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25715),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D1_obuft_iopad (
            .OE(N__79989),
            .DIN(N__79988),
            .DOUT(N__79987),
            .PACKAGEPIN(D1));
    defparam D1_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D1_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D1_obuft_preio (
            .PADOEN(N__79989),
            .PADOUT(N__79988),
            .PADIN(N__79987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35112),
            .DIN0(),
            .DOUT0(N__69074),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A12_obuf_iopad (
            .OE(N__79980),
            .DIN(N__79979),
            .DOUT(N__79978),
            .PACKAGEPIN(A12));
    defparam A12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A12_obuf_preio (
            .PADOEN(N__79980),
            .PADOUT(N__79979),
            .PADIN(N__79978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_OUT_obuf_4_iopad (
            .OE(N__79971),
            .DIN(N__79970),
            .DOUT(N__79969),
            .PACKAGEPIN(BUFFER_DATA_OUT[4]));
    defparam BUFFER_DATA_OUT_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_OUT_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_DATA_OUT_obuf_4_preio (
            .PADOEN(N__79971),
            .PADOUT(N__79970),
            .PADIN(N__79969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33763),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_DATA_IN_ibuf_4_iopad (
            .OE(N__79962),
            .DIN(N__79961),
            .DOUT(N__79960),
            .PACKAGEPIN(BUFFER_DATA_IN[4]));
    defparam BUFFER_DATA_IN_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_DATA_IN_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO BUFFER_DATA_IN_ibuf_4_preio (
            .PADOEN(N__79962),
            .PADOUT(N__79961),
            .PADIN(N__79960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(gpuOut_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A0_obuf_iopad (
            .OE(N__79953),
            .DIN(N__79952),
            .DOUT(N__79951),
            .PACKAGEPIN(A0));
    defparam A0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam A0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO A0_obuf_preio (
            .PADOEN(N__79953),
            .PADOUT(N__79952),
            .PADIN(N__79951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31334),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CE_obuf_iopad (
            .OE(N__79944),
            .DIN(N__79943),
            .DOUT(N__79942),
            .PACKAGEPIN(CE));
    defparam CE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CE_obuf_preio (
            .PADOEN(N__79944),
            .PADOUT(N__79943),
            .PADIN(N__79942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32494),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D14_obuft_iopad (
            .OE(N__79935),
            .DIN(N__79934),
            .DOUT(N__79933),
            .PACKAGEPIN(D14));
    defparam D14_obuft_preio.NEG_TRIGGER=1'b0;
    defparam D14_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO D14_obuft_preio (
            .PADOEN(N__79935),
            .PADOUT(N__79934),
            .PADIN(N__79933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35026),
            .DIN0(),
            .DOUT0(N__39751),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFFER_ADDRESS_obuf_2_iopad (
            .OE(N__79926),
            .DIN(N__79925),
            .DOUT(N__79924),
            .PACKAGEPIN(BUFFER_ADDRESS[2]));
    defparam BUFFER_ADDRESS_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam BUFFER_ADDRESS_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFFER_ADDRESS_obuf_2_preio (
            .PADOEN(N__79926),
            .PADOUT(N__79925),
            .PADIN(N__79924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29108),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__20304 (
            .O(N__79907),
            .I(N__79904));
    LocalMux I__20303 (
            .O(N__79904),
            .I(N__79901));
    Odrv4 I__20302 (
            .O(N__79901),
            .I(\PROM.ROMDATA.m331_ns ));
    InMux I__20301 (
            .O(N__79898),
            .I(N__79892));
    InMux I__20300 (
            .O(N__79897),
            .I(N__79887));
    InMux I__20299 (
            .O(N__79896),
            .I(N__79884));
    InMux I__20298 (
            .O(N__79895),
            .I(N__79875));
    LocalMux I__20297 (
            .O(N__79892),
            .I(N__79867));
    CascadeMux I__20296 (
            .O(N__79891),
            .I(N__79863));
    CascadeMux I__20295 (
            .O(N__79890),
            .I(N__79854));
    LocalMux I__20294 (
            .O(N__79887),
            .I(N__79851));
    LocalMux I__20293 (
            .O(N__79884),
            .I(N__79847));
    InMux I__20292 (
            .O(N__79883),
            .I(N__79835));
    InMux I__20291 (
            .O(N__79882),
            .I(N__79819));
    InMux I__20290 (
            .O(N__79881),
            .I(N__79819));
    InMux I__20289 (
            .O(N__79880),
            .I(N__79819));
    InMux I__20288 (
            .O(N__79879),
            .I(N__79819));
    InMux I__20287 (
            .O(N__79878),
            .I(N__79819));
    LocalMux I__20286 (
            .O(N__79875),
            .I(N__79815));
    InMux I__20285 (
            .O(N__79874),
            .I(N__79812));
    InMux I__20284 (
            .O(N__79873),
            .I(N__79809));
    InMux I__20283 (
            .O(N__79872),
            .I(N__79801));
    InMux I__20282 (
            .O(N__79871),
            .I(N__79801));
    InMux I__20281 (
            .O(N__79870),
            .I(N__79801));
    Span4Mux_v I__20280 (
            .O(N__79867),
            .I(N__79798));
    InMux I__20279 (
            .O(N__79866),
            .I(N__79795));
    InMux I__20278 (
            .O(N__79863),
            .I(N__79792));
    InMux I__20277 (
            .O(N__79862),
            .I(N__79789));
    CascadeMux I__20276 (
            .O(N__79861),
            .I(N__79784));
    InMux I__20275 (
            .O(N__79860),
            .I(N__79778));
    InMux I__20274 (
            .O(N__79859),
            .I(N__79778));
    InMux I__20273 (
            .O(N__79858),
            .I(N__79775));
    InMux I__20272 (
            .O(N__79857),
            .I(N__79772));
    InMux I__20271 (
            .O(N__79854),
            .I(N__79769));
    Span4Mux_v I__20270 (
            .O(N__79851),
            .I(N__79766));
    InMux I__20269 (
            .O(N__79850),
            .I(N__79763));
    Span4Mux_v I__20268 (
            .O(N__79847),
            .I(N__79758));
    InMux I__20267 (
            .O(N__79846),
            .I(N__79755));
    InMux I__20266 (
            .O(N__79845),
            .I(N__79752));
    InMux I__20265 (
            .O(N__79844),
            .I(N__79748));
    InMux I__20264 (
            .O(N__79843),
            .I(N__79744));
    InMux I__20263 (
            .O(N__79842),
            .I(N__79741));
    InMux I__20262 (
            .O(N__79841),
            .I(N__79738));
    InMux I__20261 (
            .O(N__79840),
            .I(N__79735));
    InMux I__20260 (
            .O(N__79839),
            .I(N__79732));
    InMux I__20259 (
            .O(N__79838),
            .I(N__79729));
    LocalMux I__20258 (
            .O(N__79835),
            .I(N__79726));
    InMux I__20257 (
            .O(N__79834),
            .I(N__79723));
    InMux I__20256 (
            .O(N__79833),
            .I(N__79716));
    InMux I__20255 (
            .O(N__79832),
            .I(N__79716));
    InMux I__20254 (
            .O(N__79831),
            .I(N__79716));
    CascadeMux I__20253 (
            .O(N__79830),
            .I(N__79711));
    LocalMux I__20252 (
            .O(N__79819),
            .I(N__79708));
    InMux I__20251 (
            .O(N__79818),
            .I(N__79705));
    Span4Mux_v I__20250 (
            .O(N__79815),
            .I(N__79698));
    LocalMux I__20249 (
            .O(N__79812),
            .I(N__79698));
    LocalMux I__20248 (
            .O(N__79809),
            .I(N__79698));
    InMux I__20247 (
            .O(N__79808),
            .I(N__79695));
    LocalMux I__20246 (
            .O(N__79801),
            .I(N__79692));
    Sp12to4 I__20245 (
            .O(N__79798),
            .I(N__79683));
    LocalMux I__20244 (
            .O(N__79795),
            .I(N__79683));
    LocalMux I__20243 (
            .O(N__79792),
            .I(N__79683));
    LocalMux I__20242 (
            .O(N__79789),
            .I(N__79683));
    InMux I__20241 (
            .O(N__79788),
            .I(N__79678));
    InMux I__20240 (
            .O(N__79787),
            .I(N__79678));
    InMux I__20239 (
            .O(N__79784),
            .I(N__79675));
    InMux I__20238 (
            .O(N__79783),
            .I(N__79672));
    LocalMux I__20237 (
            .O(N__79778),
            .I(N__79667));
    LocalMux I__20236 (
            .O(N__79775),
            .I(N__79667));
    LocalMux I__20235 (
            .O(N__79772),
            .I(N__79662));
    LocalMux I__20234 (
            .O(N__79769),
            .I(N__79662));
    Span4Mux_h I__20233 (
            .O(N__79766),
            .I(N__79657));
    LocalMux I__20232 (
            .O(N__79763),
            .I(N__79657));
    InMux I__20231 (
            .O(N__79762),
            .I(N__79652));
    InMux I__20230 (
            .O(N__79761),
            .I(N__79652));
    Span4Mux_h I__20229 (
            .O(N__79758),
            .I(N__79649));
    LocalMux I__20228 (
            .O(N__79755),
            .I(N__79644));
    LocalMux I__20227 (
            .O(N__79752),
            .I(N__79644));
    InMux I__20226 (
            .O(N__79751),
            .I(N__79641));
    LocalMux I__20225 (
            .O(N__79748),
            .I(N__79638));
    InMux I__20224 (
            .O(N__79747),
            .I(N__79635));
    LocalMux I__20223 (
            .O(N__79744),
            .I(N__79628));
    LocalMux I__20222 (
            .O(N__79741),
            .I(N__79628));
    LocalMux I__20221 (
            .O(N__79738),
            .I(N__79628));
    LocalMux I__20220 (
            .O(N__79735),
            .I(N__79621));
    LocalMux I__20219 (
            .O(N__79732),
            .I(N__79621));
    LocalMux I__20218 (
            .O(N__79729),
            .I(N__79621));
    Span4Mux_v I__20217 (
            .O(N__79726),
            .I(N__79614));
    LocalMux I__20216 (
            .O(N__79723),
            .I(N__79614));
    LocalMux I__20215 (
            .O(N__79716),
            .I(N__79614));
    InMux I__20214 (
            .O(N__79715),
            .I(N__79610));
    InMux I__20213 (
            .O(N__79714),
            .I(N__79605));
    InMux I__20212 (
            .O(N__79711),
            .I(N__79605));
    Span4Mux_v I__20211 (
            .O(N__79708),
            .I(N__79598));
    LocalMux I__20210 (
            .O(N__79705),
            .I(N__79598));
    Span4Mux_h I__20209 (
            .O(N__79698),
            .I(N__79598));
    LocalMux I__20208 (
            .O(N__79695),
            .I(N__79591));
    Span12Mux_h I__20207 (
            .O(N__79692),
            .I(N__79591));
    Span12Mux_h I__20206 (
            .O(N__79683),
            .I(N__79591));
    LocalMux I__20205 (
            .O(N__79678),
            .I(N__79584));
    LocalMux I__20204 (
            .O(N__79675),
            .I(N__79584));
    LocalMux I__20203 (
            .O(N__79672),
            .I(N__79584));
    Span12Mux_s11_v I__20202 (
            .O(N__79667),
            .I(N__79581));
    Span4Mux_v I__20201 (
            .O(N__79662),
            .I(N__79578));
    Span4Mux_v I__20200 (
            .O(N__79657),
            .I(N__79573));
    LocalMux I__20199 (
            .O(N__79652),
            .I(N__79573));
    Span4Mux_h I__20198 (
            .O(N__79649),
            .I(N__79556));
    Span4Mux_v I__20197 (
            .O(N__79644),
            .I(N__79556));
    LocalMux I__20196 (
            .O(N__79641),
            .I(N__79556));
    Span4Mux_v I__20195 (
            .O(N__79638),
            .I(N__79556));
    LocalMux I__20194 (
            .O(N__79635),
            .I(N__79556));
    Span4Mux_v I__20193 (
            .O(N__79628),
            .I(N__79556));
    Span4Mux_v I__20192 (
            .O(N__79621),
            .I(N__79556));
    Span4Mux_h I__20191 (
            .O(N__79614),
            .I(N__79556));
    InMux I__20190 (
            .O(N__79613),
            .I(N__79553));
    LocalMux I__20189 (
            .O(N__79610),
            .I(progRomAddress_5));
    LocalMux I__20188 (
            .O(N__79605),
            .I(progRomAddress_5));
    Odrv4 I__20187 (
            .O(N__79598),
            .I(progRomAddress_5));
    Odrv12 I__20186 (
            .O(N__79591),
            .I(progRomAddress_5));
    Odrv4 I__20185 (
            .O(N__79584),
            .I(progRomAddress_5));
    Odrv12 I__20184 (
            .O(N__79581),
            .I(progRomAddress_5));
    Odrv4 I__20183 (
            .O(N__79578),
            .I(progRomAddress_5));
    Odrv4 I__20182 (
            .O(N__79573),
            .I(progRomAddress_5));
    Odrv4 I__20181 (
            .O(N__79556),
            .I(progRomAddress_5));
    LocalMux I__20180 (
            .O(N__79553),
            .I(progRomAddress_5));
    CascadeMux I__20179 (
            .O(N__79532),
            .I(N__79524));
    CascadeMux I__20178 (
            .O(N__79531),
            .I(N__79519));
    CascadeMux I__20177 (
            .O(N__79530),
            .I(N__79516));
    CascadeMux I__20176 (
            .O(N__79529),
            .I(N__79511));
    CascadeMux I__20175 (
            .O(N__79528),
            .I(N__79508));
    CascadeMux I__20174 (
            .O(N__79527),
            .I(N__79504));
    InMux I__20173 (
            .O(N__79524),
            .I(N__79490));
    InMux I__20172 (
            .O(N__79523),
            .I(N__79490));
    InMux I__20171 (
            .O(N__79522),
            .I(N__79483));
    InMux I__20170 (
            .O(N__79519),
            .I(N__79474));
    InMux I__20169 (
            .O(N__79516),
            .I(N__79474));
    InMux I__20168 (
            .O(N__79515),
            .I(N__79474));
    InMux I__20167 (
            .O(N__79514),
            .I(N__79474));
    InMux I__20166 (
            .O(N__79511),
            .I(N__79469));
    InMux I__20165 (
            .O(N__79508),
            .I(N__79469));
    InMux I__20164 (
            .O(N__79507),
            .I(N__79464));
    InMux I__20163 (
            .O(N__79504),
            .I(N__79464));
    InMux I__20162 (
            .O(N__79503),
            .I(N__79461));
    InMux I__20161 (
            .O(N__79502),
            .I(N__79458));
    InMux I__20160 (
            .O(N__79501),
            .I(N__79447));
    InMux I__20159 (
            .O(N__79500),
            .I(N__79447));
    InMux I__20158 (
            .O(N__79499),
            .I(N__79440));
    InMux I__20157 (
            .O(N__79498),
            .I(N__79440));
    InMux I__20156 (
            .O(N__79497),
            .I(N__79440));
    CascadeMux I__20155 (
            .O(N__79496),
            .I(N__79437));
    CascadeMux I__20154 (
            .O(N__79495),
            .I(N__79434));
    LocalMux I__20153 (
            .O(N__79490),
            .I(N__79428));
    CascadeMux I__20152 (
            .O(N__79489),
            .I(N__79425));
    CascadeMux I__20151 (
            .O(N__79488),
            .I(N__79422));
    InMux I__20150 (
            .O(N__79487),
            .I(N__79408));
    InMux I__20149 (
            .O(N__79486),
            .I(N__79405));
    LocalMux I__20148 (
            .O(N__79483),
            .I(N__79398));
    LocalMux I__20147 (
            .O(N__79474),
            .I(N__79398));
    LocalMux I__20146 (
            .O(N__79469),
            .I(N__79398));
    LocalMux I__20145 (
            .O(N__79464),
            .I(N__79395));
    LocalMux I__20144 (
            .O(N__79461),
            .I(N__79392));
    LocalMux I__20143 (
            .O(N__79458),
            .I(N__79388));
    InMux I__20142 (
            .O(N__79457),
            .I(N__79381));
    InMux I__20141 (
            .O(N__79456),
            .I(N__79381));
    InMux I__20140 (
            .O(N__79455),
            .I(N__79381));
    InMux I__20139 (
            .O(N__79454),
            .I(N__79378));
    InMux I__20138 (
            .O(N__79453),
            .I(N__79373));
    InMux I__20137 (
            .O(N__79452),
            .I(N__79373));
    LocalMux I__20136 (
            .O(N__79447),
            .I(N__79370));
    LocalMux I__20135 (
            .O(N__79440),
            .I(N__79367));
    InMux I__20134 (
            .O(N__79437),
            .I(N__79358));
    InMux I__20133 (
            .O(N__79434),
            .I(N__79358));
    InMux I__20132 (
            .O(N__79433),
            .I(N__79358));
    InMux I__20131 (
            .O(N__79432),
            .I(N__79358));
    InMux I__20130 (
            .O(N__79431),
            .I(N__79355));
    Span4Mux_v I__20129 (
            .O(N__79428),
            .I(N__79352));
    InMux I__20128 (
            .O(N__79425),
            .I(N__79343));
    InMux I__20127 (
            .O(N__79422),
            .I(N__79343));
    InMux I__20126 (
            .O(N__79421),
            .I(N__79343));
    InMux I__20125 (
            .O(N__79420),
            .I(N__79343));
    InMux I__20124 (
            .O(N__79419),
            .I(N__79336));
    InMux I__20123 (
            .O(N__79418),
            .I(N__79336));
    CascadeMux I__20122 (
            .O(N__79417),
            .I(N__79333));
    InMux I__20121 (
            .O(N__79416),
            .I(N__79328));
    InMux I__20120 (
            .O(N__79415),
            .I(N__79328));
    CascadeMux I__20119 (
            .O(N__79414),
            .I(N__79324));
    CascadeMux I__20118 (
            .O(N__79413),
            .I(N__79315));
    InMux I__20117 (
            .O(N__79412),
            .I(N__79309));
    InMux I__20116 (
            .O(N__79411),
            .I(N__79309));
    LocalMux I__20115 (
            .O(N__79408),
            .I(N__79306));
    LocalMux I__20114 (
            .O(N__79405),
            .I(N__79301));
    Span4Mux_v I__20113 (
            .O(N__79398),
            .I(N__79301));
    Span4Mux_v I__20112 (
            .O(N__79395),
            .I(N__79294));
    Span4Mux_v I__20111 (
            .O(N__79392),
            .I(N__79290));
    InMux I__20110 (
            .O(N__79391),
            .I(N__79287));
    Span4Mux_h I__20109 (
            .O(N__79388),
            .I(N__79277));
    LocalMux I__20108 (
            .O(N__79381),
            .I(N__79277));
    LocalMux I__20107 (
            .O(N__79378),
            .I(N__79277));
    LocalMux I__20106 (
            .O(N__79373),
            .I(N__79277));
    Span4Mux_v I__20105 (
            .O(N__79370),
            .I(N__79274));
    Span4Mux_h I__20104 (
            .O(N__79367),
            .I(N__79269));
    LocalMux I__20103 (
            .O(N__79358),
            .I(N__79269));
    LocalMux I__20102 (
            .O(N__79355),
            .I(N__79262));
    Span4Mux_h I__20101 (
            .O(N__79352),
            .I(N__79262));
    LocalMux I__20100 (
            .O(N__79343),
            .I(N__79262));
    InMux I__20099 (
            .O(N__79342),
            .I(N__79259));
    InMux I__20098 (
            .O(N__79341),
            .I(N__79256));
    LocalMux I__20097 (
            .O(N__79336),
            .I(N__79253));
    InMux I__20096 (
            .O(N__79333),
            .I(N__79250));
    LocalMux I__20095 (
            .O(N__79328),
            .I(N__79245));
    InMux I__20094 (
            .O(N__79327),
            .I(N__79238));
    InMux I__20093 (
            .O(N__79324),
            .I(N__79238));
    InMux I__20092 (
            .O(N__79323),
            .I(N__79238));
    InMux I__20091 (
            .O(N__79322),
            .I(N__79233));
    InMux I__20090 (
            .O(N__79321),
            .I(N__79233));
    InMux I__20089 (
            .O(N__79320),
            .I(N__79228));
    InMux I__20088 (
            .O(N__79319),
            .I(N__79228));
    InMux I__20087 (
            .O(N__79318),
            .I(N__79223));
    InMux I__20086 (
            .O(N__79315),
            .I(N__79223));
    InMux I__20085 (
            .O(N__79314),
            .I(N__79220));
    LocalMux I__20084 (
            .O(N__79309),
            .I(N__79217));
    Span4Mux_v I__20083 (
            .O(N__79306),
            .I(N__79214));
    Span4Mux_h I__20082 (
            .O(N__79301),
            .I(N__79211));
    InMux I__20081 (
            .O(N__79300),
            .I(N__79204));
    InMux I__20080 (
            .O(N__79299),
            .I(N__79201));
    InMux I__20079 (
            .O(N__79298),
            .I(N__79196));
    InMux I__20078 (
            .O(N__79297),
            .I(N__79196));
    Span4Mux_h I__20077 (
            .O(N__79294),
            .I(N__79193));
    InMux I__20076 (
            .O(N__79293),
            .I(N__79190));
    Span4Mux_h I__20075 (
            .O(N__79290),
            .I(N__79185));
    LocalMux I__20074 (
            .O(N__79287),
            .I(N__79185));
    InMux I__20073 (
            .O(N__79286),
            .I(N__79182));
    Span4Mux_v I__20072 (
            .O(N__79277),
            .I(N__79179));
    Span4Mux_h I__20071 (
            .O(N__79274),
            .I(N__79176));
    Span4Mux_h I__20070 (
            .O(N__79269),
            .I(N__79171));
    Span4Mux_h I__20069 (
            .O(N__79262),
            .I(N__79171));
    LocalMux I__20068 (
            .O(N__79259),
            .I(N__79162));
    LocalMux I__20067 (
            .O(N__79256),
            .I(N__79162));
    Span4Mux_h I__20066 (
            .O(N__79253),
            .I(N__79162));
    LocalMux I__20065 (
            .O(N__79250),
            .I(N__79162));
    InMux I__20064 (
            .O(N__79249),
            .I(N__79157));
    InMux I__20063 (
            .O(N__79248),
            .I(N__79157));
    Span4Mux_v I__20062 (
            .O(N__79245),
            .I(N__79150));
    LocalMux I__20061 (
            .O(N__79238),
            .I(N__79150));
    LocalMux I__20060 (
            .O(N__79233),
            .I(N__79150));
    LocalMux I__20059 (
            .O(N__79228),
            .I(N__79143));
    LocalMux I__20058 (
            .O(N__79223),
            .I(N__79143));
    LocalMux I__20057 (
            .O(N__79220),
            .I(N__79143));
    Span4Mux_v I__20056 (
            .O(N__79217),
            .I(N__79139));
    Span4Mux_h I__20055 (
            .O(N__79214),
            .I(N__79134));
    Span4Mux_h I__20054 (
            .O(N__79211),
            .I(N__79134));
    InMux I__20053 (
            .O(N__79210),
            .I(N__79131));
    InMux I__20052 (
            .O(N__79209),
            .I(N__79126));
    InMux I__20051 (
            .O(N__79208),
            .I(N__79126));
    InMux I__20050 (
            .O(N__79207),
            .I(N__79123));
    LocalMux I__20049 (
            .O(N__79204),
            .I(N__79116));
    LocalMux I__20048 (
            .O(N__79201),
            .I(N__79116));
    LocalMux I__20047 (
            .O(N__79196),
            .I(N__79116));
    Span4Mux_h I__20046 (
            .O(N__79193),
            .I(N__79111));
    LocalMux I__20045 (
            .O(N__79190),
            .I(N__79111));
    Span4Mux_v I__20044 (
            .O(N__79185),
            .I(N__79104));
    LocalMux I__20043 (
            .O(N__79182),
            .I(N__79104));
    Span4Mux_h I__20042 (
            .O(N__79179),
            .I(N__79104));
    Span4Mux_h I__20041 (
            .O(N__79176),
            .I(N__79091));
    Span4Mux_v I__20040 (
            .O(N__79171),
            .I(N__79091));
    Span4Mux_v I__20039 (
            .O(N__79162),
            .I(N__79091));
    LocalMux I__20038 (
            .O(N__79157),
            .I(N__79091));
    Span4Mux_h I__20037 (
            .O(N__79150),
            .I(N__79091));
    Span4Mux_v I__20036 (
            .O(N__79143),
            .I(N__79091));
    InMux I__20035 (
            .O(N__79142),
            .I(N__79088));
    Odrv4 I__20034 (
            .O(N__79139),
            .I(progRomAddress_6));
    Odrv4 I__20033 (
            .O(N__79134),
            .I(progRomAddress_6));
    LocalMux I__20032 (
            .O(N__79131),
            .I(progRomAddress_6));
    LocalMux I__20031 (
            .O(N__79126),
            .I(progRomAddress_6));
    LocalMux I__20030 (
            .O(N__79123),
            .I(progRomAddress_6));
    Odrv4 I__20029 (
            .O(N__79116),
            .I(progRomAddress_6));
    Odrv4 I__20028 (
            .O(N__79111),
            .I(progRomAddress_6));
    Odrv4 I__20027 (
            .O(N__79104),
            .I(progRomAddress_6));
    Odrv4 I__20026 (
            .O(N__79091),
            .I(progRomAddress_6));
    LocalMux I__20025 (
            .O(N__79088),
            .I(progRomAddress_6));
    CascadeMux I__20024 (
            .O(N__79067),
            .I(\PROM.ROMDATA.m343_ns_1_cascade_ ));
    CascadeMux I__20023 (
            .O(N__79064),
            .I(N__79061));
    InMux I__20022 (
            .O(N__79061),
            .I(N__79058));
    LocalMux I__20021 (
            .O(N__79058),
            .I(N__79055));
    Span4Mux_h I__20020 (
            .O(N__79055),
            .I(N__79052));
    Odrv4 I__20019 (
            .O(N__79052),
            .I(\PROM.ROMDATA.m343_ns ));
    CascadeMux I__20018 (
            .O(N__79049),
            .I(N__79045));
    CascadeMux I__20017 (
            .O(N__79048),
            .I(N__79040));
    InMux I__20016 (
            .O(N__79045),
            .I(N__79037));
    InMux I__20015 (
            .O(N__79044),
            .I(N__79034));
    CascadeMux I__20014 (
            .O(N__79043),
            .I(N__79030));
    InMux I__20013 (
            .O(N__79040),
            .I(N__79027));
    LocalMux I__20012 (
            .O(N__79037),
            .I(N__79024));
    LocalMux I__20011 (
            .O(N__79034),
            .I(N__79021));
    InMux I__20010 (
            .O(N__79033),
            .I(N__79016));
    InMux I__20009 (
            .O(N__79030),
            .I(N__79016));
    LocalMux I__20008 (
            .O(N__79027),
            .I(N__79011));
    Span4Mux_h I__20007 (
            .O(N__79024),
            .I(N__79011));
    Span4Mux_v I__20006 (
            .O(N__79021),
            .I(N__79006));
    LocalMux I__20005 (
            .O(N__79016),
            .I(N__79006));
    Span4Mux_v I__20004 (
            .O(N__79011),
            .I(N__79001));
    Span4Mux_h I__20003 (
            .O(N__79006),
            .I(N__79001));
    Odrv4 I__20002 (
            .O(N__79001),
            .I(\PROM.ROMDATA.m4 ));
    InMux I__20001 (
            .O(N__78998),
            .I(N__78990));
    InMux I__20000 (
            .O(N__78997),
            .I(N__78985));
    InMux I__19999 (
            .O(N__78996),
            .I(N__78981));
    InMux I__19998 (
            .O(N__78995),
            .I(N__78977));
    InMux I__19997 (
            .O(N__78994),
            .I(N__78972));
    InMux I__19996 (
            .O(N__78993),
            .I(N__78972));
    LocalMux I__19995 (
            .O(N__78990),
            .I(N__78969));
    InMux I__19994 (
            .O(N__78989),
            .I(N__78966));
    InMux I__19993 (
            .O(N__78988),
            .I(N__78963));
    LocalMux I__19992 (
            .O(N__78985),
            .I(N__78960));
    InMux I__19991 (
            .O(N__78984),
            .I(N__78957));
    LocalMux I__19990 (
            .O(N__78981),
            .I(N__78952));
    InMux I__19989 (
            .O(N__78980),
            .I(N__78949));
    LocalMux I__19988 (
            .O(N__78977),
            .I(N__78944));
    LocalMux I__19987 (
            .O(N__78972),
            .I(N__78944));
    Span4Mux_v I__19986 (
            .O(N__78969),
            .I(N__78940));
    LocalMux I__19985 (
            .O(N__78966),
            .I(N__78937));
    LocalMux I__19984 (
            .O(N__78963),
            .I(N__78934));
    Span4Mux_v I__19983 (
            .O(N__78960),
            .I(N__78929));
    LocalMux I__19982 (
            .O(N__78957),
            .I(N__78929));
    InMux I__19981 (
            .O(N__78956),
            .I(N__78924));
    InMux I__19980 (
            .O(N__78955),
            .I(N__78924));
    Span4Mux_h I__19979 (
            .O(N__78952),
            .I(N__78921));
    LocalMux I__19978 (
            .O(N__78949),
            .I(N__78918));
    Span4Mux_v I__19977 (
            .O(N__78944),
            .I(N__78915));
    InMux I__19976 (
            .O(N__78943),
            .I(N__78912));
    Span4Mux_h I__19975 (
            .O(N__78940),
            .I(N__78905));
    Span4Mux_v I__19974 (
            .O(N__78937),
            .I(N__78905));
    Span4Mux_v I__19973 (
            .O(N__78934),
            .I(N__78905));
    Span4Mux_h I__19972 (
            .O(N__78929),
            .I(N__78900));
    LocalMux I__19971 (
            .O(N__78924),
            .I(N__78900));
    Odrv4 I__19970 (
            .O(N__78921),
            .I(\PROM.ROMDATA.N_28_i ));
    Odrv4 I__19969 (
            .O(N__78918),
            .I(\PROM.ROMDATA.N_28_i ));
    Odrv4 I__19968 (
            .O(N__78915),
            .I(\PROM.ROMDATA.N_28_i ));
    LocalMux I__19967 (
            .O(N__78912),
            .I(\PROM.ROMDATA.N_28_i ));
    Odrv4 I__19966 (
            .O(N__78905),
            .I(\PROM.ROMDATA.N_28_i ));
    Odrv4 I__19965 (
            .O(N__78900),
            .I(\PROM.ROMDATA.N_28_i ));
    InMux I__19964 (
            .O(N__78887),
            .I(N__78884));
    LocalMux I__19963 (
            .O(N__78884),
            .I(N__78881));
    Span12Mux_s10_h I__19962 (
            .O(N__78881),
            .I(N__78878));
    Odrv12 I__19961 (
            .O(N__78878),
            .I(\PROM.ROMDATA.m183 ));
    CascadeMux I__19960 (
            .O(N__78875),
            .I(\PROM.ROMDATA.m334_ns_1_cascade_ ));
    CascadeMux I__19959 (
            .O(N__78872),
            .I(N__78869));
    InMux I__19958 (
            .O(N__78869),
            .I(N__78866));
    LocalMux I__19957 (
            .O(N__78866),
            .I(\PROM.ROMDATA.i3_mux_0 ));
    CascadeMux I__19956 (
            .O(N__78863),
            .I(N__78846));
    CascadeMux I__19955 (
            .O(N__78862),
            .I(N__78824));
    CascadeMux I__19954 (
            .O(N__78861),
            .I(N__78820));
    CascadeMux I__19953 (
            .O(N__78860),
            .I(N__78815));
    InMux I__19952 (
            .O(N__78859),
            .I(N__78799));
    InMux I__19951 (
            .O(N__78858),
            .I(N__78799));
    InMux I__19950 (
            .O(N__78857),
            .I(N__78799));
    InMux I__19949 (
            .O(N__78856),
            .I(N__78780));
    InMux I__19948 (
            .O(N__78855),
            .I(N__78780));
    InMux I__19947 (
            .O(N__78854),
            .I(N__78780));
    InMux I__19946 (
            .O(N__78853),
            .I(N__78770));
    InMux I__19945 (
            .O(N__78852),
            .I(N__78761));
    InMux I__19944 (
            .O(N__78851),
            .I(N__78761));
    InMux I__19943 (
            .O(N__78850),
            .I(N__78754));
    InMux I__19942 (
            .O(N__78849),
            .I(N__78754));
    InMux I__19941 (
            .O(N__78846),
            .I(N__78754));
    CascadeMux I__19940 (
            .O(N__78845),
            .I(N__78750));
    CascadeMux I__19939 (
            .O(N__78844),
            .I(N__78747));
    InMux I__19938 (
            .O(N__78843),
            .I(N__78741));
    InMux I__19937 (
            .O(N__78842),
            .I(N__78738));
    InMux I__19936 (
            .O(N__78841),
            .I(N__78724));
    InMux I__19935 (
            .O(N__78840),
            .I(N__78721));
    CascadeMux I__19934 (
            .O(N__78839),
            .I(N__78715));
    InMux I__19933 (
            .O(N__78838),
            .I(N__78705));
    InMux I__19932 (
            .O(N__78837),
            .I(N__78705));
    InMux I__19931 (
            .O(N__78836),
            .I(N__78705));
    CascadeMux I__19930 (
            .O(N__78835),
            .I(N__78701));
    CascadeMux I__19929 (
            .O(N__78834),
            .I(N__78697));
    CascadeMux I__19928 (
            .O(N__78833),
            .I(N__78689));
    InMux I__19927 (
            .O(N__78832),
            .I(N__78680));
    InMux I__19926 (
            .O(N__78831),
            .I(N__78680));
    InMux I__19925 (
            .O(N__78830),
            .I(N__78672));
    InMux I__19924 (
            .O(N__78829),
            .I(N__78672));
    InMux I__19923 (
            .O(N__78828),
            .I(N__78663));
    InMux I__19922 (
            .O(N__78827),
            .I(N__78663));
    InMux I__19921 (
            .O(N__78824),
            .I(N__78663));
    InMux I__19920 (
            .O(N__78823),
            .I(N__78663));
    InMux I__19919 (
            .O(N__78820),
            .I(N__78652));
    InMux I__19918 (
            .O(N__78819),
            .I(N__78652));
    InMux I__19917 (
            .O(N__78818),
            .I(N__78652));
    InMux I__19916 (
            .O(N__78815),
            .I(N__78652));
    InMux I__19915 (
            .O(N__78814),
            .I(N__78652));
    InMux I__19914 (
            .O(N__78813),
            .I(N__78641));
    InMux I__19913 (
            .O(N__78812),
            .I(N__78641));
    InMux I__19912 (
            .O(N__78811),
            .I(N__78641));
    InMux I__19911 (
            .O(N__78810),
            .I(N__78641));
    InMux I__19910 (
            .O(N__78809),
            .I(N__78641));
    InMux I__19909 (
            .O(N__78808),
            .I(N__78631));
    InMux I__19908 (
            .O(N__78807),
            .I(N__78626));
    InMux I__19907 (
            .O(N__78806),
            .I(N__78626));
    LocalMux I__19906 (
            .O(N__78799),
            .I(N__78622));
    InMux I__19905 (
            .O(N__78798),
            .I(N__78613));
    InMux I__19904 (
            .O(N__78797),
            .I(N__78613));
    InMux I__19903 (
            .O(N__78796),
            .I(N__78613));
    InMux I__19902 (
            .O(N__78795),
            .I(N__78613));
    InMux I__19901 (
            .O(N__78794),
            .I(N__78606));
    InMux I__19900 (
            .O(N__78793),
            .I(N__78606));
    InMux I__19899 (
            .O(N__78792),
            .I(N__78606));
    InMux I__19898 (
            .O(N__78791),
            .I(N__78597));
    InMux I__19897 (
            .O(N__78790),
            .I(N__78597));
    InMux I__19896 (
            .O(N__78789),
            .I(N__78597));
    InMux I__19895 (
            .O(N__78788),
            .I(N__78597));
    InMux I__19894 (
            .O(N__78787),
            .I(N__78594));
    LocalMux I__19893 (
            .O(N__78780),
            .I(N__78591));
    InMux I__19892 (
            .O(N__78779),
            .I(N__78588));
    InMux I__19891 (
            .O(N__78778),
            .I(N__78583));
    InMux I__19890 (
            .O(N__78777),
            .I(N__78583));
    InMux I__19889 (
            .O(N__78776),
            .I(N__78574));
    InMux I__19888 (
            .O(N__78775),
            .I(N__78574));
    InMux I__19887 (
            .O(N__78774),
            .I(N__78574));
    InMux I__19886 (
            .O(N__78773),
            .I(N__78574));
    LocalMux I__19885 (
            .O(N__78770),
            .I(N__78570));
    InMux I__19884 (
            .O(N__78769),
            .I(N__78560));
    InMux I__19883 (
            .O(N__78768),
            .I(N__78560));
    InMux I__19882 (
            .O(N__78767),
            .I(N__78560));
    InMux I__19881 (
            .O(N__78766),
            .I(N__78560));
    LocalMux I__19880 (
            .O(N__78761),
            .I(N__78555));
    LocalMux I__19879 (
            .O(N__78754),
            .I(N__78555));
    InMux I__19878 (
            .O(N__78753),
            .I(N__78552));
    InMux I__19877 (
            .O(N__78750),
            .I(N__78547));
    InMux I__19876 (
            .O(N__78747),
            .I(N__78547));
    InMux I__19875 (
            .O(N__78746),
            .I(N__78544));
    InMux I__19874 (
            .O(N__78745),
            .I(N__78537));
    InMux I__19873 (
            .O(N__78744),
            .I(N__78537));
    LocalMux I__19872 (
            .O(N__78741),
            .I(N__78532));
    LocalMux I__19871 (
            .O(N__78738),
            .I(N__78532));
    InMux I__19870 (
            .O(N__78737),
            .I(N__78523));
    InMux I__19869 (
            .O(N__78736),
            .I(N__78523));
    InMux I__19868 (
            .O(N__78735),
            .I(N__78523));
    InMux I__19867 (
            .O(N__78734),
            .I(N__78523));
    InMux I__19866 (
            .O(N__78733),
            .I(N__78516));
    InMux I__19865 (
            .O(N__78732),
            .I(N__78516));
    InMux I__19864 (
            .O(N__78731),
            .I(N__78516));
    InMux I__19863 (
            .O(N__78730),
            .I(N__78507));
    InMux I__19862 (
            .O(N__78729),
            .I(N__78507));
    InMux I__19861 (
            .O(N__78728),
            .I(N__78507));
    InMux I__19860 (
            .O(N__78727),
            .I(N__78507));
    LocalMux I__19859 (
            .O(N__78724),
            .I(N__78502));
    LocalMux I__19858 (
            .O(N__78721),
            .I(N__78499));
    InMux I__19857 (
            .O(N__78720),
            .I(N__78496));
    InMux I__19856 (
            .O(N__78719),
            .I(N__78489));
    InMux I__19855 (
            .O(N__78718),
            .I(N__78489));
    InMux I__19854 (
            .O(N__78715),
            .I(N__78489));
    InMux I__19853 (
            .O(N__78714),
            .I(N__78484));
    InMux I__19852 (
            .O(N__78713),
            .I(N__78484));
    InMux I__19851 (
            .O(N__78712),
            .I(N__78479));
    LocalMux I__19850 (
            .O(N__78705),
            .I(N__78476));
    CascadeMux I__19849 (
            .O(N__78704),
            .I(N__78469));
    InMux I__19848 (
            .O(N__78701),
            .I(N__78457));
    InMux I__19847 (
            .O(N__78700),
            .I(N__78457));
    InMux I__19846 (
            .O(N__78697),
            .I(N__78457));
    InMux I__19845 (
            .O(N__78696),
            .I(N__78457));
    InMux I__19844 (
            .O(N__78695),
            .I(N__78457));
    InMux I__19843 (
            .O(N__78694),
            .I(N__78454));
    InMux I__19842 (
            .O(N__78693),
            .I(N__78447));
    InMux I__19841 (
            .O(N__78692),
            .I(N__78447));
    InMux I__19840 (
            .O(N__78689),
            .I(N__78447));
    InMux I__19839 (
            .O(N__78688),
            .I(N__78442));
    InMux I__19838 (
            .O(N__78687),
            .I(N__78442));
    InMux I__19837 (
            .O(N__78686),
            .I(N__78437));
    InMux I__19836 (
            .O(N__78685),
            .I(N__78437));
    LocalMux I__19835 (
            .O(N__78680),
            .I(N__78434));
    InMux I__19834 (
            .O(N__78679),
            .I(N__78431));
    InMux I__19833 (
            .O(N__78678),
            .I(N__78426));
    InMux I__19832 (
            .O(N__78677),
            .I(N__78426));
    LocalMux I__19831 (
            .O(N__78672),
            .I(N__78417));
    LocalMux I__19830 (
            .O(N__78663),
            .I(N__78417));
    LocalMux I__19829 (
            .O(N__78652),
            .I(N__78417));
    LocalMux I__19828 (
            .O(N__78641),
            .I(N__78417));
    InMux I__19827 (
            .O(N__78640),
            .I(N__78410));
    InMux I__19826 (
            .O(N__78639),
            .I(N__78410));
    InMux I__19825 (
            .O(N__78638),
            .I(N__78410));
    InMux I__19824 (
            .O(N__78637),
            .I(N__78407));
    InMux I__19823 (
            .O(N__78636),
            .I(N__78399));
    InMux I__19822 (
            .O(N__78635),
            .I(N__78399));
    InMux I__19821 (
            .O(N__78634),
            .I(N__78396));
    LocalMux I__19820 (
            .O(N__78631),
            .I(N__78391));
    LocalMux I__19819 (
            .O(N__78626),
            .I(N__78391));
    InMux I__19818 (
            .O(N__78625),
            .I(N__78388));
    Span4Mux_h I__19817 (
            .O(N__78622),
            .I(N__78379));
    LocalMux I__19816 (
            .O(N__78613),
            .I(N__78379));
    LocalMux I__19815 (
            .O(N__78606),
            .I(N__78379));
    LocalMux I__19814 (
            .O(N__78597),
            .I(N__78379));
    LocalMux I__19813 (
            .O(N__78594),
            .I(N__78372));
    Span4Mux_v I__19812 (
            .O(N__78591),
            .I(N__78372));
    LocalMux I__19811 (
            .O(N__78588),
            .I(N__78372));
    LocalMux I__19810 (
            .O(N__78583),
            .I(N__78369));
    LocalMux I__19809 (
            .O(N__78574),
            .I(N__78366));
    CascadeMux I__19808 (
            .O(N__78573),
            .I(N__78363));
    Span4Mux_v I__19807 (
            .O(N__78570),
            .I(N__78355));
    InMux I__19806 (
            .O(N__78569),
            .I(N__78352));
    LocalMux I__19805 (
            .O(N__78560),
            .I(N__78345));
    Span4Mux_h I__19804 (
            .O(N__78555),
            .I(N__78345));
    LocalMux I__19803 (
            .O(N__78552),
            .I(N__78345));
    LocalMux I__19802 (
            .O(N__78547),
            .I(N__78340));
    LocalMux I__19801 (
            .O(N__78544),
            .I(N__78340));
    CascadeMux I__19800 (
            .O(N__78543),
            .I(N__78316));
    InMux I__19799 (
            .O(N__78542),
            .I(N__78312));
    LocalMux I__19798 (
            .O(N__78537),
            .I(N__78305));
    Span4Mux_h I__19797 (
            .O(N__78532),
            .I(N__78305));
    LocalMux I__19796 (
            .O(N__78523),
            .I(N__78305));
    LocalMux I__19795 (
            .O(N__78516),
            .I(N__78300));
    LocalMux I__19794 (
            .O(N__78507),
            .I(N__78300));
    InMux I__19793 (
            .O(N__78506),
            .I(N__78295));
    InMux I__19792 (
            .O(N__78505),
            .I(N__78295));
    Span4Mux_h I__19791 (
            .O(N__78502),
            .I(N__78290));
    Span4Mux_h I__19790 (
            .O(N__78499),
            .I(N__78290));
    LocalMux I__19789 (
            .O(N__78496),
            .I(N__78287));
    LocalMux I__19788 (
            .O(N__78489),
            .I(N__78282));
    LocalMux I__19787 (
            .O(N__78484),
            .I(N__78282));
    InMux I__19786 (
            .O(N__78483),
            .I(N__78277));
    InMux I__19785 (
            .O(N__78482),
            .I(N__78277));
    LocalMux I__19784 (
            .O(N__78479),
            .I(N__78272));
    Span4Mux_v I__19783 (
            .O(N__78476),
            .I(N__78272));
    InMux I__19782 (
            .O(N__78475),
            .I(N__78265));
    InMux I__19781 (
            .O(N__78474),
            .I(N__78265));
    InMux I__19780 (
            .O(N__78473),
            .I(N__78265));
    InMux I__19779 (
            .O(N__78472),
            .I(N__78258));
    InMux I__19778 (
            .O(N__78469),
            .I(N__78258));
    InMux I__19777 (
            .O(N__78468),
            .I(N__78258));
    LocalMux I__19776 (
            .O(N__78457),
            .I(N__78237));
    LocalMux I__19775 (
            .O(N__78454),
            .I(N__78237));
    LocalMux I__19774 (
            .O(N__78447),
            .I(N__78237));
    LocalMux I__19773 (
            .O(N__78442),
            .I(N__78237));
    LocalMux I__19772 (
            .O(N__78437),
            .I(N__78237));
    Span4Mux_h I__19771 (
            .O(N__78434),
            .I(N__78237));
    LocalMux I__19770 (
            .O(N__78431),
            .I(N__78237));
    LocalMux I__19769 (
            .O(N__78426),
            .I(N__78237));
    Span4Mux_v I__19768 (
            .O(N__78417),
            .I(N__78237));
    LocalMux I__19767 (
            .O(N__78410),
            .I(N__78237));
    LocalMux I__19766 (
            .O(N__78407),
            .I(N__78234));
    InMux I__19765 (
            .O(N__78406),
            .I(N__78227));
    InMux I__19764 (
            .O(N__78405),
            .I(N__78227));
    InMux I__19763 (
            .O(N__78404),
            .I(N__78227));
    LocalMux I__19762 (
            .O(N__78399),
            .I(N__78214));
    LocalMux I__19761 (
            .O(N__78396),
            .I(N__78214));
    Span4Mux_v I__19760 (
            .O(N__78391),
            .I(N__78214));
    LocalMux I__19759 (
            .O(N__78388),
            .I(N__78214));
    Span4Mux_v I__19758 (
            .O(N__78379),
            .I(N__78214));
    Span4Mux_h I__19757 (
            .O(N__78372),
            .I(N__78214));
    Span4Mux_h I__19756 (
            .O(N__78369),
            .I(N__78209));
    Span4Mux_v I__19755 (
            .O(N__78366),
            .I(N__78209));
    InMux I__19754 (
            .O(N__78363),
            .I(N__78206));
    InMux I__19753 (
            .O(N__78362),
            .I(N__78203));
    InMux I__19752 (
            .O(N__78361),
            .I(N__78194));
    InMux I__19751 (
            .O(N__78360),
            .I(N__78194));
    InMux I__19750 (
            .O(N__78359),
            .I(N__78194));
    InMux I__19749 (
            .O(N__78358),
            .I(N__78194));
    Span4Mux_h I__19748 (
            .O(N__78355),
            .I(N__78185));
    LocalMux I__19747 (
            .O(N__78352),
            .I(N__78185));
    Span4Mux_v I__19746 (
            .O(N__78345),
            .I(N__78185));
    Span4Mux_v I__19745 (
            .O(N__78340),
            .I(N__78185));
    InMux I__19744 (
            .O(N__78339),
            .I(N__78178));
    InMux I__19743 (
            .O(N__78338),
            .I(N__78178));
    InMux I__19742 (
            .O(N__78337),
            .I(N__78178));
    InMux I__19741 (
            .O(N__78336),
            .I(N__78169));
    InMux I__19740 (
            .O(N__78335),
            .I(N__78169));
    InMux I__19739 (
            .O(N__78334),
            .I(N__78169));
    InMux I__19738 (
            .O(N__78333),
            .I(N__78169));
    InMux I__19737 (
            .O(N__78332),
            .I(N__78160));
    InMux I__19736 (
            .O(N__78331),
            .I(N__78160));
    InMux I__19735 (
            .O(N__78330),
            .I(N__78160));
    InMux I__19734 (
            .O(N__78329),
            .I(N__78160));
    InMux I__19733 (
            .O(N__78328),
            .I(N__78151));
    InMux I__19732 (
            .O(N__78327),
            .I(N__78151));
    InMux I__19731 (
            .O(N__78326),
            .I(N__78151));
    InMux I__19730 (
            .O(N__78325),
            .I(N__78151));
    InMux I__19729 (
            .O(N__78324),
            .I(N__78142));
    InMux I__19728 (
            .O(N__78323),
            .I(N__78142));
    InMux I__19727 (
            .O(N__78322),
            .I(N__78142));
    InMux I__19726 (
            .O(N__78321),
            .I(N__78142));
    InMux I__19725 (
            .O(N__78320),
            .I(N__78133));
    InMux I__19724 (
            .O(N__78319),
            .I(N__78133));
    InMux I__19723 (
            .O(N__78316),
            .I(N__78133));
    InMux I__19722 (
            .O(N__78315),
            .I(N__78133));
    LocalMux I__19721 (
            .O(N__78312),
            .I(N__78124));
    Span4Mux_v I__19720 (
            .O(N__78305),
            .I(N__78124));
    Span4Mux_h I__19719 (
            .O(N__78300),
            .I(N__78124));
    LocalMux I__19718 (
            .O(N__78295),
            .I(N__78124));
    Span4Mux_v I__19717 (
            .O(N__78290),
            .I(N__78107));
    Span4Mux_v I__19716 (
            .O(N__78287),
            .I(N__78107));
    Span4Mux_v I__19715 (
            .O(N__78282),
            .I(N__78107));
    LocalMux I__19714 (
            .O(N__78277),
            .I(N__78107));
    Span4Mux_h I__19713 (
            .O(N__78272),
            .I(N__78107));
    LocalMux I__19712 (
            .O(N__78265),
            .I(N__78107));
    LocalMux I__19711 (
            .O(N__78258),
            .I(N__78107));
    Span4Mux_v I__19710 (
            .O(N__78237),
            .I(N__78107));
    Span4Mux_h I__19709 (
            .O(N__78234),
            .I(N__78100));
    LocalMux I__19708 (
            .O(N__78227),
            .I(N__78100));
    Span4Mux_h I__19707 (
            .O(N__78214),
            .I(N__78100));
    Odrv4 I__19706 (
            .O(N__78209),
            .I(progRomAddress_1));
    LocalMux I__19705 (
            .O(N__78206),
            .I(progRomAddress_1));
    LocalMux I__19704 (
            .O(N__78203),
            .I(progRomAddress_1));
    LocalMux I__19703 (
            .O(N__78194),
            .I(progRomAddress_1));
    Odrv4 I__19702 (
            .O(N__78185),
            .I(progRomAddress_1));
    LocalMux I__19701 (
            .O(N__78178),
            .I(progRomAddress_1));
    LocalMux I__19700 (
            .O(N__78169),
            .I(progRomAddress_1));
    LocalMux I__19699 (
            .O(N__78160),
            .I(progRomAddress_1));
    LocalMux I__19698 (
            .O(N__78151),
            .I(progRomAddress_1));
    LocalMux I__19697 (
            .O(N__78142),
            .I(progRomAddress_1));
    LocalMux I__19696 (
            .O(N__78133),
            .I(progRomAddress_1));
    Odrv4 I__19695 (
            .O(N__78124),
            .I(progRomAddress_1));
    Odrv4 I__19694 (
            .O(N__78107),
            .I(progRomAddress_1));
    Odrv4 I__19693 (
            .O(N__78100),
            .I(progRomAddress_1));
    CascadeMux I__19692 (
            .O(N__78071),
            .I(N__78056));
    CascadeMux I__19691 (
            .O(N__78070),
            .I(N__78051));
    InMux I__19690 (
            .O(N__78069),
            .I(N__78044));
    InMux I__19689 (
            .O(N__78068),
            .I(N__78044));
    InMux I__19688 (
            .O(N__78067),
            .I(N__78032));
    InMux I__19687 (
            .O(N__78066),
            .I(N__78029));
    InMux I__19686 (
            .O(N__78065),
            .I(N__78017));
    InMux I__19685 (
            .O(N__78064),
            .I(N__78012));
    InMux I__19684 (
            .O(N__78063),
            .I(N__78012));
    InMux I__19683 (
            .O(N__78062),
            .I(N__78006));
    InMux I__19682 (
            .O(N__78061),
            .I(N__78006));
    InMux I__19681 (
            .O(N__78060),
            .I(N__78003));
    InMux I__19680 (
            .O(N__78059),
            .I(N__77996));
    InMux I__19679 (
            .O(N__78056),
            .I(N__77996));
    InMux I__19678 (
            .O(N__78055),
            .I(N__77996));
    CascadeMux I__19677 (
            .O(N__78054),
            .I(N__77990));
    InMux I__19676 (
            .O(N__78051),
            .I(N__77983));
    InMux I__19675 (
            .O(N__78050),
            .I(N__77983));
    CascadeMux I__19674 (
            .O(N__78049),
            .I(N__77978));
    LocalMux I__19673 (
            .O(N__78044),
            .I(N__77970));
    CascadeMux I__19672 (
            .O(N__78043),
            .I(N__77967));
    CascadeMux I__19671 (
            .O(N__78042),
            .I(N__77962));
    InMux I__19670 (
            .O(N__78041),
            .I(N__77958));
    CascadeMux I__19669 (
            .O(N__78040),
            .I(N__77950));
    CascadeMux I__19668 (
            .O(N__78039),
            .I(N__77947));
    CascadeMux I__19667 (
            .O(N__78038),
            .I(N__77944));
    CascadeMux I__19666 (
            .O(N__78037),
            .I(N__77941));
    CascadeMux I__19665 (
            .O(N__78036),
            .I(N__77937));
    CascadeMux I__19664 (
            .O(N__78035),
            .I(N__77934));
    LocalMux I__19663 (
            .O(N__78032),
            .I(N__77929));
    LocalMux I__19662 (
            .O(N__78029),
            .I(N__77926));
    InMux I__19661 (
            .O(N__78028),
            .I(N__77921));
    InMux I__19660 (
            .O(N__78027),
            .I(N__77921));
    InMux I__19659 (
            .O(N__78026),
            .I(N__77912));
    InMux I__19658 (
            .O(N__78025),
            .I(N__77912));
    InMux I__19657 (
            .O(N__78024),
            .I(N__77912));
    InMux I__19656 (
            .O(N__78023),
            .I(N__77912));
    CascadeMux I__19655 (
            .O(N__78022),
            .I(N__77903));
    CascadeMux I__19654 (
            .O(N__78021),
            .I(N__77900));
    CascadeMux I__19653 (
            .O(N__78020),
            .I(N__77889));
    LocalMux I__19652 (
            .O(N__78017),
            .I(N__77870));
    LocalMux I__19651 (
            .O(N__78012),
            .I(N__77867));
    InMux I__19650 (
            .O(N__78011),
            .I(N__77859));
    LocalMux I__19649 (
            .O(N__78006),
            .I(N__77856));
    LocalMux I__19648 (
            .O(N__78003),
            .I(N__77853));
    LocalMux I__19647 (
            .O(N__77996),
            .I(N__77850));
    InMux I__19646 (
            .O(N__77995),
            .I(N__77847));
    CascadeMux I__19645 (
            .O(N__77994),
            .I(N__77844));
    InMux I__19644 (
            .O(N__77993),
            .I(N__77829));
    InMux I__19643 (
            .O(N__77990),
            .I(N__77829));
    InMux I__19642 (
            .O(N__77989),
            .I(N__77829));
    InMux I__19641 (
            .O(N__77988),
            .I(N__77829));
    LocalMux I__19640 (
            .O(N__77983),
            .I(N__77826));
    InMux I__19639 (
            .O(N__77982),
            .I(N__77817));
    InMux I__19638 (
            .O(N__77981),
            .I(N__77817));
    InMux I__19637 (
            .O(N__77978),
            .I(N__77817));
    InMux I__19636 (
            .O(N__77977),
            .I(N__77817));
    CascadeMux I__19635 (
            .O(N__77976),
            .I(N__77813));
    CascadeMux I__19634 (
            .O(N__77975),
            .I(N__77809));
    CascadeMux I__19633 (
            .O(N__77974),
            .I(N__77800));
    CascadeMux I__19632 (
            .O(N__77973),
            .I(N__77797));
    Span4Mux_h I__19631 (
            .O(N__77970),
            .I(N__77790));
    InMux I__19630 (
            .O(N__77967),
            .I(N__77785));
    InMux I__19629 (
            .O(N__77966),
            .I(N__77785));
    InMux I__19628 (
            .O(N__77965),
            .I(N__77778));
    InMux I__19627 (
            .O(N__77962),
            .I(N__77778));
    InMux I__19626 (
            .O(N__77961),
            .I(N__77778));
    LocalMux I__19625 (
            .O(N__77958),
            .I(N__77775));
    InMux I__19624 (
            .O(N__77957),
            .I(N__77766));
    InMux I__19623 (
            .O(N__77956),
            .I(N__77766));
    InMux I__19622 (
            .O(N__77955),
            .I(N__77766));
    InMux I__19621 (
            .O(N__77954),
            .I(N__77766));
    InMux I__19620 (
            .O(N__77953),
            .I(N__77755));
    InMux I__19619 (
            .O(N__77950),
            .I(N__77755));
    InMux I__19618 (
            .O(N__77947),
            .I(N__77755));
    InMux I__19617 (
            .O(N__77944),
            .I(N__77755));
    InMux I__19616 (
            .O(N__77941),
            .I(N__77755));
    InMux I__19615 (
            .O(N__77940),
            .I(N__77752));
    InMux I__19614 (
            .O(N__77937),
            .I(N__77745));
    InMux I__19613 (
            .O(N__77934),
            .I(N__77745));
    InMux I__19612 (
            .O(N__77933),
            .I(N__77745));
    InMux I__19611 (
            .O(N__77932),
            .I(N__77740));
    Span4Mux_h I__19610 (
            .O(N__77929),
            .I(N__77733));
    Span4Mux_v I__19609 (
            .O(N__77926),
            .I(N__77733));
    LocalMux I__19608 (
            .O(N__77921),
            .I(N__77733));
    LocalMux I__19607 (
            .O(N__77912),
            .I(N__77730));
    InMux I__19606 (
            .O(N__77911),
            .I(N__77723));
    InMux I__19605 (
            .O(N__77910),
            .I(N__77723));
    InMux I__19604 (
            .O(N__77909),
            .I(N__77723));
    InMux I__19603 (
            .O(N__77908),
            .I(N__77720));
    InMux I__19602 (
            .O(N__77907),
            .I(N__77715));
    InMux I__19601 (
            .O(N__77906),
            .I(N__77715));
    InMux I__19600 (
            .O(N__77903),
            .I(N__77708));
    InMux I__19599 (
            .O(N__77900),
            .I(N__77708));
    InMux I__19598 (
            .O(N__77899),
            .I(N__77708));
    InMux I__19597 (
            .O(N__77898),
            .I(N__77701));
    InMux I__19596 (
            .O(N__77897),
            .I(N__77701));
    InMux I__19595 (
            .O(N__77896),
            .I(N__77701));
    CascadeMux I__19594 (
            .O(N__77895),
            .I(N__77697));
    CascadeMux I__19593 (
            .O(N__77894),
            .I(N__77694));
    CascadeMux I__19592 (
            .O(N__77893),
            .I(N__77685));
    InMux I__19591 (
            .O(N__77892),
            .I(N__77682));
    InMux I__19590 (
            .O(N__77889),
            .I(N__77675));
    InMux I__19589 (
            .O(N__77888),
            .I(N__77675));
    InMux I__19588 (
            .O(N__77887),
            .I(N__77675));
    InMux I__19587 (
            .O(N__77886),
            .I(N__77668));
    InMux I__19586 (
            .O(N__77885),
            .I(N__77668));
    InMux I__19585 (
            .O(N__77884),
            .I(N__77668));
    InMux I__19584 (
            .O(N__77883),
            .I(N__77659));
    InMux I__19583 (
            .O(N__77882),
            .I(N__77659));
    InMux I__19582 (
            .O(N__77881),
            .I(N__77659));
    InMux I__19581 (
            .O(N__77880),
            .I(N__77659));
    InMux I__19580 (
            .O(N__77879),
            .I(N__77654));
    InMux I__19579 (
            .O(N__77878),
            .I(N__77654));
    InMux I__19578 (
            .O(N__77877),
            .I(N__77647));
    InMux I__19577 (
            .O(N__77876),
            .I(N__77647));
    InMux I__19576 (
            .O(N__77875),
            .I(N__77647));
    InMux I__19575 (
            .O(N__77874),
            .I(N__77642));
    InMux I__19574 (
            .O(N__77873),
            .I(N__77642));
    Span4Mux_v I__19573 (
            .O(N__77870),
            .I(N__77639));
    Span4Mux_v I__19572 (
            .O(N__77867),
            .I(N__77636));
    InMux I__19571 (
            .O(N__77866),
            .I(N__77627));
    InMux I__19570 (
            .O(N__77865),
            .I(N__77627));
    InMux I__19569 (
            .O(N__77864),
            .I(N__77627));
    InMux I__19568 (
            .O(N__77863),
            .I(N__77627));
    InMux I__19567 (
            .O(N__77862),
            .I(N__77624));
    LocalMux I__19566 (
            .O(N__77859),
            .I(N__77621));
    Span4Mux_h I__19565 (
            .O(N__77856),
            .I(N__77605));
    Span4Mux_h I__19564 (
            .O(N__77853),
            .I(N__77598));
    Span4Mux_v I__19563 (
            .O(N__77850),
            .I(N__77598));
    LocalMux I__19562 (
            .O(N__77847),
            .I(N__77598));
    InMux I__19561 (
            .O(N__77844),
            .I(N__77591));
    InMux I__19560 (
            .O(N__77843),
            .I(N__77591));
    InMux I__19559 (
            .O(N__77842),
            .I(N__77591));
    CascadeMux I__19558 (
            .O(N__77841),
            .I(N__77587));
    CascadeMux I__19557 (
            .O(N__77840),
            .I(N__77584));
    CascadeMux I__19556 (
            .O(N__77839),
            .I(N__77580));
    CascadeMux I__19555 (
            .O(N__77838),
            .I(N__77577));
    LocalMux I__19554 (
            .O(N__77829),
            .I(N__77568));
    Span4Mux_h I__19553 (
            .O(N__77826),
            .I(N__77568));
    LocalMux I__19552 (
            .O(N__77817),
            .I(N__77568));
    InMux I__19551 (
            .O(N__77816),
            .I(N__77559));
    InMux I__19550 (
            .O(N__77813),
            .I(N__77559));
    InMux I__19549 (
            .O(N__77812),
            .I(N__77559));
    InMux I__19548 (
            .O(N__77809),
            .I(N__77559));
    InMux I__19547 (
            .O(N__77808),
            .I(N__77548));
    InMux I__19546 (
            .O(N__77807),
            .I(N__77548));
    InMux I__19545 (
            .O(N__77806),
            .I(N__77548));
    InMux I__19544 (
            .O(N__77805),
            .I(N__77548));
    InMux I__19543 (
            .O(N__77804),
            .I(N__77548));
    InMux I__19542 (
            .O(N__77803),
            .I(N__77539));
    InMux I__19541 (
            .O(N__77800),
            .I(N__77539));
    InMux I__19540 (
            .O(N__77797),
            .I(N__77539));
    InMux I__19539 (
            .O(N__77796),
            .I(N__77539));
    InMux I__19538 (
            .O(N__77795),
            .I(N__77532));
    InMux I__19537 (
            .O(N__77794),
            .I(N__77532));
    InMux I__19536 (
            .O(N__77793),
            .I(N__77532));
    Span4Mux_v I__19535 (
            .O(N__77790),
            .I(N__77525));
    LocalMux I__19534 (
            .O(N__77785),
            .I(N__77525));
    LocalMux I__19533 (
            .O(N__77778),
            .I(N__77525));
    Span4Mux_h I__19532 (
            .O(N__77775),
            .I(N__77518));
    LocalMux I__19531 (
            .O(N__77766),
            .I(N__77518));
    LocalMux I__19530 (
            .O(N__77755),
            .I(N__77518));
    LocalMux I__19529 (
            .O(N__77752),
            .I(N__77515));
    LocalMux I__19528 (
            .O(N__77745),
            .I(N__77512));
    InMux I__19527 (
            .O(N__77744),
            .I(N__77507));
    InMux I__19526 (
            .O(N__77743),
            .I(N__77507));
    LocalMux I__19525 (
            .O(N__77740),
            .I(N__77498));
    Span4Mux_h I__19524 (
            .O(N__77733),
            .I(N__77498));
    Span4Mux_h I__19523 (
            .O(N__77730),
            .I(N__77498));
    LocalMux I__19522 (
            .O(N__77723),
            .I(N__77498));
    LocalMux I__19521 (
            .O(N__77720),
            .I(N__77489));
    LocalMux I__19520 (
            .O(N__77715),
            .I(N__77489));
    LocalMux I__19519 (
            .O(N__77708),
            .I(N__77489));
    LocalMux I__19518 (
            .O(N__77701),
            .I(N__77489));
    InMux I__19517 (
            .O(N__77700),
            .I(N__77480));
    InMux I__19516 (
            .O(N__77697),
            .I(N__77480));
    InMux I__19515 (
            .O(N__77694),
            .I(N__77480));
    InMux I__19514 (
            .O(N__77693),
            .I(N__77480));
    InMux I__19513 (
            .O(N__77692),
            .I(N__77473));
    InMux I__19512 (
            .O(N__77691),
            .I(N__77473));
    InMux I__19511 (
            .O(N__77690),
            .I(N__77473));
    InMux I__19510 (
            .O(N__77689),
            .I(N__77466));
    InMux I__19509 (
            .O(N__77688),
            .I(N__77466));
    InMux I__19508 (
            .O(N__77685),
            .I(N__77466));
    LocalMux I__19507 (
            .O(N__77682),
            .I(N__77459));
    LocalMux I__19506 (
            .O(N__77675),
            .I(N__77459));
    LocalMux I__19505 (
            .O(N__77668),
            .I(N__77459));
    LocalMux I__19504 (
            .O(N__77659),
            .I(N__77450));
    LocalMux I__19503 (
            .O(N__77654),
            .I(N__77450));
    LocalMux I__19502 (
            .O(N__77647),
            .I(N__77450));
    LocalMux I__19501 (
            .O(N__77642),
            .I(N__77450));
    Span4Mux_h I__19500 (
            .O(N__77639),
            .I(N__77441));
    Span4Mux_v I__19499 (
            .O(N__77636),
            .I(N__77441));
    LocalMux I__19498 (
            .O(N__77627),
            .I(N__77441));
    LocalMux I__19497 (
            .O(N__77624),
            .I(N__77441));
    Span12Mux_s11_h I__19496 (
            .O(N__77621),
            .I(N__77438));
    InMux I__19495 (
            .O(N__77620),
            .I(N__77427));
    InMux I__19494 (
            .O(N__77619),
            .I(N__77427));
    InMux I__19493 (
            .O(N__77618),
            .I(N__77427));
    InMux I__19492 (
            .O(N__77617),
            .I(N__77427));
    InMux I__19491 (
            .O(N__77616),
            .I(N__77427));
    InMux I__19490 (
            .O(N__77615),
            .I(N__77420));
    InMux I__19489 (
            .O(N__77614),
            .I(N__77420));
    InMux I__19488 (
            .O(N__77613),
            .I(N__77420));
    InMux I__19487 (
            .O(N__77612),
            .I(N__77415));
    InMux I__19486 (
            .O(N__77611),
            .I(N__77415));
    InMux I__19485 (
            .O(N__77610),
            .I(N__77408));
    InMux I__19484 (
            .O(N__77609),
            .I(N__77408));
    InMux I__19483 (
            .O(N__77608),
            .I(N__77408));
    Span4Mux_h I__19482 (
            .O(N__77605),
            .I(N__77401));
    Span4Mux_h I__19481 (
            .O(N__77598),
            .I(N__77401));
    LocalMux I__19480 (
            .O(N__77591),
            .I(N__77401));
    InMux I__19479 (
            .O(N__77590),
            .I(N__77392));
    InMux I__19478 (
            .O(N__77587),
            .I(N__77392));
    InMux I__19477 (
            .O(N__77584),
            .I(N__77392));
    InMux I__19476 (
            .O(N__77583),
            .I(N__77392));
    InMux I__19475 (
            .O(N__77580),
            .I(N__77383));
    InMux I__19474 (
            .O(N__77577),
            .I(N__77383));
    InMux I__19473 (
            .O(N__77576),
            .I(N__77383));
    InMux I__19472 (
            .O(N__77575),
            .I(N__77383));
    Span4Mux_v I__19471 (
            .O(N__77568),
            .I(N__77378));
    LocalMux I__19470 (
            .O(N__77559),
            .I(N__77378));
    LocalMux I__19469 (
            .O(N__77548),
            .I(N__77373));
    LocalMux I__19468 (
            .O(N__77539),
            .I(N__77373));
    LocalMux I__19467 (
            .O(N__77532),
            .I(N__77366));
    Span4Mux_h I__19466 (
            .O(N__77525),
            .I(N__77366));
    Span4Mux_v I__19465 (
            .O(N__77518),
            .I(N__77366));
    Span4Mux_v I__19464 (
            .O(N__77515),
            .I(N__77343));
    Span4Mux_h I__19463 (
            .O(N__77512),
            .I(N__77343));
    LocalMux I__19462 (
            .O(N__77507),
            .I(N__77343));
    Span4Mux_v I__19461 (
            .O(N__77498),
            .I(N__77343));
    Span4Mux_v I__19460 (
            .O(N__77489),
            .I(N__77343));
    LocalMux I__19459 (
            .O(N__77480),
            .I(N__77343));
    LocalMux I__19458 (
            .O(N__77473),
            .I(N__77343));
    LocalMux I__19457 (
            .O(N__77466),
            .I(N__77343));
    Span4Mux_v I__19456 (
            .O(N__77459),
            .I(N__77343));
    Span4Mux_v I__19455 (
            .O(N__77450),
            .I(N__77343));
    Span4Mux_h I__19454 (
            .O(N__77441),
            .I(N__77343));
    Odrv12 I__19453 (
            .O(N__77438),
            .I(progRomAddress_2));
    LocalMux I__19452 (
            .O(N__77427),
            .I(progRomAddress_2));
    LocalMux I__19451 (
            .O(N__77420),
            .I(progRomAddress_2));
    LocalMux I__19450 (
            .O(N__77415),
            .I(progRomAddress_2));
    LocalMux I__19449 (
            .O(N__77408),
            .I(progRomAddress_2));
    Odrv4 I__19448 (
            .O(N__77401),
            .I(progRomAddress_2));
    LocalMux I__19447 (
            .O(N__77392),
            .I(progRomAddress_2));
    LocalMux I__19446 (
            .O(N__77383),
            .I(progRomAddress_2));
    Odrv4 I__19445 (
            .O(N__77378),
            .I(progRomAddress_2));
    Odrv4 I__19444 (
            .O(N__77373),
            .I(progRomAddress_2));
    Odrv4 I__19443 (
            .O(N__77366),
            .I(progRomAddress_2));
    Odrv4 I__19442 (
            .O(N__77343),
            .I(progRomAddress_2));
    InMux I__19441 (
            .O(N__77318),
            .I(N__77305));
    InMux I__19440 (
            .O(N__77317),
            .I(N__77298));
    InMux I__19439 (
            .O(N__77316),
            .I(N__77287));
    InMux I__19438 (
            .O(N__77315),
            .I(N__77287));
    CascadeMux I__19437 (
            .O(N__77314),
            .I(N__77284));
    InMux I__19436 (
            .O(N__77313),
            .I(N__77275));
    InMux I__19435 (
            .O(N__77312),
            .I(N__77275));
    InMux I__19434 (
            .O(N__77311),
            .I(N__77268));
    InMux I__19433 (
            .O(N__77310),
            .I(N__77265));
    InMux I__19432 (
            .O(N__77309),
            .I(N__77262));
    InMux I__19431 (
            .O(N__77308),
            .I(N__77259));
    LocalMux I__19430 (
            .O(N__77305),
            .I(N__77231));
    InMux I__19429 (
            .O(N__77304),
            .I(N__77222));
    InMux I__19428 (
            .O(N__77303),
            .I(N__77222));
    InMux I__19427 (
            .O(N__77302),
            .I(N__77222));
    InMux I__19426 (
            .O(N__77301),
            .I(N__77222));
    LocalMux I__19425 (
            .O(N__77298),
            .I(N__77219));
    InMux I__19424 (
            .O(N__77297),
            .I(N__77214));
    InMux I__19423 (
            .O(N__77296),
            .I(N__77214));
    InMux I__19422 (
            .O(N__77295),
            .I(N__77205));
    InMux I__19421 (
            .O(N__77294),
            .I(N__77205));
    InMux I__19420 (
            .O(N__77293),
            .I(N__77205));
    InMux I__19419 (
            .O(N__77292),
            .I(N__77205));
    LocalMux I__19418 (
            .O(N__77287),
            .I(N__77202));
    InMux I__19417 (
            .O(N__77284),
            .I(N__77193));
    InMux I__19416 (
            .O(N__77283),
            .I(N__77176));
    InMux I__19415 (
            .O(N__77282),
            .I(N__77176));
    InMux I__19414 (
            .O(N__77281),
            .I(N__77166));
    InMux I__19413 (
            .O(N__77280),
            .I(N__77166));
    LocalMux I__19412 (
            .O(N__77275),
            .I(N__77161));
    InMux I__19411 (
            .O(N__77274),
            .I(N__77152));
    InMux I__19410 (
            .O(N__77273),
            .I(N__77152));
    InMux I__19409 (
            .O(N__77272),
            .I(N__77152));
    InMux I__19408 (
            .O(N__77271),
            .I(N__77152));
    LocalMux I__19407 (
            .O(N__77268),
            .I(N__77137));
    LocalMux I__19406 (
            .O(N__77265),
            .I(N__77132));
    LocalMux I__19405 (
            .O(N__77262),
            .I(N__77132));
    LocalMux I__19404 (
            .O(N__77259),
            .I(N__77129));
    InMux I__19403 (
            .O(N__77258),
            .I(N__77126));
    InMux I__19402 (
            .O(N__77257),
            .I(N__77109));
    InMux I__19401 (
            .O(N__77256),
            .I(N__77109));
    InMux I__19400 (
            .O(N__77255),
            .I(N__77100));
    InMux I__19399 (
            .O(N__77254),
            .I(N__77100));
    InMux I__19398 (
            .O(N__77253),
            .I(N__77100));
    InMux I__19397 (
            .O(N__77252),
            .I(N__77100));
    InMux I__19396 (
            .O(N__77251),
            .I(N__77093));
    InMux I__19395 (
            .O(N__77250),
            .I(N__77093));
    InMux I__19394 (
            .O(N__77249),
            .I(N__77093));
    InMux I__19393 (
            .O(N__77248),
            .I(N__77088));
    InMux I__19392 (
            .O(N__77247),
            .I(N__77088));
    InMux I__19391 (
            .O(N__77246),
            .I(N__77081));
    InMux I__19390 (
            .O(N__77245),
            .I(N__77081));
    InMux I__19389 (
            .O(N__77244),
            .I(N__77081));
    InMux I__19388 (
            .O(N__77243),
            .I(N__77074));
    InMux I__19387 (
            .O(N__77242),
            .I(N__77074));
    InMux I__19386 (
            .O(N__77241),
            .I(N__77074));
    InMux I__19385 (
            .O(N__77240),
            .I(N__77062));
    InMux I__19384 (
            .O(N__77239),
            .I(N__77055));
    InMux I__19383 (
            .O(N__77238),
            .I(N__77055));
    InMux I__19382 (
            .O(N__77237),
            .I(N__77055));
    InMux I__19381 (
            .O(N__77236),
            .I(N__77048));
    InMux I__19380 (
            .O(N__77235),
            .I(N__77048));
    InMux I__19379 (
            .O(N__77234),
            .I(N__77048));
    Span4Mux_h I__19378 (
            .O(N__77231),
            .I(N__77039));
    LocalMux I__19377 (
            .O(N__77222),
            .I(N__77039));
    Span4Mux_v I__19376 (
            .O(N__77219),
            .I(N__77039));
    LocalMux I__19375 (
            .O(N__77214),
            .I(N__77039));
    LocalMux I__19374 (
            .O(N__77205),
            .I(N__77034));
    Span4Mux_v I__19373 (
            .O(N__77202),
            .I(N__77034));
    InMux I__19372 (
            .O(N__77201),
            .I(N__77027));
    InMux I__19371 (
            .O(N__77200),
            .I(N__77027));
    InMux I__19370 (
            .O(N__77199),
            .I(N__77027));
    InMux I__19369 (
            .O(N__77198),
            .I(N__77020));
    InMux I__19368 (
            .O(N__77197),
            .I(N__77020));
    InMux I__19367 (
            .O(N__77196),
            .I(N__77020));
    LocalMux I__19366 (
            .O(N__77193),
            .I(N__77017));
    InMux I__19365 (
            .O(N__77192),
            .I(N__77010));
    InMux I__19364 (
            .O(N__77191),
            .I(N__77010));
    InMux I__19363 (
            .O(N__77190),
            .I(N__77010));
    InMux I__19362 (
            .O(N__77189),
            .I(N__77003));
    InMux I__19361 (
            .O(N__77188),
            .I(N__77003));
    InMux I__19360 (
            .O(N__77187),
            .I(N__77003));
    InMux I__19359 (
            .O(N__77186),
            .I(N__76998));
    InMux I__19358 (
            .O(N__77185),
            .I(N__76998));
    InMux I__19357 (
            .O(N__77184),
            .I(N__76995));
    InMux I__19356 (
            .O(N__77183),
            .I(N__76988));
    InMux I__19355 (
            .O(N__77182),
            .I(N__76988));
    InMux I__19354 (
            .O(N__77181),
            .I(N__76988));
    LocalMux I__19353 (
            .O(N__77176),
            .I(N__76985));
    InMux I__19352 (
            .O(N__77175),
            .I(N__76982));
    InMux I__19351 (
            .O(N__77174),
            .I(N__76979));
    InMux I__19350 (
            .O(N__77173),
            .I(N__76970));
    InMux I__19349 (
            .O(N__77172),
            .I(N__76970));
    InMux I__19348 (
            .O(N__77171),
            .I(N__76970));
    LocalMux I__19347 (
            .O(N__77166),
            .I(N__76967));
    InMux I__19346 (
            .O(N__77165),
            .I(N__76960));
    InMux I__19345 (
            .O(N__77164),
            .I(N__76960));
    Span4Mux_v I__19344 (
            .O(N__77161),
            .I(N__76957));
    LocalMux I__19343 (
            .O(N__77152),
            .I(N__76954));
    InMux I__19342 (
            .O(N__77151),
            .I(N__76947));
    InMux I__19341 (
            .O(N__77150),
            .I(N__76947));
    InMux I__19340 (
            .O(N__77149),
            .I(N__76947));
    InMux I__19339 (
            .O(N__77148),
            .I(N__76938));
    InMux I__19338 (
            .O(N__77147),
            .I(N__76938));
    InMux I__19337 (
            .O(N__77146),
            .I(N__76938));
    InMux I__19336 (
            .O(N__77145),
            .I(N__76938));
    InMux I__19335 (
            .O(N__77144),
            .I(N__76914));
    InMux I__19334 (
            .O(N__77143),
            .I(N__76914));
    InMux I__19333 (
            .O(N__77142),
            .I(N__76914));
    InMux I__19332 (
            .O(N__77141),
            .I(N__76914));
    InMux I__19331 (
            .O(N__77140),
            .I(N__76914));
    Span4Mux_h I__19330 (
            .O(N__77137),
            .I(N__76904));
    Span4Mux_v I__19329 (
            .O(N__77132),
            .I(N__76904));
    Span4Mux_h I__19328 (
            .O(N__77129),
            .I(N__76899));
    LocalMux I__19327 (
            .O(N__77126),
            .I(N__76899));
    InMux I__19326 (
            .O(N__77125),
            .I(N__76890));
    InMux I__19325 (
            .O(N__77124),
            .I(N__76890));
    InMux I__19324 (
            .O(N__77123),
            .I(N__76890));
    InMux I__19323 (
            .O(N__77122),
            .I(N__76890));
    InMux I__19322 (
            .O(N__77121),
            .I(N__76879));
    InMux I__19321 (
            .O(N__77120),
            .I(N__76879));
    InMux I__19320 (
            .O(N__77119),
            .I(N__76879));
    InMux I__19319 (
            .O(N__77118),
            .I(N__76879));
    InMux I__19318 (
            .O(N__77117),
            .I(N__76879));
    InMux I__19317 (
            .O(N__77116),
            .I(N__76872));
    InMux I__19316 (
            .O(N__77115),
            .I(N__76872));
    InMux I__19315 (
            .O(N__77114),
            .I(N__76872));
    LocalMux I__19314 (
            .O(N__77109),
            .I(N__76865));
    LocalMux I__19313 (
            .O(N__77100),
            .I(N__76865));
    LocalMux I__19312 (
            .O(N__77093),
            .I(N__76865));
    LocalMux I__19311 (
            .O(N__77088),
            .I(N__76858));
    LocalMux I__19310 (
            .O(N__77081),
            .I(N__76858));
    LocalMux I__19309 (
            .O(N__77074),
            .I(N__76858));
    InMux I__19308 (
            .O(N__77073),
            .I(N__76851));
    InMux I__19307 (
            .O(N__77072),
            .I(N__76851));
    InMux I__19306 (
            .O(N__77071),
            .I(N__76851));
    InMux I__19305 (
            .O(N__77070),
            .I(N__76838));
    InMux I__19304 (
            .O(N__77069),
            .I(N__76838));
    InMux I__19303 (
            .O(N__77068),
            .I(N__76838));
    InMux I__19302 (
            .O(N__77067),
            .I(N__76838));
    InMux I__19301 (
            .O(N__77066),
            .I(N__76838));
    InMux I__19300 (
            .O(N__77065),
            .I(N__76838));
    LocalMux I__19299 (
            .O(N__77062),
            .I(N__76831));
    LocalMux I__19298 (
            .O(N__77055),
            .I(N__76831));
    LocalMux I__19297 (
            .O(N__77048),
            .I(N__76831));
    Span4Mux_h I__19296 (
            .O(N__77039),
            .I(N__76822));
    Span4Mux_h I__19295 (
            .O(N__77034),
            .I(N__76822));
    LocalMux I__19294 (
            .O(N__77027),
            .I(N__76822));
    LocalMux I__19293 (
            .O(N__77020),
            .I(N__76822));
    Span4Mux_v I__19292 (
            .O(N__77017),
            .I(N__76811));
    LocalMux I__19291 (
            .O(N__77010),
            .I(N__76811));
    LocalMux I__19290 (
            .O(N__77003),
            .I(N__76811));
    LocalMux I__19289 (
            .O(N__76998),
            .I(N__76811));
    LocalMux I__19288 (
            .O(N__76995),
            .I(N__76811));
    LocalMux I__19287 (
            .O(N__76988),
            .I(N__76802));
    Span4Mux_v I__19286 (
            .O(N__76985),
            .I(N__76802));
    LocalMux I__19285 (
            .O(N__76982),
            .I(N__76802));
    LocalMux I__19284 (
            .O(N__76979),
            .I(N__76802));
    InMux I__19283 (
            .O(N__76978),
            .I(N__76797));
    InMux I__19282 (
            .O(N__76977),
            .I(N__76797));
    LocalMux I__19281 (
            .O(N__76970),
            .I(N__76792));
    Span12Mux_s10_v I__19280 (
            .O(N__76967),
            .I(N__76792));
    InMux I__19279 (
            .O(N__76966),
            .I(N__76787));
    InMux I__19278 (
            .O(N__76965),
            .I(N__76787));
    LocalMux I__19277 (
            .O(N__76960),
            .I(N__76784));
    Span4Mux_h I__19276 (
            .O(N__76957),
            .I(N__76775));
    Span4Mux_v I__19275 (
            .O(N__76954),
            .I(N__76775));
    LocalMux I__19274 (
            .O(N__76947),
            .I(N__76775));
    LocalMux I__19273 (
            .O(N__76938),
            .I(N__76775));
    InMux I__19272 (
            .O(N__76937),
            .I(N__76762));
    InMux I__19271 (
            .O(N__76936),
            .I(N__76762));
    InMux I__19270 (
            .O(N__76935),
            .I(N__76762));
    InMux I__19269 (
            .O(N__76934),
            .I(N__76762));
    InMux I__19268 (
            .O(N__76933),
            .I(N__76762));
    InMux I__19267 (
            .O(N__76932),
            .I(N__76762));
    InMux I__19266 (
            .O(N__76931),
            .I(N__76753));
    InMux I__19265 (
            .O(N__76930),
            .I(N__76753));
    InMux I__19264 (
            .O(N__76929),
            .I(N__76753));
    InMux I__19263 (
            .O(N__76928),
            .I(N__76753));
    InMux I__19262 (
            .O(N__76927),
            .I(N__76746));
    InMux I__19261 (
            .O(N__76926),
            .I(N__76746));
    InMux I__19260 (
            .O(N__76925),
            .I(N__76746));
    LocalMux I__19259 (
            .O(N__76914),
            .I(N__76743));
    InMux I__19258 (
            .O(N__76913),
            .I(N__76732));
    InMux I__19257 (
            .O(N__76912),
            .I(N__76732));
    InMux I__19256 (
            .O(N__76911),
            .I(N__76732));
    InMux I__19255 (
            .O(N__76910),
            .I(N__76732));
    InMux I__19254 (
            .O(N__76909),
            .I(N__76732));
    Span4Mux_h I__19253 (
            .O(N__76904),
            .I(N__76723));
    Span4Mux_h I__19252 (
            .O(N__76899),
            .I(N__76723));
    LocalMux I__19251 (
            .O(N__76890),
            .I(N__76723));
    LocalMux I__19250 (
            .O(N__76879),
            .I(N__76723));
    LocalMux I__19249 (
            .O(N__76872),
            .I(N__76704));
    Span4Mux_v I__19248 (
            .O(N__76865),
            .I(N__76704));
    Span4Mux_v I__19247 (
            .O(N__76858),
            .I(N__76704));
    LocalMux I__19246 (
            .O(N__76851),
            .I(N__76704));
    LocalMux I__19245 (
            .O(N__76838),
            .I(N__76704));
    Span4Mux_v I__19244 (
            .O(N__76831),
            .I(N__76704));
    Span4Mux_v I__19243 (
            .O(N__76822),
            .I(N__76704));
    Span4Mux_v I__19242 (
            .O(N__76811),
            .I(N__76704));
    Span4Mux_h I__19241 (
            .O(N__76802),
            .I(N__76704));
    LocalMux I__19240 (
            .O(N__76797),
            .I(progRomAddress_0));
    Odrv12 I__19239 (
            .O(N__76792),
            .I(progRomAddress_0));
    LocalMux I__19238 (
            .O(N__76787),
            .I(progRomAddress_0));
    Odrv4 I__19237 (
            .O(N__76784),
            .I(progRomAddress_0));
    Odrv4 I__19236 (
            .O(N__76775),
            .I(progRomAddress_0));
    LocalMux I__19235 (
            .O(N__76762),
            .I(progRomAddress_0));
    LocalMux I__19234 (
            .O(N__76753),
            .I(progRomAddress_0));
    LocalMux I__19233 (
            .O(N__76746),
            .I(progRomAddress_0));
    Odrv4 I__19232 (
            .O(N__76743),
            .I(progRomAddress_0));
    LocalMux I__19231 (
            .O(N__76732),
            .I(progRomAddress_0));
    Odrv4 I__19230 (
            .O(N__76723),
            .I(progRomAddress_0));
    Odrv4 I__19229 (
            .O(N__76704),
            .I(progRomAddress_0));
    InMux I__19228 (
            .O(N__76679),
            .I(N__76676));
    LocalMux I__19227 (
            .O(N__76676),
            .I(N__76673));
    Span4Mux_v I__19226 (
            .O(N__76673),
            .I(N__76670));
    Span4Mux_h I__19225 (
            .O(N__76670),
            .I(N__76667));
    Odrv4 I__19224 (
            .O(N__76667),
            .I(\PROM.ROMDATA.m338_bm ));
    CascadeMux I__19223 (
            .O(N__76664),
            .I(\PROM.ROMDATA.m338_am_cascade_ ));
    InMux I__19222 (
            .O(N__76661),
            .I(N__76658));
    LocalMux I__19221 (
            .O(N__76658),
            .I(\PROM.ROMDATA.m338_ns ));
    InMux I__19220 (
            .O(N__76655),
            .I(N__76652));
    LocalMux I__19219 (
            .O(N__76652),
            .I(N__76649));
    Span4Mux_h I__19218 (
            .O(N__76649),
            .I(N__76645));
    InMux I__19217 (
            .O(N__76648),
            .I(N__76642));
    Odrv4 I__19216 (
            .O(N__76645),
            .I(\PROM.ROMDATA.m246 ));
    LocalMux I__19215 (
            .O(N__76642),
            .I(\PROM.ROMDATA.m246 ));
    InMux I__19214 (
            .O(N__76637),
            .I(N__76626));
    InMux I__19213 (
            .O(N__76636),
            .I(N__76626));
    InMux I__19212 (
            .O(N__76635),
            .I(N__76626));
    CascadeMux I__19211 (
            .O(N__76634),
            .I(N__76620));
    InMux I__19210 (
            .O(N__76633),
            .I(N__76613));
    LocalMux I__19209 (
            .O(N__76626),
            .I(N__76610));
    InMux I__19208 (
            .O(N__76625),
            .I(N__76597));
    InMux I__19207 (
            .O(N__76624),
            .I(N__76594));
    CascadeMux I__19206 (
            .O(N__76623),
            .I(N__76588));
    InMux I__19205 (
            .O(N__76620),
            .I(N__76580));
    CascadeMux I__19204 (
            .O(N__76619),
            .I(N__76576));
    InMux I__19203 (
            .O(N__76618),
            .I(N__76566));
    InMux I__19202 (
            .O(N__76617),
            .I(N__76563));
    CascadeMux I__19201 (
            .O(N__76616),
            .I(N__76560));
    LocalMux I__19200 (
            .O(N__76613),
            .I(N__76554));
    Span4Mux_v I__19199 (
            .O(N__76610),
            .I(N__76554));
    InMux I__19198 (
            .O(N__76609),
            .I(N__76551));
    InMux I__19197 (
            .O(N__76608),
            .I(N__76546));
    InMux I__19196 (
            .O(N__76607),
            .I(N__76546));
    InMux I__19195 (
            .O(N__76606),
            .I(N__76541));
    InMux I__19194 (
            .O(N__76605),
            .I(N__76541));
    InMux I__19193 (
            .O(N__76604),
            .I(N__76536));
    InMux I__19192 (
            .O(N__76603),
            .I(N__76536));
    CascadeMux I__19191 (
            .O(N__76602),
            .I(N__76523));
    CascadeMux I__19190 (
            .O(N__76601),
            .I(N__76519));
    InMux I__19189 (
            .O(N__76600),
            .I(N__76516));
    LocalMux I__19188 (
            .O(N__76597),
            .I(N__76513));
    LocalMux I__19187 (
            .O(N__76594),
            .I(N__76510));
    InMux I__19186 (
            .O(N__76593),
            .I(N__76507));
    InMux I__19185 (
            .O(N__76592),
            .I(N__76504));
    InMux I__19184 (
            .O(N__76591),
            .I(N__76501));
    InMux I__19183 (
            .O(N__76588),
            .I(N__76493));
    InMux I__19182 (
            .O(N__76587),
            .I(N__76493));
    InMux I__19181 (
            .O(N__76586),
            .I(N__76486));
    InMux I__19180 (
            .O(N__76585),
            .I(N__76486));
    InMux I__19179 (
            .O(N__76584),
            .I(N__76486));
    InMux I__19178 (
            .O(N__76583),
            .I(N__76476));
    LocalMux I__19177 (
            .O(N__76580),
            .I(N__76467));
    CascadeMux I__19176 (
            .O(N__76579),
            .I(N__76464));
    InMux I__19175 (
            .O(N__76576),
            .I(N__76455));
    InMux I__19174 (
            .O(N__76575),
            .I(N__76449));
    InMux I__19173 (
            .O(N__76574),
            .I(N__76449));
    InMux I__19172 (
            .O(N__76573),
            .I(N__76441));
    InMux I__19171 (
            .O(N__76572),
            .I(N__76441));
    InMux I__19170 (
            .O(N__76571),
            .I(N__76434));
    InMux I__19169 (
            .O(N__76570),
            .I(N__76434));
    InMux I__19168 (
            .O(N__76569),
            .I(N__76434));
    LocalMux I__19167 (
            .O(N__76566),
            .I(N__76429));
    LocalMux I__19166 (
            .O(N__76563),
            .I(N__76429));
    InMux I__19165 (
            .O(N__76560),
            .I(N__76424));
    InMux I__19164 (
            .O(N__76559),
            .I(N__76424));
    Span4Mux_h I__19163 (
            .O(N__76554),
            .I(N__76421));
    LocalMux I__19162 (
            .O(N__76551),
            .I(N__76414));
    LocalMux I__19161 (
            .O(N__76546),
            .I(N__76414));
    LocalMux I__19160 (
            .O(N__76541),
            .I(N__76414));
    LocalMux I__19159 (
            .O(N__76536),
            .I(N__76411));
    InMux I__19158 (
            .O(N__76535),
            .I(N__76406));
    InMux I__19157 (
            .O(N__76534),
            .I(N__76406));
    InMux I__19156 (
            .O(N__76533),
            .I(N__76396));
    InMux I__19155 (
            .O(N__76532),
            .I(N__76396));
    InMux I__19154 (
            .O(N__76531),
            .I(N__76396));
    InMux I__19153 (
            .O(N__76530),
            .I(N__76391));
    InMux I__19152 (
            .O(N__76529),
            .I(N__76391));
    InMux I__19151 (
            .O(N__76528),
            .I(N__76388));
    InMux I__19150 (
            .O(N__76527),
            .I(N__76381));
    InMux I__19149 (
            .O(N__76526),
            .I(N__76381));
    InMux I__19148 (
            .O(N__76523),
            .I(N__76381));
    InMux I__19147 (
            .O(N__76522),
            .I(N__76378));
    InMux I__19146 (
            .O(N__76519),
            .I(N__76375));
    LocalMux I__19145 (
            .O(N__76516),
            .I(N__76369));
    Span4Mux_h I__19144 (
            .O(N__76513),
            .I(N__76362));
    Span4Mux_v I__19143 (
            .O(N__76510),
            .I(N__76362));
    LocalMux I__19142 (
            .O(N__76507),
            .I(N__76362));
    LocalMux I__19141 (
            .O(N__76504),
            .I(N__76357));
    LocalMux I__19140 (
            .O(N__76501),
            .I(N__76357));
    InMux I__19139 (
            .O(N__76500),
            .I(N__76354));
    InMux I__19138 (
            .O(N__76499),
            .I(N__76351));
    CascadeMux I__19137 (
            .O(N__76498),
            .I(N__76346));
    LocalMux I__19136 (
            .O(N__76493),
            .I(N__76341));
    LocalMux I__19135 (
            .O(N__76486),
            .I(N__76341));
    InMux I__19134 (
            .O(N__76485),
            .I(N__76336));
    InMux I__19133 (
            .O(N__76484),
            .I(N__76336));
    InMux I__19132 (
            .O(N__76483),
            .I(N__76331));
    InMux I__19131 (
            .O(N__76482),
            .I(N__76331));
    InMux I__19130 (
            .O(N__76481),
            .I(N__76326));
    InMux I__19129 (
            .O(N__76480),
            .I(N__76326));
    InMux I__19128 (
            .O(N__76479),
            .I(N__76323));
    LocalMux I__19127 (
            .O(N__76476),
            .I(N__76318));
    InMux I__19126 (
            .O(N__76475),
            .I(N__76313));
    InMux I__19125 (
            .O(N__76474),
            .I(N__76313));
    InMux I__19124 (
            .O(N__76473),
            .I(N__76310));
    InMux I__19123 (
            .O(N__76472),
            .I(N__76305));
    InMux I__19122 (
            .O(N__76471),
            .I(N__76305));
    InMux I__19121 (
            .O(N__76470),
            .I(N__76302));
    Span4Mux_h I__19120 (
            .O(N__76467),
            .I(N__76299));
    InMux I__19119 (
            .O(N__76464),
            .I(N__76294));
    InMux I__19118 (
            .O(N__76463),
            .I(N__76294));
    CascadeMux I__19117 (
            .O(N__76462),
            .I(N__76288));
    InMux I__19116 (
            .O(N__76461),
            .I(N__76277));
    InMux I__19115 (
            .O(N__76460),
            .I(N__76277));
    InMux I__19114 (
            .O(N__76459),
            .I(N__76277));
    InMux I__19113 (
            .O(N__76458),
            .I(N__76277));
    LocalMux I__19112 (
            .O(N__76455),
            .I(N__76274));
    CascadeMux I__19111 (
            .O(N__76454),
            .I(N__76265));
    LocalMux I__19110 (
            .O(N__76449),
            .I(N__76258));
    InMux I__19109 (
            .O(N__76448),
            .I(N__76251));
    InMux I__19108 (
            .O(N__76447),
            .I(N__76251));
    InMux I__19107 (
            .O(N__76446),
            .I(N__76251));
    LocalMux I__19106 (
            .O(N__76441),
            .I(N__76248));
    LocalMux I__19105 (
            .O(N__76434),
            .I(N__76241));
    Span4Mux_v I__19104 (
            .O(N__76429),
            .I(N__76241));
    LocalMux I__19103 (
            .O(N__76424),
            .I(N__76241));
    Span4Mux_h I__19102 (
            .O(N__76421),
            .I(N__76232));
    Span4Mux_v I__19101 (
            .O(N__76414),
            .I(N__76232));
    Span4Mux_v I__19100 (
            .O(N__76411),
            .I(N__76232));
    LocalMux I__19099 (
            .O(N__76406),
            .I(N__76232));
    InMux I__19098 (
            .O(N__76405),
            .I(N__76225));
    InMux I__19097 (
            .O(N__76404),
            .I(N__76225));
    InMux I__19096 (
            .O(N__76403),
            .I(N__76225));
    LocalMux I__19095 (
            .O(N__76396),
            .I(N__76222));
    LocalMux I__19094 (
            .O(N__76391),
            .I(N__76215));
    LocalMux I__19093 (
            .O(N__76388),
            .I(N__76215));
    LocalMux I__19092 (
            .O(N__76381),
            .I(N__76215));
    LocalMux I__19091 (
            .O(N__76378),
            .I(N__76210));
    LocalMux I__19090 (
            .O(N__76375),
            .I(N__76210));
    InMux I__19089 (
            .O(N__76374),
            .I(N__76203));
    InMux I__19088 (
            .O(N__76373),
            .I(N__76203));
    InMux I__19087 (
            .O(N__76372),
            .I(N__76203));
    Span4Mux_v I__19086 (
            .O(N__76369),
            .I(N__76192));
    Span4Mux_h I__19085 (
            .O(N__76362),
            .I(N__76192));
    Span4Mux_v I__19084 (
            .O(N__76357),
            .I(N__76192));
    LocalMux I__19083 (
            .O(N__76354),
            .I(N__76192));
    LocalMux I__19082 (
            .O(N__76351),
            .I(N__76192));
    InMux I__19081 (
            .O(N__76350),
            .I(N__76185));
    InMux I__19080 (
            .O(N__76349),
            .I(N__76185));
    InMux I__19079 (
            .O(N__76346),
            .I(N__76185));
    Span4Mux_h I__19078 (
            .O(N__76341),
            .I(N__76174));
    LocalMux I__19077 (
            .O(N__76336),
            .I(N__76174));
    LocalMux I__19076 (
            .O(N__76331),
            .I(N__76174));
    LocalMux I__19075 (
            .O(N__76326),
            .I(N__76174));
    LocalMux I__19074 (
            .O(N__76323),
            .I(N__76174));
    InMux I__19073 (
            .O(N__76322),
            .I(N__76168));
    InMux I__19072 (
            .O(N__76321),
            .I(N__76168));
    Span4Mux_h I__19071 (
            .O(N__76318),
            .I(N__76159));
    LocalMux I__19070 (
            .O(N__76313),
            .I(N__76159));
    LocalMux I__19069 (
            .O(N__76310),
            .I(N__76159));
    LocalMux I__19068 (
            .O(N__76305),
            .I(N__76159));
    LocalMux I__19067 (
            .O(N__76302),
            .I(N__76152));
    Span4Mux_v I__19066 (
            .O(N__76299),
            .I(N__76152));
    LocalMux I__19065 (
            .O(N__76294),
            .I(N__76152));
    InMux I__19064 (
            .O(N__76293),
            .I(N__76145));
    InMux I__19063 (
            .O(N__76292),
            .I(N__76145));
    InMux I__19062 (
            .O(N__76291),
            .I(N__76145));
    InMux I__19061 (
            .O(N__76288),
            .I(N__76142));
    InMux I__19060 (
            .O(N__76287),
            .I(N__76139));
    InMux I__19059 (
            .O(N__76286),
            .I(N__76136));
    LocalMux I__19058 (
            .O(N__76277),
            .I(N__76131));
    Span4Mux_h I__19057 (
            .O(N__76274),
            .I(N__76131));
    InMux I__19056 (
            .O(N__76273),
            .I(N__76128));
    InMux I__19055 (
            .O(N__76272),
            .I(N__76123));
    InMux I__19054 (
            .O(N__76271),
            .I(N__76123));
    InMux I__19053 (
            .O(N__76270),
            .I(N__76118));
    InMux I__19052 (
            .O(N__76269),
            .I(N__76118));
    InMux I__19051 (
            .O(N__76268),
            .I(N__76113));
    InMux I__19050 (
            .O(N__76265),
            .I(N__76113));
    InMux I__19049 (
            .O(N__76264),
            .I(N__76110));
    InMux I__19048 (
            .O(N__76263),
            .I(N__76103));
    InMux I__19047 (
            .O(N__76262),
            .I(N__76103));
    InMux I__19046 (
            .O(N__76261),
            .I(N__76103));
    Span4Mux_v I__19045 (
            .O(N__76258),
            .I(N__76098));
    LocalMux I__19044 (
            .O(N__76251),
            .I(N__76098));
    Span4Mux_v I__19043 (
            .O(N__76248),
            .I(N__76089));
    Span4Mux_h I__19042 (
            .O(N__76241),
            .I(N__76089));
    Span4Mux_h I__19041 (
            .O(N__76232),
            .I(N__76089));
    LocalMux I__19040 (
            .O(N__76225),
            .I(N__76089));
    Span4Mux_v I__19039 (
            .O(N__76222),
            .I(N__76074));
    Span4Mux_v I__19038 (
            .O(N__76215),
            .I(N__76074));
    Span4Mux_v I__19037 (
            .O(N__76210),
            .I(N__76074));
    LocalMux I__19036 (
            .O(N__76203),
            .I(N__76074));
    Span4Mux_h I__19035 (
            .O(N__76192),
            .I(N__76074));
    LocalMux I__19034 (
            .O(N__76185),
            .I(N__76074));
    Span4Mux_v I__19033 (
            .O(N__76174),
            .I(N__76074));
    InMux I__19032 (
            .O(N__76173),
            .I(N__76071));
    LocalMux I__19031 (
            .O(N__76168),
            .I(N__76062));
    Span4Mux_v I__19030 (
            .O(N__76159),
            .I(N__76062));
    Span4Mux_h I__19029 (
            .O(N__76152),
            .I(N__76062));
    LocalMux I__19028 (
            .O(N__76145),
            .I(N__76062));
    LocalMux I__19027 (
            .O(N__76142),
            .I(N__76059));
    LocalMux I__19026 (
            .O(N__76139),
            .I(progRomAddress_4));
    LocalMux I__19025 (
            .O(N__76136),
            .I(progRomAddress_4));
    Odrv4 I__19024 (
            .O(N__76131),
            .I(progRomAddress_4));
    LocalMux I__19023 (
            .O(N__76128),
            .I(progRomAddress_4));
    LocalMux I__19022 (
            .O(N__76123),
            .I(progRomAddress_4));
    LocalMux I__19021 (
            .O(N__76118),
            .I(progRomAddress_4));
    LocalMux I__19020 (
            .O(N__76113),
            .I(progRomAddress_4));
    LocalMux I__19019 (
            .O(N__76110),
            .I(progRomAddress_4));
    LocalMux I__19018 (
            .O(N__76103),
            .I(progRomAddress_4));
    Odrv4 I__19017 (
            .O(N__76098),
            .I(progRomAddress_4));
    Odrv4 I__19016 (
            .O(N__76089),
            .I(progRomAddress_4));
    Odrv4 I__19015 (
            .O(N__76074),
            .I(progRomAddress_4));
    LocalMux I__19014 (
            .O(N__76071),
            .I(progRomAddress_4));
    Odrv4 I__19013 (
            .O(N__76062),
            .I(progRomAddress_4));
    Odrv12 I__19012 (
            .O(N__76059),
            .I(progRomAddress_4));
    CascadeMux I__19011 (
            .O(N__76028),
            .I(N__76025));
    InMux I__19010 (
            .O(N__76025),
            .I(N__76022));
    LocalMux I__19009 (
            .O(N__76022),
            .I(N__76019));
    Odrv4 I__19008 (
            .O(N__76019),
            .I(\PROM.ROMDATA.m341_ns_1 ));
    CascadeMux I__19007 (
            .O(N__76016),
            .I(N__76012));
    InMux I__19006 (
            .O(N__76015),
            .I(N__76005));
    InMux I__19005 (
            .O(N__76012),
            .I(N__75997));
    InMux I__19004 (
            .O(N__76011),
            .I(N__75997));
    CascadeMux I__19003 (
            .O(N__76010),
            .I(N__75987));
    CascadeMux I__19002 (
            .O(N__76009),
            .I(N__75980));
    CascadeMux I__19001 (
            .O(N__76008),
            .I(N__75977));
    LocalMux I__19000 (
            .O(N__76005),
            .I(N__75974));
    CascadeMux I__18999 (
            .O(N__76004),
            .I(N__75970));
    CascadeMux I__18998 (
            .O(N__76003),
            .I(N__75956));
    CascadeMux I__18997 (
            .O(N__76002),
            .I(N__75951));
    LocalMux I__18996 (
            .O(N__75997),
            .I(N__75947));
    InMux I__18995 (
            .O(N__75996),
            .I(N__75942));
    InMux I__18994 (
            .O(N__75995),
            .I(N__75942));
    CascadeMux I__18993 (
            .O(N__75994),
            .I(N__75935));
    CascadeMux I__18992 (
            .O(N__75993),
            .I(N__75929));
    CascadeMux I__18991 (
            .O(N__75992),
            .I(N__75926));
    CascadeMux I__18990 (
            .O(N__75991),
            .I(N__75923));
    CascadeMux I__18989 (
            .O(N__75990),
            .I(N__75920));
    InMux I__18988 (
            .O(N__75987),
            .I(N__75896));
    CascadeMux I__18987 (
            .O(N__75986),
            .I(N__75893));
    InMux I__18986 (
            .O(N__75985),
            .I(N__75882));
    CascadeMux I__18985 (
            .O(N__75984),
            .I(N__75876));
    InMux I__18984 (
            .O(N__75983),
            .I(N__75871));
    InMux I__18983 (
            .O(N__75980),
            .I(N__75871));
    InMux I__18982 (
            .O(N__75977),
            .I(N__75868));
    Span4Mux_v I__18981 (
            .O(N__75974),
            .I(N__75865));
    InMux I__18980 (
            .O(N__75973),
            .I(N__75860));
    InMux I__18979 (
            .O(N__75970),
            .I(N__75860));
    InMux I__18978 (
            .O(N__75969),
            .I(N__75857));
    CascadeMux I__18977 (
            .O(N__75968),
            .I(N__75853));
    CascadeMux I__18976 (
            .O(N__75967),
            .I(N__75848));
    CascadeMux I__18975 (
            .O(N__75966),
            .I(N__75843));
    CascadeMux I__18974 (
            .O(N__75965),
            .I(N__75840));
    CascadeMux I__18973 (
            .O(N__75964),
            .I(N__75836));
    CascadeMux I__18972 (
            .O(N__75963),
            .I(N__75833));
    CascadeMux I__18971 (
            .O(N__75962),
            .I(N__75825));
    CascadeMux I__18970 (
            .O(N__75961),
            .I(N__75822));
    CascadeMux I__18969 (
            .O(N__75960),
            .I(N__75818));
    CascadeMux I__18968 (
            .O(N__75959),
            .I(N__75811));
    InMux I__18967 (
            .O(N__75956),
            .I(N__75805));
    CascadeMux I__18966 (
            .O(N__75955),
            .I(N__75801));
    CascadeMux I__18965 (
            .O(N__75954),
            .I(N__75796));
    InMux I__18964 (
            .O(N__75951),
            .I(N__75792));
    CascadeMux I__18963 (
            .O(N__75950),
            .I(N__75786));
    Span4Mux_h I__18962 (
            .O(N__75947),
            .I(N__75781));
    LocalMux I__18961 (
            .O(N__75942),
            .I(N__75781));
    InMux I__18960 (
            .O(N__75941),
            .I(N__75770));
    InMux I__18959 (
            .O(N__75940),
            .I(N__75770));
    InMux I__18958 (
            .O(N__75939),
            .I(N__75770));
    InMux I__18957 (
            .O(N__75938),
            .I(N__75770));
    InMux I__18956 (
            .O(N__75935),
            .I(N__75770));
    InMux I__18955 (
            .O(N__75934),
            .I(N__75763));
    InMux I__18954 (
            .O(N__75933),
            .I(N__75763));
    InMux I__18953 (
            .O(N__75932),
            .I(N__75763));
    InMux I__18952 (
            .O(N__75929),
            .I(N__75754));
    InMux I__18951 (
            .O(N__75926),
            .I(N__75754));
    InMux I__18950 (
            .O(N__75923),
            .I(N__75754));
    InMux I__18949 (
            .O(N__75920),
            .I(N__75754));
    CascadeMux I__18948 (
            .O(N__75919),
            .I(N__75751));
    CascadeMux I__18947 (
            .O(N__75918),
            .I(N__75747));
    CascadeMux I__18946 (
            .O(N__75917),
            .I(N__75743));
    CascadeMux I__18945 (
            .O(N__75916),
            .I(N__75740));
    CascadeMux I__18944 (
            .O(N__75915),
            .I(N__75737));
    CascadeMux I__18943 (
            .O(N__75914),
            .I(N__75733));
    CascadeMux I__18942 (
            .O(N__75913),
            .I(N__75730));
    CascadeMux I__18941 (
            .O(N__75912),
            .I(N__75727));
    CascadeMux I__18940 (
            .O(N__75911),
            .I(N__75722));
    CascadeMux I__18939 (
            .O(N__75910),
            .I(N__75715));
    CascadeMux I__18938 (
            .O(N__75909),
            .I(N__75712));
    InMux I__18937 (
            .O(N__75908),
            .I(N__75705));
    InMux I__18936 (
            .O(N__75907),
            .I(N__75702));
    InMux I__18935 (
            .O(N__75906),
            .I(N__75695));
    InMux I__18934 (
            .O(N__75905),
            .I(N__75695));
    InMux I__18933 (
            .O(N__75904),
            .I(N__75695));
    CascadeMux I__18932 (
            .O(N__75903),
            .I(N__75692));
    CascadeMux I__18931 (
            .O(N__75902),
            .I(N__75689));
    CascadeMux I__18930 (
            .O(N__75901),
            .I(N__75685));
    CascadeMux I__18929 (
            .O(N__75900),
            .I(N__75681));
    CascadeMux I__18928 (
            .O(N__75899),
            .I(N__75677));
    LocalMux I__18927 (
            .O(N__75896),
            .I(N__75673));
    InMux I__18926 (
            .O(N__75893),
            .I(N__75665));
    InMux I__18925 (
            .O(N__75892),
            .I(N__75660));
    InMux I__18924 (
            .O(N__75891),
            .I(N__75660));
    CascadeMux I__18923 (
            .O(N__75890),
            .I(N__75656));
    CascadeMux I__18922 (
            .O(N__75889),
            .I(N__75650));
    CascadeMux I__18921 (
            .O(N__75888),
            .I(N__75647));
    CascadeMux I__18920 (
            .O(N__75887),
            .I(N__75642));
    CascadeMux I__18919 (
            .O(N__75886),
            .I(N__75639));
    CascadeMux I__18918 (
            .O(N__75885),
            .I(N__75632));
    LocalMux I__18917 (
            .O(N__75882),
            .I(N__75627));
    InMux I__18916 (
            .O(N__75881),
            .I(N__75620));
    InMux I__18915 (
            .O(N__75880),
            .I(N__75620));
    InMux I__18914 (
            .O(N__75879),
            .I(N__75620));
    InMux I__18913 (
            .O(N__75876),
            .I(N__75616));
    LocalMux I__18912 (
            .O(N__75871),
            .I(N__75606));
    LocalMux I__18911 (
            .O(N__75868),
            .I(N__75606));
    Span4Mux_h I__18910 (
            .O(N__75865),
            .I(N__75599));
    LocalMux I__18909 (
            .O(N__75860),
            .I(N__75599));
    LocalMux I__18908 (
            .O(N__75857),
            .I(N__75599));
    InMux I__18907 (
            .O(N__75856),
            .I(N__75594));
    InMux I__18906 (
            .O(N__75853),
            .I(N__75587));
    InMux I__18905 (
            .O(N__75852),
            .I(N__75587));
    InMux I__18904 (
            .O(N__75851),
            .I(N__75587));
    InMux I__18903 (
            .O(N__75848),
            .I(N__75580));
    InMux I__18902 (
            .O(N__75847),
            .I(N__75580));
    InMux I__18901 (
            .O(N__75846),
            .I(N__75580));
    InMux I__18900 (
            .O(N__75843),
            .I(N__75577));
    InMux I__18899 (
            .O(N__75840),
            .I(N__75570));
    InMux I__18898 (
            .O(N__75839),
            .I(N__75570));
    InMux I__18897 (
            .O(N__75836),
            .I(N__75570));
    InMux I__18896 (
            .O(N__75833),
            .I(N__75561));
    InMux I__18895 (
            .O(N__75832),
            .I(N__75561));
    InMux I__18894 (
            .O(N__75831),
            .I(N__75561));
    InMux I__18893 (
            .O(N__75830),
            .I(N__75561));
    InMux I__18892 (
            .O(N__75829),
            .I(N__75556));
    InMux I__18891 (
            .O(N__75828),
            .I(N__75556));
    InMux I__18890 (
            .O(N__75825),
            .I(N__75551));
    InMux I__18889 (
            .O(N__75822),
            .I(N__75551));
    InMux I__18888 (
            .O(N__75821),
            .I(N__75546));
    InMux I__18887 (
            .O(N__75818),
            .I(N__75546));
    InMux I__18886 (
            .O(N__75817),
            .I(N__75541));
    InMux I__18885 (
            .O(N__75816),
            .I(N__75541));
    InMux I__18884 (
            .O(N__75815),
            .I(N__75535));
    CascadeMux I__18883 (
            .O(N__75814),
            .I(N__75530));
    InMux I__18882 (
            .O(N__75811),
            .I(N__75521));
    InMux I__18881 (
            .O(N__75810),
            .I(N__75521));
    InMux I__18880 (
            .O(N__75809),
            .I(N__75516));
    InMux I__18879 (
            .O(N__75808),
            .I(N__75516));
    LocalMux I__18878 (
            .O(N__75805),
            .I(N__75513));
    InMux I__18877 (
            .O(N__75804),
            .I(N__75502));
    InMux I__18876 (
            .O(N__75801),
            .I(N__75502));
    InMux I__18875 (
            .O(N__75800),
            .I(N__75502));
    InMux I__18874 (
            .O(N__75799),
            .I(N__75502));
    InMux I__18873 (
            .O(N__75796),
            .I(N__75502));
    CascadeMux I__18872 (
            .O(N__75795),
            .I(N__75496));
    LocalMux I__18871 (
            .O(N__75792),
            .I(N__75493));
    InMux I__18870 (
            .O(N__75791),
            .I(N__75490));
    InMux I__18869 (
            .O(N__75790),
            .I(N__75483));
    InMux I__18868 (
            .O(N__75789),
            .I(N__75483));
    InMux I__18867 (
            .O(N__75786),
            .I(N__75483));
    Span4Mux_h I__18866 (
            .O(N__75781),
            .I(N__75474));
    LocalMux I__18865 (
            .O(N__75770),
            .I(N__75474));
    LocalMux I__18864 (
            .O(N__75763),
            .I(N__75474));
    LocalMux I__18863 (
            .O(N__75754),
            .I(N__75474));
    InMux I__18862 (
            .O(N__75751),
            .I(N__75467));
    InMux I__18861 (
            .O(N__75750),
            .I(N__75467));
    InMux I__18860 (
            .O(N__75747),
            .I(N__75467));
    InMux I__18859 (
            .O(N__75746),
            .I(N__75460));
    InMux I__18858 (
            .O(N__75743),
            .I(N__75460));
    InMux I__18857 (
            .O(N__75740),
            .I(N__75460));
    InMux I__18856 (
            .O(N__75737),
            .I(N__75453));
    InMux I__18855 (
            .O(N__75736),
            .I(N__75453));
    InMux I__18854 (
            .O(N__75733),
            .I(N__75453));
    InMux I__18853 (
            .O(N__75730),
            .I(N__75446));
    InMux I__18852 (
            .O(N__75727),
            .I(N__75446));
    InMux I__18851 (
            .O(N__75726),
            .I(N__75446));
    InMux I__18850 (
            .O(N__75725),
            .I(N__75439));
    InMux I__18849 (
            .O(N__75722),
            .I(N__75439));
    InMux I__18848 (
            .O(N__75721),
            .I(N__75439));
    InMux I__18847 (
            .O(N__75720),
            .I(N__75430));
    InMux I__18846 (
            .O(N__75719),
            .I(N__75430));
    InMux I__18845 (
            .O(N__75718),
            .I(N__75430));
    InMux I__18844 (
            .O(N__75715),
            .I(N__75430));
    InMux I__18843 (
            .O(N__75712),
            .I(N__75425));
    InMux I__18842 (
            .O(N__75711),
            .I(N__75425));
    CascadeMux I__18841 (
            .O(N__75710),
            .I(N__75419));
    CascadeMux I__18840 (
            .O(N__75709),
            .I(N__75416));
    InMux I__18839 (
            .O(N__75708),
            .I(N__75413));
    LocalMux I__18838 (
            .O(N__75705),
            .I(N__75410));
    LocalMux I__18837 (
            .O(N__75702),
            .I(N__75407));
    LocalMux I__18836 (
            .O(N__75695),
            .I(N__75404));
    InMux I__18835 (
            .O(N__75692),
            .I(N__75401));
    InMux I__18834 (
            .O(N__75689),
            .I(N__75394));
    InMux I__18833 (
            .O(N__75688),
            .I(N__75394));
    InMux I__18832 (
            .O(N__75685),
            .I(N__75394));
    InMux I__18831 (
            .O(N__75684),
            .I(N__75385));
    InMux I__18830 (
            .O(N__75681),
            .I(N__75385));
    InMux I__18829 (
            .O(N__75680),
            .I(N__75385));
    InMux I__18828 (
            .O(N__75677),
            .I(N__75385));
    CascadeMux I__18827 (
            .O(N__75676),
            .I(N__75380));
    Span4Mux_h I__18826 (
            .O(N__75673),
            .I(N__75377));
    InMux I__18825 (
            .O(N__75672),
            .I(N__75366));
    InMux I__18824 (
            .O(N__75671),
            .I(N__75366));
    InMux I__18823 (
            .O(N__75670),
            .I(N__75366));
    InMux I__18822 (
            .O(N__75669),
            .I(N__75366));
    InMux I__18821 (
            .O(N__75668),
            .I(N__75366));
    LocalMux I__18820 (
            .O(N__75665),
            .I(N__75361));
    LocalMux I__18819 (
            .O(N__75660),
            .I(N__75361));
    InMux I__18818 (
            .O(N__75659),
            .I(N__75348));
    InMux I__18817 (
            .O(N__75656),
            .I(N__75348));
    InMux I__18816 (
            .O(N__75655),
            .I(N__75348));
    InMux I__18815 (
            .O(N__75654),
            .I(N__75348));
    InMux I__18814 (
            .O(N__75653),
            .I(N__75348));
    InMux I__18813 (
            .O(N__75650),
            .I(N__75348));
    InMux I__18812 (
            .O(N__75647),
            .I(N__75339));
    InMux I__18811 (
            .O(N__75646),
            .I(N__75339));
    InMux I__18810 (
            .O(N__75645),
            .I(N__75339));
    InMux I__18809 (
            .O(N__75642),
            .I(N__75339));
    InMux I__18808 (
            .O(N__75639),
            .I(N__75336));
    InMux I__18807 (
            .O(N__75638),
            .I(N__75329));
    InMux I__18806 (
            .O(N__75637),
            .I(N__75329));
    InMux I__18805 (
            .O(N__75636),
            .I(N__75329));
    InMux I__18804 (
            .O(N__75635),
            .I(N__75320));
    InMux I__18803 (
            .O(N__75632),
            .I(N__75320));
    InMux I__18802 (
            .O(N__75631),
            .I(N__75320));
    InMux I__18801 (
            .O(N__75630),
            .I(N__75320));
    Span4Mux_v I__18800 (
            .O(N__75627),
            .I(N__75317));
    LocalMux I__18799 (
            .O(N__75620),
            .I(N__75314));
    InMux I__18798 (
            .O(N__75619),
            .I(N__75311));
    LocalMux I__18797 (
            .O(N__75616),
            .I(N__75308));
    CascadeMux I__18796 (
            .O(N__75615),
            .I(N__75300));
    CascadeMux I__18795 (
            .O(N__75614),
            .I(N__75296));
    CascadeMux I__18794 (
            .O(N__75613),
            .I(N__75293));
    CascadeMux I__18793 (
            .O(N__75612),
            .I(N__75288));
    CascadeMux I__18792 (
            .O(N__75611),
            .I(N__75284));
    Span4Mux_v I__18791 (
            .O(N__75606),
            .I(N__75280));
    Span4Mux_v I__18790 (
            .O(N__75599),
            .I(N__75277));
    InMux I__18789 (
            .O(N__75598),
            .I(N__75272));
    InMux I__18788 (
            .O(N__75597),
            .I(N__75272));
    LocalMux I__18787 (
            .O(N__75594),
            .I(N__75263));
    LocalMux I__18786 (
            .O(N__75587),
            .I(N__75263));
    LocalMux I__18785 (
            .O(N__75580),
            .I(N__75263));
    LocalMux I__18784 (
            .O(N__75577),
            .I(N__75263));
    LocalMux I__18783 (
            .O(N__75570),
            .I(N__75258));
    LocalMux I__18782 (
            .O(N__75561),
            .I(N__75258));
    LocalMux I__18781 (
            .O(N__75556),
            .I(N__75249));
    LocalMux I__18780 (
            .O(N__75551),
            .I(N__75249));
    LocalMux I__18779 (
            .O(N__75546),
            .I(N__75249));
    LocalMux I__18778 (
            .O(N__75541),
            .I(N__75249));
    CascadeMux I__18777 (
            .O(N__75540),
            .I(N__75244));
    CascadeMux I__18776 (
            .O(N__75539),
            .I(N__75240));
    CascadeMux I__18775 (
            .O(N__75538),
            .I(N__75237));
    LocalMux I__18774 (
            .O(N__75535),
            .I(N__75231));
    InMux I__18773 (
            .O(N__75534),
            .I(N__75224));
    InMux I__18772 (
            .O(N__75533),
            .I(N__75224));
    InMux I__18771 (
            .O(N__75530),
            .I(N__75224));
    InMux I__18770 (
            .O(N__75529),
            .I(N__75215));
    InMux I__18769 (
            .O(N__75528),
            .I(N__75215));
    InMux I__18768 (
            .O(N__75527),
            .I(N__75215));
    InMux I__18767 (
            .O(N__75526),
            .I(N__75215));
    LocalMux I__18766 (
            .O(N__75521),
            .I(N__75212));
    LocalMux I__18765 (
            .O(N__75516),
            .I(N__75205));
    Span4Mux_v I__18764 (
            .O(N__75513),
            .I(N__75205));
    LocalMux I__18763 (
            .O(N__75502),
            .I(N__75205));
    InMux I__18762 (
            .O(N__75501),
            .I(N__75196));
    InMux I__18761 (
            .O(N__75500),
            .I(N__75196));
    InMux I__18760 (
            .O(N__75499),
            .I(N__75196));
    InMux I__18759 (
            .O(N__75496),
            .I(N__75196));
    Span4Mux_h I__18758 (
            .O(N__75493),
            .I(N__75179));
    LocalMux I__18757 (
            .O(N__75490),
            .I(N__75179));
    LocalMux I__18756 (
            .O(N__75483),
            .I(N__75179));
    Span4Mux_v I__18755 (
            .O(N__75474),
            .I(N__75179));
    LocalMux I__18754 (
            .O(N__75467),
            .I(N__75179));
    LocalMux I__18753 (
            .O(N__75460),
            .I(N__75179));
    LocalMux I__18752 (
            .O(N__75453),
            .I(N__75179));
    LocalMux I__18751 (
            .O(N__75446),
            .I(N__75179));
    LocalMux I__18750 (
            .O(N__75439),
            .I(N__75172));
    LocalMux I__18749 (
            .O(N__75430),
            .I(N__75172));
    LocalMux I__18748 (
            .O(N__75425),
            .I(N__75172));
    InMux I__18747 (
            .O(N__75424),
            .I(N__75161));
    InMux I__18746 (
            .O(N__75423),
            .I(N__75161));
    InMux I__18745 (
            .O(N__75422),
            .I(N__75161));
    InMux I__18744 (
            .O(N__75419),
            .I(N__75161));
    InMux I__18743 (
            .O(N__75416),
            .I(N__75161));
    LocalMux I__18742 (
            .O(N__75413),
            .I(N__75158));
    Span4Mux_h I__18741 (
            .O(N__75410),
            .I(N__75151));
    Span4Mux_v I__18740 (
            .O(N__75407),
            .I(N__75151));
    Span4Mux_h I__18739 (
            .O(N__75404),
            .I(N__75151));
    LocalMux I__18738 (
            .O(N__75401),
            .I(N__75144));
    LocalMux I__18737 (
            .O(N__75394),
            .I(N__75144));
    LocalMux I__18736 (
            .O(N__75385),
            .I(N__75144));
    InMux I__18735 (
            .O(N__75384),
            .I(N__75137));
    InMux I__18734 (
            .O(N__75383),
            .I(N__75137));
    InMux I__18733 (
            .O(N__75380),
            .I(N__75137));
    Span4Mux_v I__18732 (
            .O(N__75377),
            .I(N__75126));
    LocalMux I__18731 (
            .O(N__75366),
            .I(N__75126));
    Span4Mux_h I__18730 (
            .O(N__75361),
            .I(N__75126));
    LocalMux I__18729 (
            .O(N__75348),
            .I(N__75126));
    LocalMux I__18728 (
            .O(N__75339),
            .I(N__75126));
    LocalMux I__18727 (
            .O(N__75336),
            .I(N__75123));
    LocalMux I__18726 (
            .O(N__75329),
            .I(N__75118));
    LocalMux I__18725 (
            .O(N__75320),
            .I(N__75118));
    Span4Mux_h I__18724 (
            .O(N__75317),
            .I(N__75109));
    Span4Mux_v I__18723 (
            .O(N__75314),
            .I(N__75109));
    LocalMux I__18722 (
            .O(N__75311),
            .I(N__75109));
    Span4Mux_v I__18721 (
            .O(N__75308),
            .I(N__75109));
    InMux I__18720 (
            .O(N__75307),
            .I(N__75106));
    InMux I__18719 (
            .O(N__75306),
            .I(N__75101));
    InMux I__18718 (
            .O(N__75305),
            .I(N__75101));
    InMux I__18717 (
            .O(N__75304),
            .I(N__75090));
    InMux I__18716 (
            .O(N__75303),
            .I(N__75090));
    InMux I__18715 (
            .O(N__75300),
            .I(N__75090));
    InMux I__18714 (
            .O(N__75299),
            .I(N__75090));
    InMux I__18713 (
            .O(N__75296),
            .I(N__75090));
    InMux I__18712 (
            .O(N__75293),
            .I(N__75083));
    InMux I__18711 (
            .O(N__75292),
            .I(N__75083));
    InMux I__18710 (
            .O(N__75291),
            .I(N__75083));
    InMux I__18709 (
            .O(N__75288),
            .I(N__75074));
    InMux I__18708 (
            .O(N__75287),
            .I(N__75074));
    InMux I__18707 (
            .O(N__75284),
            .I(N__75074));
    InMux I__18706 (
            .O(N__75283),
            .I(N__75074));
    Span4Mux_h I__18705 (
            .O(N__75280),
            .I(N__75061));
    Span4Mux_h I__18704 (
            .O(N__75277),
            .I(N__75061));
    LocalMux I__18703 (
            .O(N__75272),
            .I(N__75061));
    Span4Mux_v I__18702 (
            .O(N__75263),
            .I(N__75061));
    Span4Mux_v I__18701 (
            .O(N__75258),
            .I(N__75061));
    Span4Mux_v I__18700 (
            .O(N__75249),
            .I(N__75061));
    InMux I__18699 (
            .O(N__75248),
            .I(N__75050));
    InMux I__18698 (
            .O(N__75247),
            .I(N__75050));
    InMux I__18697 (
            .O(N__75244),
            .I(N__75050));
    InMux I__18696 (
            .O(N__75243),
            .I(N__75050));
    InMux I__18695 (
            .O(N__75240),
            .I(N__75050));
    InMux I__18694 (
            .O(N__75237),
            .I(N__75041));
    InMux I__18693 (
            .O(N__75236),
            .I(N__75041));
    InMux I__18692 (
            .O(N__75235),
            .I(N__75041));
    InMux I__18691 (
            .O(N__75234),
            .I(N__75041));
    Span4Mux_h I__18690 (
            .O(N__75231),
            .I(N__75034));
    LocalMux I__18689 (
            .O(N__75224),
            .I(N__75034));
    LocalMux I__18688 (
            .O(N__75215),
            .I(N__75034));
    Span4Mux_h I__18687 (
            .O(N__75212),
            .I(N__75021));
    Span4Mux_v I__18686 (
            .O(N__75205),
            .I(N__75021));
    LocalMux I__18685 (
            .O(N__75196),
            .I(N__75021));
    Span4Mux_v I__18684 (
            .O(N__75179),
            .I(N__75021));
    Span4Mux_v I__18683 (
            .O(N__75172),
            .I(N__75021));
    LocalMux I__18682 (
            .O(N__75161),
            .I(N__75021));
    Span4Mux_h I__18681 (
            .O(N__75158),
            .I(N__75010));
    Span4Mux_h I__18680 (
            .O(N__75151),
            .I(N__75010));
    Span4Mux_h I__18679 (
            .O(N__75144),
            .I(N__75010));
    LocalMux I__18678 (
            .O(N__75137),
            .I(N__75010));
    Span4Mux_h I__18677 (
            .O(N__75126),
            .I(N__75010));
    Span4Mux_h I__18676 (
            .O(N__75123),
            .I(N__75003));
    Span4Mux_h I__18675 (
            .O(N__75118),
            .I(N__75003));
    Span4Mux_h I__18674 (
            .O(N__75109),
            .I(N__75003));
    LocalMux I__18673 (
            .O(N__75106),
            .I(progRomAddress_3));
    LocalMux I__18672 (
            .O(N__75101),
            .I(progRomAddress_3));
    LocalMux I__18671 (
            .O(N__75090),
            .I(progRomAddress_3));
    LocalMux I__18670 (
            .O(N__75083),
            .I(progRomAddress_3));
    LocalMux I__18669 (
            .O(N__75074),
            .I(progRomAddress_3));
    Odrv4 I__18668 (
            .O(N__75061),
            .I(progRomAddress_3));
    LocalMux I__18667 (
            .O(N__75050),
            .I(progRomAddress_3));
    LocalMux I__18666 (
            .O(N__75041),
            .I(progRomAddress_3));
    Odrv4 I__18665 (
            .O(N__75034),
            .I(progRomAddress_3));
    Odrv4 I__18664 (
            .O(N__75021),
            .I(progRomAddress_3));
    Odrv4 I__18663 (
            .O(N__75010),
            .I(progRomAddress_3));
    Odrv4 I__18662 (
            .O(N__75003),
            .I(progRomAddress_3));
    InMux I__18661 (
            .O(N__74978),
            .I(N__74975));
    LocalMux I__18660 (
            .O(N__74975),
            .I(\PROM.ROMDATA.m341_ns ));
    InMux I__18659 (
            .O(N__74972),
            .I(N__74969));
    LocalMux I__18658 (
            .O(N__74969),
            .I(N__74966));
    Odrv4 I__18657 (
            .O(N__74966),
            .I(\PROM.ROMDATA.m347 ));
    InMux I__18656 (
            .O(N__74963),
            .I(N__74959));
    InMux I__18655 (
            .O(N__74962),
            .I(N__74956));
    LocalMux I__18654 (
            .O(N__74959),
            .I(N__74953));
    LocalMux I__18653 (
            .O(N__74956),
            .I(N__74950));
    Odrv4 I__18652 (
            .O(N__74953),
            .I(\PROM.ROMDATA.m112 ));
    Odrv4 I__18651 (
            .O(N__74950),
            .I(\PROM.ROMDATA.m112 ));
    InMux I__18650 (
            .O(N__74945),
            .I(N__74942));
    LocalMux I__18649 (
            .O(N__74942),
            .I(\PROM.ROMDATA.m349_am ));
    CascadeMux I__18648 (
            .O(N__74939),
            .I(\PROM.ROMDATA.m349_bm_cascade_ ));
    InMux I__18647 (
            .O(N__74936),
            .I(N__74933));
    LocalMux I__18646 (
            .O(N__74933),
            .I(\PROM.ROMDATA.m349_ns ));
    CascadeMux I__18645 (
            .O(N__74930),
            .I(\PROM.ROMDATA.m331_bm_cascade_ ));
    InMux I__18644 (
            .O(N__74927),
            .I(N__74924));
    LocalMux I__18643 (
            .O(N__74924),
            .I(N__74921));
    Span4Mux_v I__18642 (
            .O(N__74921),
            .I(N__74918));
    Odrv4 I__18641 (
            .O(N__74918),
            .I(\PROM.ROMDATA.m323_bm ));
    CascadeMux I__18640 (
            .O(N__74915),
            .I(\PROM.ROMDATA.m323_am_cascade_ ));
    InMux I__18639 (
            .O(N__74912),
            .I(N__74909));
    LocalMux I__18638 (
            .O(N__74909),
            .I(N__74906));
    Odrv12 I__18637 (
            .O(N__74906),
            .I(\PROM.ROMDATA.m323_ns ));
    CascadeMux I__18636 (
            .O(N__74903),
            .I(N__74899));
    CascadeMux I__18635 (
            .O(N__74902),
            .I(N__74896));
    InMux I__18634 (
            .O(N__74899),
            .I(N__74891));
    InMux I__18633 (
            .O(N__74896),
            .I(N__74883));
    InMux I__18632 (
            .O(N__74895),
            .I(N__74879));
    CascadeMux I__18631 (
            .O(N__74894),
            .I(N__74876));
    LocalMux I__18630 (
            .O(N__74891),
            .I(N__74873));
    InMux I__18629 (
            .O(N__74890),
            .I(N__74870));
    CascadeMux I__18628 (
            .O(N__74889),
            .I(N__74867));
    CascadeMux I__18627 (
            .O(N__74888),
            .I(N__74864));
    CascadeMux I__18626 (
            .O(N__74887),
            .I(N__74861));
    CascadeMux I__18625 (
            .O(N__74886),
            .I(N__74857));
    LocalMux I__18624 (
            .O(N__74883),
            .I(N__74850));
    InMux I__18623 (
            .O(N__74882),
            .I(N__74847));
    LocalMux I__18622 (
            .O(N__74879),
            .I(N__74844));
    InMux I__18621 (
            .O(N__74876),
            .I(N__74841));
    Span4Mux_v I__18620 (
            .O(N__74873),
            .I(N__74838));
    LocalMux I__18619 (
            .O(N__74870),
            .I(N__74835));
    InMux I__18618 (
            .O(N__74867),
            .I(N__74827));
    InMux I__18617 (
            .O(N__74864),
            .I(N__74827));
    InMux I__18616 (
            .O(N__74861),
            .I(N__74817));
    InMux I__18615 (
            .O(N__74860),
            .I(N__74817));
    InMux I__18614 (
            .O(N__74857),
            .I(N__74817));
    InMux I__18613 (
            .O(N__74856),
            .I(N__74812));
    InMux I__18612 (
            .O(N__74855),
            .I(N__74809));
    InMux I__18611 (
            .O(N__74854),
            .I(N__74804));
    InMux I__18610 (
            .O(N__74853),
            .I(N__74804));
    Span4Mux_v I__18609 (
            .O(N__74850),
            .I(N__74801));
    LocalMux I__18608 (
            .O(N__74847),
            .I(N__74798));
    Span4Mux_h I__18607 (
            .O(N__74844),
            .I(N__74793));
    LocalMux I__18606 (
            .O(N__74841),
            .I(N__74793));
    Span4Mux_h I__18605 (
            .O(N__74838),
            .I(N__74788));
    Span4Mux_h I__18604 (
            .O(N__74835),
            .I(N__74788));
    InMux I__18603 (
            .O(N__74834),
            .I(N__74785));
    InMux I__18602 (
            .O(N__74833),
            .I(N__74782));
    CascadeMux I__18601 (
            .O(N__74832),
            .I(N__74779));
    LocalMux I__18600 (
            .O(N__74827),
            .I(N__74775));
    CascadeMux I__18599 (
            .O(N__74826),
            .I(N__74772));
    CascadeMux I__18598 (
            .O(N__74825),
            .I(N__74768));
    CascadeMux I__18597 (
            .O(N__74824),
            .I(N__74765));
    LocalMux I__18596 (
            .O(N__74817),
            .I(N__74762));
    CascadeMux I__18595 (
            .O(N__74816),
            .I(N__74759));
    InMux I__18594 (
            .O(N__74815),
            .I(N__74756));
    LocalMux I__18593 (
            .O(N__74812),
            .I(N__74753));
    LocalMux I__18592 (
            .O(N__74809),
            .I(N__74750));
    LocalMux I__18591 (
            .O(N__74804),
            .I(N__74739));
    Span4Mux_h I__18590 (
            .O(N__74801),
            .I(N__74739));
    Span4Mux_v I__18589 (
            .O(N__74798),
            .I(N__74739));
    Span4Mux_v I__18588 (
            .O(N__74793),
            .I(N__74739));
    Span4Mux_h I__18587 (
            .O(N__74788),
            .I(N__74739));
    LocalMux I__18586 (
            .O(N__74785),
            .I(N__74736));
    LocalMux I__18585 (
            .O(N__74782),
            .I(N__74733));
    InMux I__18584 (
            .O(N__74779),
            .I(N__74730));
    InMux I__18583 (
            .O(N__74778),
            .I(N__74727));
    Span4Mux_v I__18582 (
            .O(N__74775),
            .I(N__74724));
    InMux I__18581 (
            .O(N__74772),
            .I(N__74715));
    InMux I__18580 (
            .O(N__74771),
            .I(N__74715));
    InMux I__18579 (
            .O(N__74768),
            .I(N__74715));
    InMux I__18578 (
            .O(N__74765),
            .I(N__74715));
    Span4Mux_v I__18577 (
            .O(N__74762),
            .I(N__74712));
    InMux I__18576 (
            .O(N__74759),
            .I(N__74709));
    LocalMux I__18575 (
            .O(N__74756),
            .I(N__74706));
    Span4Mux_h I__18574 (
            .O(N__74753),
            .I(N__74703));
    Span4Mux_v I__18573 (
            .O(N__74750),
            .I(N__74700));
    Span4Mux_h I__18572 (
            .O(N__74739),
            .I(N__74697));
    Span4Mux_v I__18571 (
            .O(N__74736),
            .I(N__74694));
    Span4Mux_v I__18570 (
            .O(N__74733),
            .I(N__74691));
    LocalMux I__18569 (
            .O(N__74730),
            .I(N__74686));
    LocalMux I__18568 (
            .O(N__74727),
            .I(N__74686));
    Span4Mux_v I__18567 (
            .O(N__74724),
            .I(N__74683));
    LocalMux I__18566 (
            .O(N__74715),
            .I(N__74674));
    Sp12to4 I__18565 (
            .O(N__74712),
            .I(N__74674));
    LocalMux I__18564 (
            .O(N__74709),
            .I(N__74674));
    Span4Mux_h I__18563 (
            .O(N__74706),
            .I(N__74671));
    Span4Mux_v I__18562 (
            .O(N__74703),
            .I(N__74666));
    Span4Mux_h I__18561 (
            .O(N__74700),
            .I(N__74666));
    Span4Mux_v I__18560 (
            .O(N__74697),
            .I(N__74663));
    Span4Mux_v I__18559 (
            .O(N__74694),
            .I(N__74658));
    Span4Mux_h I__18558 (
            .O(N__74691),
            .I(N__74658));
    Span4Mux_h I__18557 (
            .O(N__74686),
            .I(N__74655));
    Span4Mux_h I__18556 (
            .O(N__74683),
            .I(N__74652));
    InMux I__18555 (
            .O(N__74682),
            .I(N__74649));
    InMux I__18554 (
            .O(N__74681),
            .I(N__74646));
    Span12Mux_h I__18553 (
            .O(N__74674),
            .I(N__74643));
    Span4Mux_h I__18552 (
            .O(N__74671),
            .I(N__74636));
    Span4Mux_h I__18551 (
            .O(N__74666),
            .I(N__74636));
    Span4Mux_v I__18550 (
            .O(N__74663),
            .I(N__74636));
    Span4Mux_h I__18549 (
            .O(N__74658),
            .I(N__74629));
    Span4Mux_v I__18548 (
            .O(N__74655),
            .I(N__74629));
    Span4Mux_h I__18547 (
            .O(N__74652),
            .I(N__74629));
    LocalMux I__18546 (
            .O(N__74649),
            .I(aluParams_1));
    LocalMux I__18545 (
            .O(N__74646),
            .I(aluParams_1));
    Odrv12 I__18544 (
            .O(N__74643),
            .I(aluParams_1));
    Odrv4 I__18543 (
            .O(N__74636),
            .I(aluParams_1));
    Odrv4 I__18542 (
            .O(N__74629),
            .I(aluParams_1));
    InMux I__18541 (
            .O(N__74618),
            .I(N__74615));
    LocalMux I__18540 (
            .O(N__74615),
            .I(N__74612));
    Odrv12 I__18539 (
            .O(N__74612),
            .I(\ALU.un14_log_0_0_15 ));
    InMux I__18538 (
            .O(N__74609),
            .I(N__74604));
    InMux I__18537 (
            .O(N__74608),
            .I(N__74600));
    InMux I__18536 (
            .O(N__74607),
            .I(N__74597));
    LocalMux I__18535 (
            .O(N__74604),
            .I(N__74593));
    InMux I__18534 (
            .O(N__74603),
            .I(N__74590));
    LocalMux I__18533 (
            .O(N__74600),
            .I(N__74587));
    LocalMux I__18532 (
            .O(N__74597),
            .I(N__74584));
    InMux I__18531 (
            .O(N__74596),
            .I(N__74581));
    Span4Mux_h I__18530 (
            .O(N__74593),
            .I(N__74578));
    LocalMux I__18529 (
            .O(N__74590),
            .I(N__74575));
    Span12Mux_v I__18528 (
            .O(N__74587),
            .I(N__74572));
    Span4Mux_v I__18527 (
            .O(N__74584),
            .I(N__74566));
    LocalMux I__18526 (
            .O(N__74581),
            .I(N__74563));
    Span4Mux_h I__18525 (
            .O(N__74578),
            .I(N__74560));
    Span12Mux_s11_h I__18524 (
            .O(N__74575),
            .I(N__74555));
    Span12Mux_h I__18523 (
            .O(N__74572),
            .I(N__74555));
    InMux I__18522 (
            .O(N__74571),
            .I(N__74548));
    InMux I__18521 (
            .O(N__74570),
            .I(N__74548));
    InMux I__18520 (
            .O(N__74569),
            .I(N__74548));
    Span4Mux_v I__18519 (
            .O(N__74566),
            .I(N__74545));
    Span4Mux_h I__18518 (
            .O(N__74563),
            .I(N__74542));
    Span4Mux_h I__18517 (
            .O(N__74560),
            .I(N__74539));
    Odrv12 I__18516 (
            .O(N__74555),
            .I(\ALU.status_19_14 ));
    LocalMux I__18515 (
            .O(N__74548),
            .I(\ALU.status_19_14 ));
    Odrv4 I__18514 (
            .O(N__74545),
            .I(\ALU.status_19_14 ));
    Odrv4 I__18513 (
            .O(N__74542),
            .I(\ALU.status_19_14 ));
    Odrv4 I__18512 (
            .O(N__74539),
            .I(\ALU.status_19_14 ));
    InMux I__18511 (
            .O(N__74528),
            .I(N__74525));
    LocalMux I__18510 (
            .O(N__74525),
            .I(N__74521));
    InMux I__18509 (
            .O(N__74524),
            .I(N__74518));
    Span4Mux_h I__18508 (
            .O(N__74521),
            .I(N__74515));
    LocalMux I__18507 (
            .O(N__74518),
            .I(N__74512));
    Odrv4 I__18506 (
            .O(N__74515),
            .I(\ALU.N_586 ));
    Odrv12 I__18505 (
            .O(N__74512),
            .I(\ALU.N_586 ));
    InMux I__18504 (
            .O(N__74507),
            .I(N__74504));
    LocalMux I__18503 (
            .O(N__74504),
            .I(\PROM.ROMDATA.m331_am ));
    InMux I__18502 (
            .O(N__74501),
            .I(N__74498));
    LocalMux I__18501 (
            .O(N__74498),
            .I(\PROM.ROMDATA.m357_bm ));
    CascadeMux I__18500 (
            .O(N__74495),
            .I(\PROM.ROMDATA.m357_am_cascade_ ));
    InMux I__18499 (
            .O(N__74492),
            .I(N__74484));
    InMux I__18498 (
            .O(N__74491),
            .I(N__74481));
    InMux I__18497 (
            .O(N__74490),
            .I(N__74477));
    InMux I__18496 (
            .O(N__74489),
            .I(N__74474));
    InMux I__18495 (
            .O(N__74488),
            .I(N__74471));
    InMux I__18494 (
            .O(N__74487),
            .I(N__74468));
    LocalMux I__18493 (
            .O(N__74484),
            .I(N__74465));
    LocalMux I__18492 (
            .O(N__74481),
            .I(N__74462));
    InMux I__18491 (
            .O(N__74480),
            .I(N__74459));
    LocalMux I__18490 (
            .O(N__74477),
            .I(N__74454));
    LocalMux I__18489 (
            .O(N__74474),
            .I(N__74454));
    LocalMux I__18488 (
            .O(N__74471),
            .I(N__74451));
    LocalMux I__18487 (
            .O(N__74468),
            .I(N__74448));
    Span4Mux_v I__18486 (
            .O(N__74465),
            .I(N__74444));
    Span4Mux_v I__18485 (
            .O(N__74462),
            .I(N__74439));
    LocalMux I__18484 (
            .O(N__74459),
            .I(N__74439));
    Span4Mux_v I__18483 (
            .O(N__74454),
            .I(N__74434));
    Span4Mux_v I__18482 (
            .O(N__74451),
            .I(N__74434));
    Span4Mux_v I__18481 (
            .O(N__74448),
            .I(N__74431));
    InMux I__18480 (
            .O(N__74447),
            .I(N__74428));
    Span4Mux_v I__18479 (
            .O(N__74444),
            .I(N__74423));
    Span4Mux_h I__18478 (
            .O(N__74439),
            .I(N__74423));
    Span4Mux_h I__18477 (
            .O(N__74434),
            .I(N__74416));
    Span4Mux_h I__18476 (
            .O(N__74431),
            .I(N__74416));
    LocalMux I__18475 (
            .O(N__74428),
            .I(N__74416));
    Odrv4 I__18474 (
            .O(N__74423),
            .I(\PROM.ROMDATA.m178 ));
    Odrv4 I__18473 (
            .O(N__74416),
            .I(\PROM.ROMDATA.m178 ));
    CascadeMux I__18472 (
            .O(N__74411),
            .I(N__74407));
    InMux I__18471 (
            .O(N__74410),
            .I(N__74403));
    InMux I__18470 (
            .O(N__74407),
            .I(N__74400));
    InMux I__18469 (
            .O(N__74406),
            .I(N__74397));
    LocalMux I__18468 (
            .O(N__74403),
            .I(N__74394));
    LocalMux I__18467 (
            .O(N__74400),
            .I(N__74391));
    LocalMux I__18466 (
            .O(N__74397),
            .I(N__74386));
    Span12Mux_h I__18465 (
            .O(N__74394),
            .I(N__74386));
    Span4Mux_v I__18464 (
            .O(N__74391),
            .I(N__74383));
    Odrv12 I__18463 (
            .O(N__74386),
            .I(\PROM.ROMDATA.m287 ));
    Odrv4 I__18462 (
            .O(N__74383),
            .I(\PROM.ROMDATA.m287 ));
    InMux I__18461 (
            .O(N__74378),
            .I(N__74375));
    LocalMux I__18460 (
            .O(N__74375),
            .I(N__74372));
    Span4Mux_h I__18459 (
            .O(N__74372),
            .I(N__74369));
    Span4Mux_h I__18458 (
            .O(N__74369),
            .I(N__74366));
    Odrv4 I__18457 (
            .O(N__74366),
            .I(\PROM.ROMDATA.m294_ns ));
    CascadeMux I__18456 (
            .O(N__74363),
            .I(\PROM.ROMDATA.m290_cascade_ ));
    CascadeMux I__18455 (
            .O(N__74360),
            .I(N__74357));
    InMux I__18454 (
            .O(N__74357),
            .I(N__74354));
    LocalMux I__18453 (
            .O(N__74354),
            .I(N__74351));
    Odrv4 I__18452 (
            .O(N__74351),
            .I(\PROM.ROMDATA.m303_ns_1 ));
    InMux I__18451 (
            .O(N__74348),
            .I(N__74345));
    LocalMux I__18450 (
            .O(N__74345),
            .I(N__74342));
    Odrv4 I__18449 (
            .O(N__74342),
            .I(\PROM.ROMDATA.m361_ns ));
    CascadeMux I__18448 (
            .O(N__74339),
            .I(N__74336));
    InMux I__18447 (
            .O(N__74336),
            .I(N__74333));
    LocalMux I__18446 (
            .O(N__74333),
            .I(\PROM.ROMDATA.m357_ns ));
    InMux I__18445 (
            .O(N__74330),
            .I(N__74324));
    InMux I__18444 (
            .O(N__74329),
            .I(N__74324));
    LocalMux I__18443 (
            .O(N__74324),
            .I(N__74321));
    Sp12to4 I__18442 (
            .O(N__74321),
            .I(N__74318));
    Span12Mux_h I__18441 (
            .O(N__74318),
            .I(N__74315));
    Odrv12 I__18440 (
            .O(N__74315),
            .I(\PROM.ROMDATA.m363_ns ));
    CascadeMux I__18439 (
            .O(N__74312),
            .I(\PROM.ROMDATA.m353_am_cascade_ ));
    InMux I__18438 (
            .O(N__74309),
            .I(N__74306));
    LocalMux I__18437 (
            .O(N__74306),
            .I(N__74303));
    Span4Mux_v I__18436 (
            .O(N__74303),
            .I(N__74300));
    Span4Mux_h I__18435 (
            .O(N__74300),
            .I(N__74297));
    Odrv4 I__18434 (
            .O(N__74297),
            .I(\PROM.ROMDATA.m353_bm ));
    CascadeMux I__18433 (
            .O(N__74294),
            .I(\PROM.ROMDATA.m353_ns_cascade_ ));
    InMux I__18432 (
            .O(N__74291),
            .I(N__74288));
    LocalMux I__18431 (
            .O(N__74288),
            .I(\PROM.ROMDATA.m363_ns_1 ));
    CascadeMux I__18430 (
            .O(N__74285),
            .I(N__74282));
    InMux I__18429 (
            .O(N__74282),
            .I(N__74279));
    LocalMux I__18428 (
            .O(N__74279),
            .I(N__74276));
    Span4Mux_v I__18427 (
            .O(N__74276),
            .I(N__74273));
    Odrv4 I__18426 (
            .O(N__74273),
            .I(\PROM.ROMDATA.m373 ));
    InMux I__18425 (
            .O(N__74270),
            .I(N__74267));
    LocalMux I__18424 (
            .O(N__74267),
            .I(N__74264));
    Span4Mux_v I__18423 (
            .O(N__74264),
            .I(N__74261));
    Odrv4 I__18422 (
            .O(N__74261),
            .I(\PROM.ROMDATA.m298_ns ));
    InMux I__18421 (
            .O(N__74258),
            .I(N__74255));
    LocalMux I__18420 (
            .O(N__74255),
            .I(N__74252));
    Span4Mux_h I__18419 (
            .O(N__74252),
            .I(N__74249));
    Odrv4 I__18418 (
            .O(N__74249),
            .I(\PROM.ROMDATA.m303_ns ));
    InMux I__18417 (
            .O(N__74246),
            .I(N__74243));
    LocalMux I__18416 (
            .O(N__74243),
            .I(N__74240));
    Span4Mux_v I__18415 (
            .O(N__74240),
            .I(N__74236));
    InMux I__18414 (
            .O(N__74239),
            .I(N__74233));
    Span4Mux_h I__18413 (
            .O(N__74236),
            .I(N__74230));
    LocalMux I__18412 (
            .O(N__74233),
            .I(\PROM.ROMDATA.m262 ));
    Odrv4 I__18411 (
            .O(N__74230),
            .I(\PROM.ROMDATA.m262 ));
    InMux I__18410 (
            .O(N__74225),
            .I(N__74222));
    LocalMux I__18409 (
            .O(N__74222),
            .I(N__74219));
    Span4Mux_h I__18408 (
            .O(N__74219),
            .I(N__74216));
    Odrv4 I__18407 (
            .O(N__74216),
            .I(\PROM.ROMDATA.m422_ns ));
    InMux I__18406 (
            .O(N__74213),
            .I(N__74207));
    InMux I__18405 (
            .O(N__74212),
            .I(N__74207));
    LocalMux I__18404 (
            .O(N__74207),
            .I(N__74204));
    Span4Mux_h I__18403 (
            .O(N__74204),
            .I(N__74201));
    Span4Mux_h I__18402 (
            .O(N__74201),
            .I(N__74198));
    Span4Mux_h I__18401 (
            .O(N__74198),
            .I(N__74195));
    Odrv4 I__18400 (
            .O(N__74195),
            .I(\PROM.ROMDATA.m424 ));
    InMux I__18399 (
            .O(N__74192),
            .I(N__74189));
    LocalMux I__18398 (
            .O(N__74189),
            .I(\PROM.ROMDATA.m361_bm ));
    InMux I__18397 (
            .O(N__74186),
            .I(N__74182));
    InMux I__18396 (
            .O(N__74185),
            .I(N__74179));
    LocalMux I__18395 (
            .O(N__74182),
            .I(N__74176));
    LocalMux I__18394 (
            .O(N__74179),
            .I(\PROM.ROMDATA.m127 ));
    Odrv12 I__18393 (
            .O(N__74176),
            .I(\PROM.ROMDATA.m127 ));
    InMux I__18392 (
            .O(N__74171),
            .I(N__74168));
    LocalMux I__18391 (
            .O(N__74168),
            .I(\PROM.ROMDATA.m128 ));
    CascadeMux I__18390 (
            .O(N__74165),
            .I(\PROM.ROMDATA.m137_am_cascade_ ));
    InMux I__18389 (
            .O(N__74162),
            .I(N__74159));
    LocalMux I__18388 (
            .O(N__74159),
            .I(\PROM.ROMDATA.m137_bm ));
    InMux I__18387 (
            .O(N__74156),
            .I(N__74153));
    LocalMux I__18386 (
            .O(N__74153),
            .I(\PROM.ROMDATA.m147_am ));
    InMux I__18385 (
            .O(N__74150),
            .I(N__74147));
    LocalMux I__18384 (
            .O(N__74147),
            .I(N__74144));
    Odrv4 I__18383 (
            .O(N__74144),
            .I(\PROM.ROMDATA.m147_bm ));
    CascadeMux I__18382 (
            .O(N__74141),
            .I(\PROM.ROMDATA.m148_ns_1_cascade_ ));
    InMux I__18381 (
            .O(N__74138),
            .I(N__74135));
    LocalMux I__18380 (
            .O(N__74135),
            .I(N__74132));
    Odrv12 I__18379 (
            .O(N__74132),
            .I(\PROM.ROMDATA.m148_ns ));
    InMux I__18378 (
            .O(N__74129),
            .I(N__74126));
    LocalMux I__18377 (
            .O(N__74126),
            .I(N__74122));
    InMux I__18376 (
            .O(N__74125),
            .I(N__74119));
    Span4Mux_v I__18375 (
            .O(N__74122),
            .I(N__74116));
    LocalMux I__18374 (
            .O(N__74119),
            .I(N__74111));
    Span4Mux_h I__18373 (
            .O(N__74116),
            .I(N__74111));
    Odrv4 I__18372 (
            .O(N__74111),
            .I(\PROM.ROMDATA.m292 ));
    CascadeMux I__18371 (
            .O(N__74108),
            .I(N__74105));
    InMux I__18370 (
            .O(N__74105),
            .I(N__74102));
    LocalMux I__18369 (
            .O(N__74102),
            .I(N__74099));
    Span12Mux_v I__18368 (
            .O(N__74099),
            .I(N__74096));
    Odrv12 I__18367 (
            .O(N__74096),
            .I(\PROM.ROMDATA.m299 ));
    InMux I__18366 (
            .O(N__74093),
            .I(N__74090));
    LocalMux I__18365 (
            .O(N__74090),
            .I(\PROM.ROMDATA.m301 ));
    InMux I__18364 (
            .O(N__74087),
            .I(N__74084));
    LocalMux I__18363 (
            .O(N__74084),
            .I(N__74081));
    Span4Mux_v I__18362 (
            .O(N__74081),
            .I(N__74078));
    Span4Mux_h I__18361 (
            .O(N__74078),
            .I(N__74075));
    Odrv4 I__18360 (
            .O(N__74075),
            .I(\PROM.ROMDATA.m488_ns_1 ));
    InMux I__18359 (
            .O(N__74072),
            .I(N__74062));
    InMux I__18358 (
            .O(N__74071),
            .I(N__74058));
    InMux I__18357 (
            .O(N__74070),
            .I(N__74053));
    InMux I__18356 (
            .O(N__74069),
            .I(N__74053));
    InMux I__18355 (
            .O(N__74068),
            .I(N__74050));
    InMux I__18354 (
            .O(N__74067),
            .I(N__74045));
    InMux I__18353 (
            .O(N__74066),
            .I(N__74045));
    InMux I__18352 (
            .O(N__74065),
            .I(N__74042));
    LocalMux I__18351 (
            .O(N__74062),
            .I(N__74039));
    InMux I__18350 (
            .O(N__74061),
            .I(N__74034));
    LocalMux I__18349 (
            .O(N__74058),
            .I(N__74031));
    LocalMux I__18348 (
            .O(N__74053),
            .I(N__74024));
    LocalMux I__18347 (
            .O(N__74050),
            .I(N__74024));
    LocalMux I__18346 (
            .O(N__74045),
            .I(N__74024));
    LocalMux I__18345 (
            .O(N__74042),
            .I(N__74020));
    Span4Mux_v I__18344 (
            .O(N__74039),
            .I(N__74017));
    InMux I__18343 (
            .O(N__74038),
            .I(N__74012));
    InMux I__18342 (
            .O(N__74037),
            .I(N__74012));
    LocalMux I__18341 (
            .O(N__74034),
            .I(N__74008));
    Span4Mux_v I__18340 (
            .O(N__74031),
            .I(N__74004));
    Span4Mux_v I__18339 (
            .O(N__74024),
            .I(N__74001));
    InMux I__18338 (
            .O(N__74023),
            .I(N__73998));
    Span4Mux_v I__18337 (
            .O(N__74020),
            .I(N__73994));
    Span4Mux_h I__18336 (
            .O(N__74017),
            .I(N__73989));
    LocalMux I__18335 (
            .O(N__74012),
            .I(N__73989));
    InMux I__18334 (
            .O(N__74011),
            .I(N__73986));
    Span4Mux_v I__18333 (
            .O(N__74008),
            .I(N__73983));
    InMux I__18332 (
            .O(N__74007),
            .I(N__73980));
    Span4Mux_h I__18331 (
            .O(N__74004),
            .I(N__73977));
    Span4Mux_h I__18330 (
            .O(N__74001),
            .I(N__73972));
    LocalMux I__18329 (
            .O(N__73998),
            .I(N__73972));
    InMux I__18328 (
            .O(N__73997),
            .I(N__73969));
    Span4Mux_h I__18327 (
            .O(N__73994),
            .I(N__73964));
    Span4Mux_h I__18326 (
            .O(N__73989),
            .I(N__73964));
    LocalMux I__18325 (
            .O(N__73986),
            .I(N__73959));
    Span4Mux_h I__18324 (
            .O(N__73983),
            .I(N__73959));
    LocalMux I__18323 (
            .O(N__73980),
            .I(m125_e));
    Odrv4 I__18322 (
            .O(N__73977),
            .I(m125_e));
    Odrv4 I__18321 (
            .O(N__73972),
            .I(m125_e));
    LocalMux I__18320 (
            .O(N__73969),
            .I(m125_e));
    Odrv4 I__18319 (
            .O(N__73964),
            .I(m125_e));
    Odrv4 I__18318 (
            .O(N__73959),
            .I(m125_e));
    CascadeMux I__18317 (
            .O(N__73946),
            .I(N__73942));
    InMux I__18316 (
            .O(N__73945),
            .I(N__73937));
    InMux I__18315 (
            .O(N__73942),
            .I(N__73937));
    LocalMux I__18314 (
            .O(N__73937),
            .I(N__73934));
    Span4Mux_v I__18313 (
            .O(N__73934),
            .I(N__73931));
    Span4Mux_h I__18312 (
            .O(N__73931),
            .I(N__73928));
    Span4Mux_h I__18311 (
            .O(N__73928),
            .I(N__73925));
    Span4Mux_h I__18310 (
            .O(N__73925),
            .I(N__73922));
    Odrv4 I__18309 (
            .O(N__73922),
            .I(\PROM.ROMDATA.N_570_mux ));
    CascadeMux I__18308 (
            .O(N__73919),
            .I(N__73915));
    CascadeMux I__18307 (
            .O(N__73918),
            .I(N__73912));
    InMux I__18306 (
            .O(N__73915),
            .I(N__73906));
    InMux I__18305 (
            .O(N__73912),
            .I(N__73906));
    CascadeMux I__18304 (
            .O(N__73911),
            .I(N__73902));
    LocalMux I__18303 (
            .O(N__73906),
            .I(N__73899));
    InMux I__18302 (
            .O(N__73905),
            .I(N__73896));
    InMux I__18301 (
            .O(N__73902),
            .I(N__73893));
    Span4Mux_v I__18300 (
            .O(N__73899),
            .I(N__73886));
    LocalMux I__18299 (
            .O(N__73896),
            .I(N__73886));
    LocalMux I__18298 (
            .O(N__73893),
            .I(N__73883));
    CascadeMux I__18297 (
            .O(N__73892),
            .I(N__73880));
    CascadeMux I__18296 (
            .O(N__73891),
            .I(N__73877));
    Span4Mux_v I__18295 (
            .O(N__73886),
            .I(N__73874));
    Span4Mux_h I__18294 (
            .O(N__73883),
            .I(N__73870));
    InMux I__18293 (
            .O(N__73880),
            .I(N__73867));
    InMux I__18292 (
            .O(N__73877),
            .I(N__73864));
    Span4Mux_h I__18291 (
            .O(N__73874),
            .I(N__73861));
    CascadeMux I__18290 (
            .O(N__73873),
            .I(N__73858));
    Span4Mux_v I__18289 (
            .O(N__73870),
            .I(N__73852));
    LocalMux I__18288 (
            .O(N__73867),
            .I(N__73852));
    LocalMux I__18287 (
            .O(N__73864),
            .I(N__73849));
    Span4Mux_h I__18286 (
            .O(N__73861),
            .I(N__73846));
    InMux I__18285 (
            .O(N__73858),
            .I(N__73841));
    InMux I__18284 (
            .O(N__73857),
            .I(N__73841));
    Span4Mux_h I__18283 (
            .O(N__73852),
            .I(N__73838));
    Odrv12 I__18282 (
            .O(N__73849),
            .I(\PROM.ROMDATA.m2 ));
    Odrv4 I__18281 (
            .O(N__73846),
            .I(\PROM.ROMDATA.m2 ));
    LocalMux I__18280 (
            .O(N__73841),
            .I(\PROM.ROMDATA.m2 ));
    Odrv4 I__18279 (
            .O(N__73838),
            .I(\PROM.ROMDATA.m2 ));
    InMux I__18278 (
            .O(N__73829),
            .I(N__73826));
    LocalMux I__18277 (
            .O(N__73826),
            .I(N__73823));
    Odrv4 I__18276 (
            .O(N__73823),
            .I(\PROM.ROMDATA.m493_am ));
    InMux I__18275 (
            .O(N__73820),
            .I(N__73817));
    LocalMux I__18274 (
            .O(N__73817),
            .I(N__73814));
    Span4Mux_v I__18273 (
            .O(N__73814),
            .I(N__73805));
    InMux I__18272 (
            .O(N__73813),
            .I(N__73800));
    InMux I__18271 (
            .O(N__73812),
            .I(N__73800));
    InMux I__18270 (
            .O(N__73811),
            .I(N__73797));
    InMux I__18269 (
            .O(N__73810),
            .I(N__73794));
    InMux I__18268 (
            .O(N__73809),
            .I(N__73791));
    InMux I__18267 (
            .O(N__73808),
            .I(N__73788));
    Span4Mux_h I__18266 (
            .O(N__73805),
            .I(N__73784));
    LocalMux I__18265 (
            .O(N__73800),
            .I(N__73781));
    LocalMux I__18264 (
            .O(N__73797),
            .I(N__73778));
    LocalMux I__18263 (
            .O(N__73794),
            .I(N__73773));
    LocalMux I__18262 (
            .O(N__73791),
            .I(N__73773));
    LocalMux I__18261 (
            .O(N__73788),
            .I(N__73770));
    InMux I__18260 (
            .O(N__73787),
            .I(N__73767));
    Span4Mux_h I__18259 (
            .O(N__73784),
            .I(N__73761));
    Span4Mux_v I__18258 (
            .O(N__73781),
            .I(N__73761));
    Span4Mux_v I__18257 (
            .O(N__73778),
            .I(N__73752));
    Span4Mux_v I__18256 (
            .O(N__73773),
            .I(N__73752));
    Span4Mux_v I__18255 (
            .O(N__73770),
            .I(N__73752));
    LocalMux I__18254 (
            .O(N__73767),
            .I(N__73752));
    InMux I__18253 (
            .O(N__73766),
            .I(N__73749));
    Odrv4 I__18252 (
            .O(N__73761),
            .I(CONTROL_addrstack_reto_1));
    Odrv4 I__18251 (
            .O(N__73752),
            .I(CONTROL_addrstack_reto_1));
    LocalMux I__18250 (
            .O(N__73749),
            .I(CONTROL_addrstack_reto_1));
    CascadeMux I__18249 (
            .O(N__73742),
            .I(N__73737));
    CascadeMux I__18248 (
            .O(N__73741),
            .I(N__73734));
    CascadeMux I__18247 (
            .O(N__73740),
            .I(N__73731));
    InMux I__18246 (
            .O(N__73737),
            .I(N__73725));
    InMux I__18245 (
            .O(N__73734),
            .I(N__73722));
    InMux I__18244 (
            .O(N__73731),
            .I(N__73716));
    CascadeMux I__18243 (
            .O(N__73730),
            .I(N__73713));
    InMux I__18242 (
            .O(N__73729),
            .I(N__73707));
    InMux I__18241 (
            .O(N__73728),
            .I(N__73707));
    LocalMux I__18240 (
            .O(N__73725),
            .I(N__73702));
    LocalMux I__18239 (
            .O(N__73722),
            .I(N__73702));
    InMux I__18238 (
            .O(N__73721),
            .I(N__73697));
    InMux I__18237 (
            .O(N__73720),
            .I(N__73697));
    CascadeMux I__18236 (
            .O(N__73719),
            .I(N__73694));
    LocalMux I__18235 (
            .O(N__73716),
            .I(N__73691));
    InMux I__18234 (
            .O(N__73713),
            .I(N__73688));
    InMux I__18233 (
            .O(N__73712),
            .I(N__73683));
    LocalMux I__18232 (
            .O(N__73707),
            .I(N__73680));
    Span4Mux_v I__18231 (
            .O(N__73702),
            .I(N__73672));
    LocalMux I__18230 (
            .O(N__73697),
            .I(N__73672));
    InMux I__18229 (
            .O(N__73694),
            .I(N__73669));
    Span4Mux_v I__18228 (
            .O(N__73691),
            .I(N__73665));
    LocalMux I__18227 (
            .O(N__73688),
            .I(N__73662));
    InMux I__18226 (
            .O(N__73687),
            .I(N__73658));
    InMux I__18225 (
            .O(N__73686),
            .I(N__73655));
    LocalMux I__18224 (
            .O(N__73683),
            .I(N__73652));
    Span4Mux_v I__18223 (
            .O(N__73680),
            .I(N__73649));
    InMux I__18222 (
            .O(N__73679),
            .I(N__73642));
    InMux I__18221 (
            .O(N__73678),
            .I(N__73642));
    InMux I__18220 (
            .O(N__73677),
            .I(N__73642));
    Span4Mux_h I__18219 (
            .O(N__73672),
            .I(N__73637));
    LocalMux I__18218 (
            .O(N__73669),
            .I(N__73637));
    InMux I__18217 (
            .O(N__73668),
            .I(N__73633));
    Span4Mux_h I__18216 (
            .O(N__73665),
            .I(N__73628));
    Span4Mux_v I__18215 (
            .O(N__73662),
            .I(N__73628));
    CascadeMux I__18214 (
            .O(N__73661),
            .I(N__73624));
    LocalMux I__18213 (
            .O(N__73658),
            .I(N__73619));
    LocalMux I__18212 (
            .O(N__73655),
            .I(N__73619));
    Span4Mux_v I__18211 (
            .O(N__73652),
            .I(N__73614));
    Span4Mux_h I__18210 (
            .O(N__73649),
            .I(N__73614));
    LocalMux I__18209 (
            .O(N__73642),
            .I(N__73611));
    Span4Mux_v I__18208 (
            .O(N__73637),
            .I(N__73608));
    InMux I__18207 (
            .O(N__73636),
            .I(N__73605));
    LocalMux I__18206 (
            .O(N__73633),
            .I(N__73600));
    Sp12to4 I__18205 (
            .O(N__73628),
            .I(N__73600));
    InMux I__18204 (
            .O(N__73627),
            .I(N__73595));
    InMux I__18203 (
            .O(N__73624),
            .I(N__73595));
    Span4Mux_v I__18202 (
            .O(N__73619),
            .I(N__73588));
    Span4Mux_h I__18201 (
            .O(N__73614),
            .I(N__73588));
    Span4Mux_v I__18200 (
            .O(N__73611),
            .I(N__73588));
    Span4Mux_h I__18199 (
            .O(N__73608),
            .I(N__73585));
    LocalMux I__18198 (
            .O(N__73605),
            .I(CONTROL_programCounter11_reto));
    Odrv12 I__18197 (
            .O(N__73600),
            .I(CONTROL_programCounter11_reto));
    LocalMux I__18196 (
            .O(N__73595),
            .I(CONTROL_programCounter11_reto));
    Odrv4 I__18195 (
            .O(N__73588),
            .I(CONTROL_programCounter11_reto));
    Odrv4 I__18194 (
            .O(N__73585),
            .I(CONTROL_programCounter11_reto));
    InMux I__18193 (
            .O(N__73574),
            .I(N__73569));
    CascadeMux I__18192 (
            .O(N__73573),
            .I(N__73566));
    InMux I__18191 (
            .O(N__73572),
            .I(N__73562));
    LocalMux I__18190 (
            .O(N__73569),
            .I(N__73559));
    InMux I__18189 (
            .O(N__73566),
            .I(N__73554));
    InMux I__18188 (
            .O(N__73565),
            .I(N__73554));
    LocalMux I__18187 (
            .O(N__73562),
            .I(N__73549));
    Span4Mux_v I__18186 (
            .O(N__73559),
            .I(N__73546));
    LocalMux I__18185 (
            .O(N__73554),
            .I(N__73543));
    InMux I__18184 (
            .O(N__73553),
            .I(N__73539));
    InMux I__18183 (
            .O(N__73552),
            .I(N__73536));
    Span4Mux_v I__18182 (
            .O(N__73549),
            .I(N__73533));
    Sp12to4 I__18181 (
            .O(N__73546),
            .I(N__73530));
    Span4Mux_h I__18180 (
            .O(N__73543),
            .I(N__73527));
    InMux I__18179 (
            .O(N__73542),
            .I(N__73524));
    LocalMux I__18178 (
            .O(N__73539),
            .I(N__73519));
    LocalMux I__18177 (
            .O(N__73536),
            .I(N__73519));
    Span4Mux_h I__18176 (
            .O(N__73533),
            .I(N__73516));
    Odrv12 I__18175 (
            .O(N__73530),
            .I(N_416));
    Odrv4 I__18174 (
            .O(N__73527),
            .I(N_416));
    LocalMux I__18173 (
            .O(N__73524),
            .I(N_416));
    Odrv4 I__18172 (
            .O(N__73519),
            .I(N_416));
    Odrv4 I__18171 (
            .O(N__73516),
            .I(N_416));
    InMux I__18170 (
            .O(N__73505),
            .I(N__73498));
    InMux I__18169 (
            .O(N__73504),
            .I(N__73498));
    InMux I__18168 (
            .O(N__73503),
            .I(N__73495));
    LocalMux I__18167 (
            .O(N__73498),
            .I(N__73492));
    LocalMux I__18166 (
            .O(N__73495),
            .I(N__73488));
    Span4Mux_h I__18165 (
            .O(N__73492),
            .I(N__73485));
    InMux I__18164 (
            .O(N__73491),
            .I(N__73482));
    Span4Mux_h I__18163 (
            .O(N__73488),
            .I(N__73475));
    Span4Mux_h I__18162 (
            .O(N__73485),
            .I(N__73475));
    LocalMux I__18161 (
            .O(N__73482),
            .I(N__73475));
    Span4Mux_v I__18160 (
            .O(N__73475),
            .I(N__73472));
    Odrv4 I__18159 (
            .O(N__73472),
            .I(\PROM.ROMDATA.m1 ));
    CascadeMux I__18158 (
            .O(N__73469),
            .I(N__73466));
    InMux I__18157 (
            .O(N__73466),
            .I(N__73463));
    LocalMux I__18156 (
            .O(N__73463),
            .I(N__73460));
    Span4Mux_h I__18155 (
            .O(N__73460),
            .I(N__73457));
    Odrv4 I__18154 (
            .O(N__73457),
            .I(\PROM.ROMDATA.m493_bm ));
    InMux I__18153 (
            .O(N__73454),
            .I(N__73451));
    LocalMux I__18152 (
            .O(N__73451),
            .I(\PROM.ROMDATA.m361_am ));
    CascadeMux I__18151 (
            .O(N__73448),
            .I(N__73445));
    InMux I__18150 (
            .O(N__73445),
            .I(N__73442));
    LocalMux I__18149 (
            .O(N__73442),
            .I(N__73439));
    Odrv4 I__18148 (
            .O(N__73439),
            .I(\PROM.ROMDATA.m211_ns_N_2L1 ));
    CascadeMux I__18147 (
            .O(N__73436),
            .I(\PROM.ROMDATA.m211_ns_cascade_ ));
    InMux I__18146 (
            .O(N__73433),
            .I(N__73430));
    LocalMux I__18145 (
            .O(N__73430),
            .I(N__73427));
    Span4Mux_h I__18144 (
            .O(N__73427),
            .I(N__73424));
    Span4Mux_h I__18143 (
            .O(N__73424),
            .I(N__73421));
    Odrv4 I__18142 (
            .O(N__73421),
            .I(\PROM.ROMDATA.m221cf0_1 ));
    InMux I__18141 (
            .O(N__73418),
            .I(N__73415));
    LocalMux I__18140 (
            .O(N__73415),
            .I(\PROM.ROMDATA.m211_ns ));
    CascadeMux I__18139 (
            .O(N__73412),
            .I(N__73409));
    InMux I__18138 (
            .O(N__73409),
            .I(N__73406));
    LocalMux I__18137 (
            .O(N__73406),
            .I(N__73403));
    Span4Mux_v I__18136 (
            .O(N__73403),
            .I(N__73400));
    Sp12to4 I__18135 (
            .O(N__73400),
            .I(N__73397));
    Odrv12 I__18134 (
            .O(N__73397),
            .I(\PROM.ROMDATA.m221cf1_1 ));
    CascadeMux I__18133 (
            .O(N__73394),
            .I(N__73391));
    InMux I__18132 (
            .O(N__73391),
            .I(N__73388));
    LocalMux I__18131 (
            .O(N__73388),
            .I(N__73385));
    Span4Mux_v I__18130 (
            .O(N__73385),
            .I(N__73382));
    Span4Mux_h I__18129 (
            .O(N__73382),
            .I(N__73379));
    Sp12to4 I__18128 (
            .O(N__73379),
            .I(N__73376));
    Odrv12 I__18127 (
            .O(N__73376),
            .I(\PROM.ROMDATA.m369 ));
    CascadeMux I__18126 (
            .O(N__73373),
            .I(N__73370));
    InMux I__18125 (
            .O(N__73370),
            .I(N__73367));
    LocalMux I__18124 (
            .O(N__73367),
            .I(N__73364));
    Span4Mux_h I__18123 (
            .O(N__73364),
            .I(N__73361));
    Span4Mux_v I__18122 (
            .O(N__73361),
            .I(N__73358));
    Odrv4 I__18121 (
            .O(N__73358),
            .I(\PROM.ROMDATA.m60 ));
    InMux I__18120 (
            .O(N__73355),
            .I(N__73352));
    LocalMux I__18119 (
            .O(N__73352),
            .I(N__73349));
    Span4Mux_v I__18118 (
            .O(N__73349),
            .I(N__73345));
    InMux I__18117 (
            .O(N__73348),
            .I(N__73342));
    Span4Mux_h I__18116 (
            .O(N__73345),
            .I(N__73339));
    LocalMux I__18115 (
            .O(N__73342),
            .I(N__73336));
    Span4Mux_h I__18114 (
            .O(N__73339),
            .I(N__73333));
    Span4Mux_v I__18113 (
            .O(N__73336),
            .I(N__73330));
    Span4Mux_h I__18112 (
            .O(N__73333),
            .I(N__73327));
    Span4Mux_h I__18111 (
            .O(N__73330),
            .I(N__73324));
    Odrv4 I__18110 (
            .O(N__73327),
            .I(\CONTROL.programCounter_1_7 ));
    Odrv4 I__18109 (
            .O(N__73324),
            .I(\CONTROL.programCounter_1_7 ));
    InMux I__18108 (
            .O(N__73319),
            .I(N__73316));
    LocalMux I__18107 (
            .O(N__73316),
            .I(N__73313));
    Span4Mux_h I__18106 (
            .O(N__73313),
            .I(N__73310));
    Span4Mux_h I__18105 (
            .O(N__73310),
            .I(N__73307));
    Odrv4 I__18104 (
            .O(N__73307),
            .I(\CONTROL.programCounter_1_reto_7 ));
    InMux I__18103 (
            .O(N__73304),
            .I(N__73299));
    InMux I__18102 (
            .O(N__73303),
            .I(N__73294));
    InMux I__18101 (
            .O(N__73302),
            .I(N__73294));
    LocalMux I__18100 (
            .O(N__73299),
            .I(N__73287));
    LocalMux I__18099 (
            .O(N__73294),
            .I(N__73283));
    ClkMux I__18098 (
            .O(N__73293),
            .I(N__72833));
    ClkMux I__18097 (
            .O(N__73292),
            .I(N__72833));
    ClkMux I__18096 (
            .O(N__73291),
            .I(N__72833));
    ClkMux I__18095 (
            .O(N__73290),
            .I(N__72833));
    Glb2LocalMux I__18094 (
            .O(N__73287),
            .I(N__72833));
    ClkMux I__18093 (
            .O(N__73286),
            .I(N__72833));
    Glb2LocalMux I__18092 (
            .O(N__73283),
            .I(N__72833));
    ClkMux I__18091 (
            .O(N__73282),
            .I(N__72833));
    ClkMux I__18090 (
            .O(N__73281),
            .I(N__72833));
    ClkMux I__18089 (
            .O(N__73280),
            .I(N__72833));
    ClkMux I__18088 (
            .O(N__73279),
            .I(N__72833));
    ClkMux I__18087 (
            .O(N__73278),
            .I(N__72833));
    ClkMux I__18086 (
            .O(N__73277),
            .I(N__72833));
    ClkMux I__18085 (
            .O(N__73276),
            .I(N__72833));
    ClkMux I__18084 (
            .O(N__73275),
            .I(N__72833));
    ClkMux I__18083 (
            .O(N__73274),
            .I(N__72833));
    ClkMux I__18082 (
            .O(N__73273),
            .I(N__72833));
    ClkMux I__18081 (
            .O(N__73272),
            .I(N__72833));
    ClkMux I__18080 (
            .O(N__73271),
            .I(N__72833));
    ClkMux I__18079 (
            .O(N__73270),
            .I(N__72833));
    ClkMux I__18078 (
            .O(N__73269),
            .I(N__72833));
    ClkMux I__18077 (
            .O(N__73268),
            .I(N__72833));
    ClkMux I__18076 (
            .O(N__73267),
            .I(N__72833));
    ClkMux I__18075 (
            .O(N__73266),
            .I(N__72833));
    ClkMux I__18074 (
            .O(N__73265),
            .I(N__72833));
    ClkMux I__18073 (
            .O(N__73264),
            .I(N__72833));
    ClkMux I__18072 (
            .O(N__73263),
            .I(N__72833));
    ClkMux I__18071 (
            .O(N__73262),
            .I(N__72833));
    ClkMux I__18070 (
            .O(N__73261),
            .I(N__72833));
    ClkMux I__18069 (
            .O(N__73260),
            .I(N__72833));
    ClkMux I__18068 (
            .O(N__73259),
            .I(N__72833));
    ClkMux I__18067 (
            .O(N__73258),
            .I(N__72833));
    ClkMux I__18066 (
            .O(N__73257),
            .I(N__72833));
    ClkMux I__18065 (
            .O(N__73256),
            .I(N__72833));
    ClkMux I__18064 (
            .O(N__73255),
            .I(N__72833));
    ClkMux I__18063 (
            .O(N__73254),
            .I(N__72833));
    ClkMux I__18062 (
            .O(N__73253),
            .I(N__72833));
    ClkMux I__18061 (
            .O(N__73252),
            .I(N__72833));
    ClkMux I__18060 (
            .O(N__73251),
            .I(N__72833));
    ClkMux I__18059 (
            .O(N__73250),
            .I(N__72833));
    ClkMux I__18058 (
            .O(N__73249),
            .I(N__72833));
    ClkMux I__18057 (
            .O(N__73248),
            .I(N__72833));
    ClkMux I__18056 (
            .O(N__73247),
            .I(N__72833));
    ClkMux I__18055 (
            .O(N__73246),
            .I(N__72833));
    ClkMux I__18054 (
            .O(N__73245),
            .I(N__72833));
    ClkMux I__18053 (
            .O(N__73244),
            .I(N__72833));
    ClkMux I__18052 (
            .O(N__73243),
            .I(N__72833));
    ClkMux I__18051 (
            .O(N__73242),
            .I(N__72833));
    ClkMux I__18050 (
            .O(N__73241),
            .I(N__72833));
    ClkMux I__18049 (
            .O(N__73240),
            .I(N__72833));
    ClkMux I__18048 (
            .O(N__73239),
            .I(N__72833));
    ClkMux I__18047 (
            .O(N__73238),
            .I(N__72833));
    ClkMux I__18046 (
            .O(N__73237),
            .I(N__72833));
    ClkMux I__18045 (
            .O(N__73236),
            .I(N__72833));
    ClkMux I__18044 (
            .O(N__73235),
            .I(N__72833));
    ClkMux I__18043 (
            .O(N__73234),
            .I(N__72833));
    ClkMux I__18042 (
            .O(N__73233),
            .I(N__72833));
    ClkMux I__18041 (
            .O(N__73232),
            .I(N__72833));
    ClkMux I__18040 (
            .O(N__73231),
            .I(N__72833));
    ClkMux I__18039 (
            .O(N__73230),
            .I(N__72833));
    ClkMux I__18038 (
            .O(N__73229),
            .I(N__72833));
    ClkMux I__18037 (
            .O(N__73228),
            .I(N__72833));
    ClkMux I__18036 (
            .O(N__73227),
            .I(N__72833));
    ClkMux I__18035 (
            .O(N__73226),
            .I(N__72833));
    ClkMux I__18034 (
            .O(N__73225),
            .I(N__72833));
    ClkMux I__18033 (
            .O(N__73224),
            .I(N__72833));
    ClkMux I__18032 (
            .O(N__73223),
            .I(N__72833));
    ClkMux I__18031 (
            .O(N__73222),
            .I(N__72833));
    ClkMux I__18030 (
            .O(N__73221),
            .I(N__72833));
    ClkMux I__18029 (
            .O(N__73220),
            .I(N__72833));
    ClkMux I__18028 (
            .O(N__73219),
            .I(N__72833));
    ClkMux I__18027 (
            .O(N__73218),
            .I(N__72833));
    ClkMux I__18026 (
            .O(N__73217),
            .I(N__72833));
    ClkMux I__18025 (
            .O(N__73216),
            .I(N__72833));
    ClkMux I__18024 (
            .O(N__73215),
            .I(N__72833));
    ClkMux I__18023 (
            .O(N__73214),
            .I(N__72833));
    ClkMux I__18022 (
            .O(N__73213),
            .I(N__72833));
    ClkMux I__18021 (
            .O(N__73212),
            .I(N__72833));
    ClkMux I__18020 (
            .O(N__73211),
            .I(N__72833));
    ClkMux I__18019 (
            .O(N__73210),
            .I(N__72833));
    ClkMux I__18018 (
            .O(N__73209),
            .I(N__72833));
    ClkMux I__18017 (
            .O(N__73208),
            .I(N__72833));
    ClkMux I__18016 (
            .O(N__73207),
            .I(N__72833));
    ClkMux I__18015 (
            .O(N__73206),
            .I(N__72833));
    ClkMux I__18014 (
            .O(N__73205),
            .I(N__72833));
    ClkMux I__18013 (
            .O(N__73204),
            .I(N__72833));
    ClkMux I__18012 (
            .O(N__73203),
            .I(N__72833));
    ClkMux I__18011 (
            .O(N__73202),
            .I(N__72833));
    ClkMux I__18010 (
            .O(N__73201),
            .I(N__72833));
    ClkMux I__18009 (
            .O(N__73200),
            .I(N__72833));
    ClkMux I__18008 (
            .O(N__73199),
            .I(N__72833));
    ClkMux I__18007 (
            .O(N__73198),
            .I(N__72833));
    ClkMux I__18006 (
            .O(N__73197),
            .I(N__72833));
    ClkMux I__18005 (
            .O(N__73196),
            .I(N__72833));
    ClkMux I__18004 (
            .O(N__73195),
            .I(N__72833));
    ClkMux I__18003 (
            .O(N__73194),
            .I(N__72833));
    ClkMux I__18002 (
            .O(N__73193),
            .I(N__72833));
    ClkMux I__18001 (
            .O(N__73192),
            .I(N__72833));
    ClkMux I__18000 (
            .O(N__73191),
            .I(N__72833));
    ClkMux I__17999 (
            .O(N__73190),
            .I(N__72833));
    ClkMux I__17998 (
            .O(N__73189),
            .I(N__72833));
    ClkMux I__17997 (
            .O(N__73188),
            .I(N__72833));
    ClkMux I__17996 (
            .O(N__73187),
            .I(N__72833));
    ClkMux I__17995 (
            .O(N__73186),
            .I(N__72833));
    ClkMux I__17994 (
            .O(N__73185),
            .I(N__72833));
    ClkMux I__17993 (
            .O(N__73184),
            .I(N__72833));
    ClkMux I__17992 (
            .O(N__73183),
            .I(N__72833));
    ClkMux I__17991 (
            .O(N__73182),
            .I(N__72833));
    ClkMux I__17990 (
            .O(N__73181),
            .I(N__72833));
    ClkMux I__17989 (
            .O(N__73180),
            .I(N__72833));
    ClkMux I__17988 (
            .O(N__73179),
            .I(N__72833));
    ClkMux I__17987 (
            .O(N__73178),
            .I(N__72833));
    ClkMux I__17986 (
            .O(N__73177),
            .I(N__72833));
    ClkMux I__17985 (
            .O(N__73176),
            .I(N__72833));
    ClkMux I__17984 (
            .O(N__73175),
            .I(N__72833));
    ClkMux I__17983 (
            .O(N__73174),
            .I(N__72833));
    ClkMux I__17982 (
            .O(N__73173),
            .I(N__72833));
    ClkMux I__17981 (
            .O(N__73172),
            .I(N__72833));
    ClkMux I__17980 (
            .O(N__73171),
            .I(N__72833));
    ClkMux I__17979 (
            .O(N__73170),
            .I(N__72833));
    ClkMux I__17978 (
            .O(N__73169),
            .I(N__72833));
    ClkMux I__17977 (
            .O(N__73168),
            .I(N__72833));
    ClkMux I__17976 (
            .O(N__73167),
            .I(N__72833));
    ClkMux I__17975 (
            .O(N__73166),
            .I(N__72833));
    ClkMux I__17974 (
            .O(N__73165),
            .I(N__72833));
    ClkMux I__17973 (
            .O(N__73164),
            .I(N__72833));
    ClkMux I__17972 (
            .O(N__73163),
            .I(N__72833));
    ClkMux I__17971 (
            .O(N__73162),
            .I(N__72833));
    ClkMux I__17970 (
            .O(N__73161),
            .I(N__72833));
    ClkMux I__17969 (
            .O(N__73160),
            .I(N__72833));
    ClkMux I__17968 (
            .O(N__73159),
            .I(N__72833));
    ClkMux I__17967 (
            .O(N__73158),
            .I(N__72833));
    ClkMux I__17966 (
            .O(N__73157),
            .I(N__72833));
    ClkMux I__17965 (
            .O(N__73156),
            .I(N__72833));
    ClkMux I__17964 (
            .O(N__73155),
            .I(N__72833));
    ClkMux I__17963 (
            .O(N__73154),
            .I(N__72833));
    ClkMux I__17962 (
            .O(N__73153),
            .I(N__72833));
    ClkMux I__17961 (
            .O(N__73152),
            .I(N__72833));
    ClkMux I__17960 (
            .O(N__73151),
            .I(N__72833));
    ClkMux I__17959 (
            .O(N__73150),
            .I(N__72833));
    ClkMux I__17958 (
            .O(N__73149),
            .I(N__72833));
    ClkMux I__17957 (
            .O(N__73148),
            .I(N__72833));
    ClkMux I__17956 (
            .O(N__73147),
            .I(N__72833));
    ClkMux I__17955 (
            .O(N__73146),
            .I(N__72833));
    ClkMux I__17954 (
            .O(N__73145),
            .I(N__72833));
    ClkMux I__17953 (
            .O(N__73144),
            .I(N__72833));
    ClkMux I__17952 (
            .O(N__73143),
            .I(N__72833));
    ClkMux I__17951 (
            .O(N__73142),
            .I(N__72833));
    ClkMux I__17950 (
            .O(N__73141),
            .I(N__72833));
    ClkMux I__17949 (
            .O(N__73140),
            .I(N__72833));
    ClkMux I__17948 (
            .O(N__73139),
            .I(N__72833));
    ClkMux I__17947 (
            .O(N__73138),
            .I(N__72833));
    GlobalMux I__17946 (
            .O(N__72833),
            .I(N__72830));
    gio2CtrlBuf I__17945 (
            .O(N__72830),
            .I(CLK_c_g));
    InMux I__17944 (
            .O(N__72827),
            .I(N__72824));
    LocalMux I__17943 (
            .O(N__72824),
            .I(N__72821));
    Span4Mux_v I__17942 (
            .O(N__72821),
            .I(N__72818));
    Odrv4 I__17941 (
            .O(N__72818),
            .I(\PROM.ROMDATA.m181 ));
    InMux I__17940 (
            .O(N__72815),
            .I(N__72812));
    LocalMux I__17939 (
            .O(N__72812),
            .I(\PROM.ROMDATA.m480_bm ));
    CascadeMux I__17938 (
            .O(N__72809),
            .I(\PROM.ROMDATA.m480_am_cascade_ ));
    InMux I__17937 (
            .O(N__72806),
            .I(N__72803));
    LocalMux I__17936 (
            .O(N__72803),
            .I(N__72800));
    Span4Mux_h I__17935 (
            .O(N__72800),
            .I(N__72797));
    Span4Mux_h I__17934 (
            .O(N__72797),
            .I(N__72794));
    Odrv4 I__17933 (
            .O(N__72794),
            .I(\PROM.ROMDATA.N_551_mux ));
    CascadeMux I__17932 (
            .O(N__72791),
            .I(N__72786));
    CascadeMux I__17931 (
            .O(N__72790),
            .I(N__72781));
    CascadeMux I__17930 (
            .O(N__72789),
            .I(N__72778));
    InMux I__17929 (
            .O(N__72786),
            .I(N__72761));
    InMux I__17928 (
            .O(N__72785),
            .I(N__72761));
    InMux I__17927 (
            .O(N__72784),
            .I(N__72761));
    InMux I__17926 (
            .O(N__72781),
            .I(N__72752));
    InMux I__17925 (
            .O(N__72778),
            .I(N__72752));
    InMux I__17924 (
            .O(N__72777),
            .I(N__72752));
    InMux I__17923 (
            .O(N__72776),
            .I(N__72752));
    InMux I__17922 (
            .O(N__72775),
            .I(N__72749));
    InMux I__17921 (
            .O(N__72774),
            .I(N__72746));
    InMux I__17920 (
            .O(N__72773),
            .I(N__72743));
    CascadeMux I__17919 (
            .O(N__72772),
            .I(N__72738));
    InMux I__17918 (
            .O(N__72771),
            .I(N__72732));
    InMux I__17917 (
            .O(N__72770),
            .I(N__72732));
    CascadeMux I__17916 (
            .O(N__72769),
            .I(N__72717));
    CascadeMux I__17915 (
            .O(N__72768),
            .I(N__72714));
    LocalMux I__17914 (
            .O(N__72761),
            .I(N__72707));
    LocalMux I__17913 (
            .O(N__72752),
            .I(N__72707));
    LocalMux I__17912 (
            .O(N__72749),
            .I(N__72704));
    LocalMux I__17911 (
            .O(N__72746),
            .I(N__72699));
    LocalMux I__17910 (
            .O(N__72743),
            .I(N__72699));
    CascadeMux I__17909 (
            .O(N__72742),
            .I(N__72685));
    InMux I__17908 (
            .O(N__72741),
            .I(N__72676));
    InMux I__17907 (
            .O(N__72738),
            .I(N__72676));
    InMux I__17906 (
            .O(N__72737),
            .I(N__72673));
    LocalMux I__17905 (
            .O(N__72732),
            .I(N__72669));
    InMux I__17904 (
            .O(N__72731),
            .I(N__72666));
    InMux I__17903 (
            .O(N__72730),
            .I(N__72657));
    InMux I__17902 (
            .O(N__72729),
            .I(N__72657));
    InMux I__17901 (
            .O(N__72728),
            .I(N__72657));
    InMux I__17900 (
            .O(N__72727),
            .I(N__72657));
    CascadeMux I__17899 (
            .O(N__72726),
            .I(N__72652));
    CascadeMux I__17898 (
            .O(N__72725),
            .I(N__72649));
    InMux I__17897 (
            .O(N__72724),
            .I(N__72637));
    InMux I__17896 (
            .O(N__72723),
            .I(N__72637));
    InMux I__17895 (
            .O(N__72722),
            .I(N__72637));
    InMux I__17894 (
            .O(N__72721),
            .I(N__72637));
    InMux I__17893 (
            .O(N__72720),
            .I(N__72637));
    InMux I__17892 (
            .O(N__72717),
            .I(N__72630));
    InMux I__17891 (
            .O(N__72714),
            .I(N__72630));
    InMux I__17890 (
            .O(N__72713),
            .I(N__72630));
    InMux I__17889 (
            .O(N__72712),
            .I(N__72627));
    Span4Mux_v I__17888 (
            .O(N__72707),
            .I(N__72619));
    Span4Mux_v I__17887 (
            .O(N__72704),
            .I(N__72619));
    Span4Mux_v I__17886 (
            .O(N__72699),
            .I(N__72619));
    CascadeMux I__17885 (
            .O(N__72698),
            .I(N__72615));
    InMux I__17884 (
            .O(N__72697),
            .I(N__72612));
    InMux I__17883 (
            .O(N__72696),
            .I(N__72609));
    InMux I__17882 (
            .O(N__72695),
            .I(N__72603));
    InMux I__17881 (
            .O(N__72694),
            .I(N__72600));
    InMux I__17880 (
            .O(N__72693),
            .I(N__72597));
    InMux I__17879 (
            .O(N__72692),
            .I(N__72588));
    InMux I__17878 (
            .O(N__72691),
            .I(N__72588));
    InMux I__17877 (
            .O(N__72690),
            .I(N__72588));
    InMux I__17876 (
            .O(N__72689),
            .I(N__72588));
    InMux I__17875 (
            .O(N__72688),
            .I(N__72583));
    InMux I__17874 (
            .O(N__72685),
            .I(N__72583));
    InMux I__17873 (
            .O(N__72684),
            .I(N__72580));
    InMux I__17872 (
            .O(N__72683),
            .I(N__72577));
    InMux I__17871 (
            .O(N__72682),
            .I(N__72572));
    InMux I__17870 (
            .O(N__72681),
            .I(N__72572));
    LocalMux I__17869 (
            .O(N__72676),
            .I(N__72567));
    LocalMux I__17868 (
            .O(N__72673),
            .I(N__72567));
    CascadeMux I__17867 (
            .O(N__72672),
            .I(N__72564));
    Span4Mux_h I__17866 (
            .O(N__72669),
            .I(N__72560));
    LocalMux I__17865 (
            .O(N__72666),
            .I(N__72557));
    LocalMux I__17864 (
            .O(N__72657),
            .I(N__72554));
    InMux I__17863 (
            .O(N__72656),
            .I(N__72549));
    InMux I__17862 (
            .O(N__72655),
            .I(N__72549));
    InMux I__17861 (
            .O(N__72652),
            .I(N__72546));
    InMux I__17860 (
            .O(N__72649),
            .I(N__72541));
    InMux I__17859 (
            .O(N__72648),
            .I(N__72541));
    LocalMux I__17858 (
            .O(N__72637),
            .I(N__72538));
    LocalMux I__17857 (
            .O(N__72630),
            .I(N__72535));
    LocalMux I__17856 (
            .O(N__72627),
            .I(N__72532));
    CascadeMux I__17855 (
            .O(N__72626),
            .I(N__72529));
    Span4Mux_h I__17854 (
            .O(N__72619),
            .I(N__72526));
    InMux I__17853 (
            .O(N__72618),
            .I(N__72523));
    InMux I__17852 (
            .O(N__72615),
            .I(N__72520));
    LocalMux I__17851 (
            .O(N__72612),
            .I(N__72515));
    LocalMux I__17850 (
            .O(N__72609),
            .I(N__72515));
    InMux I__17849 (
            .O(N__72608),
            .I(N__72512));
    CascadeMux I__17848 (
            .O(N__72607),
            .I(N__72508));
    CascadeMux I__17847 (
            .O(N__72606),
            .I(N__72505));
    LocalMux I__17846 (
            .O(N__72603),
            .I(N__72500));
    LocalMux I__17845 (
            .O(N__72600),
            .I(N__72495));
    LocalMux I__17844 (
            .O(N__72597),
            .I(N__72495));
    LocalMux I__17843 (
            .O(N__72588),
            .I(N__72490));
    LocalMux I__17842 (
            .O(N__72583),
            .I(N__72490));
    LocalMux I__17841 (
            .O(N__72580),
            .I(N__72485));
    LocalMux I__17840 (
            .O(N__72577),
            .I(N__72485));
    LocalMux I__17839 (
            .O(N__72572),
            .I(N__72480));
    Span4Mux_v I__17838 (
            .O(N__72567),
            .I(N__72480));
    InMux I__17837 (
            .O(N__72564),
            .I(N__72475));
    InMux I__17836 (
            .O(N__72563),
            .I(N__72475));
    Span4Mux_v I__17835 (
            .O(N__72560),
            .I(N__72470));
    Span4Mux_v I__17834 (
            .O(N__72557),
            .I(N__72470));
    Span4Mux_v I__17833 (
            .O(N__72554),
            .I(N__72461));
    LocalMux I__17832 (
            .O(N__72549),
            .I(N__72461));
    LocalMux I__17831 (
            .O(N__72546),
            .I(N__72461));
    LocalMux I__17830 (
            .O(N__72541),
            .I(N__72461));
    Span4Mux_v I__17829 (
            .O(N__72538),
            .I(N__72454));
    Span4Mux_h I__17828 (
            .O(N__72535),
            .I(N__72454));
    Span4Mux_h I__17827 (
            .O(N__72532),
            .I(N__72454));
    InMux I__17826 (
            .O(N__72529),
            .I(N__72451));
    Span4Mux_h I__17825 (
            .O(N__72526),
            .I(N__72446));
    LocalMux I__17824 (
            .O(N__72523),
            .I(N__72446));
    LocalMux I__17823 (
            .O(N__72520),
            .I(N__72439));
    Span12Mux_h I__17822 (
            .O(N__72515),
            .I(N__72439));
    LocalMux I__17821 (
            .O(N__72512),
            .I(N__72439));
    InMux I__17820 (
            .O(N__72511),
            .I(N__72436));
    InMux I__17819 (
            .O(N__72508),
            .I(N__72433));
    InMux I__17818 (
            .O(N__72505),
            .I(N__72430));
    InMux I__17817 (
            .O(N__72504),
            .I(N__72427));
    InMux I__17816 (
            .O(N__72503),
            .I(N__72424));
    Span4Mux_h I__17815 (
            .O(N__72500),
            .I(N__72415));
    Span4Mux_v I__17814 (
            .O(N__72495),
            .I(N__72415));
    Span4Mux_v I__17813 (
            .O(N__72490),
            .I(N__72415));
    Span4Mux_h I__17812 (
            .O(N__72485),
            .I(N__72415));
    Span4Mux_h I__17811 (
            .O(N__72480),
            .I(N__72404));
    LocalMux I__17810 (
            .O(N__72475),
            .I(N__72404));
    Span4Mux_h I__17809 (
            .O(N__72470),
            .I(N__72404));
    Span4Mux_v I__17808 (
            .O(N__72461),
            .I(N__72404));
    Span4Mux_v I__17807 (
            .O(N__72454),
            .I(N__72404));
    LocalMux I__17806 (
            .O(N__72451),
            .I(progRomAddress_7));
    Odrv4 I__17805 (
            .O(N__72446),
            .I(progRomAddress_7));
    Odrv12 I__17804 (
            .O(N__72439),
            .I(progRomAddress_7));
    LocalMux I__17803 (
            .O(N__72436),
            .I(progRomAddress_7));
    LocalMux I__17802 (
            .O(N__72433),
            .I(progRomAddress_7));
    LocalMux I__17801 (
            .O(N__72430),
            .I(progRomAddress_7));
    LocalMux I__17800 (
            .O(N__72427),
            .I(progRomAddress_7));
    LocalMux I__17799 (
            .O(N__72424),
            .I(progRomAddress_7));
    Odrv4 I__17798 (
            .O(N__72415),
            .I(progRomAddress_7));
    Odrv4 I__17797 (
            .O(N__72404),
            .I(progRomAddress_7));
    CascadeMux I__17796 (
            .O(N__72383),
            .I(\PROM.ROMDATA.m480_ns_cascade_ ));
    InMux I__17795 (
            .O(N__72380),
            .I(N__72377));
    LocalMux I__17794 (
            .O(N__72377),
            .I(N__72373));
    InMux I__17793 (
            .O(N__72376),
            .I(N__72370));
    Span4Mux_h I__17792 (
            .O(N__72373),
            .I(N__72367));
    LocalMux I__17791 (
            .O(N__72370),
            .I(N__72364));
    Span4Mux_h I__17790 (
            .O(N__72367),
            .I(N__72361));
    Span12Mux_h I__17789 (
            .O(N__72364),
            .I(N__72358));
    Odrv4 I__17788 (
            .O(N__72361),
            .I(PROM_ROMDATA_dintern_25ro));
    Odrv12 I__17787 (
            .O(N__72358),
            .I(PROM_ROMDATA_dintern_25ro));
    InMux I__17786 (
            .O(N__72353),
            .I(N__72349));
    InMux I__17785 (
            .O(N__72352),
            .I(N__72345));
    LocalMux I__17784 (
            .O(N__72349),
            .I(N__72342));
    InMux I__17783 (
            .O(N__72348),
            .I(N__72339));
    LocalMux I__17782 (
            .O(N__72345),
            .I(N__72336));
    Span4Mux_h I__17781 (
            .O(N__72342),
            .I(N__72331));
    LocalMux I__17780 (
            .O(N__72339),
            .I(N__72331));
    Span4Mux_h I__17779 (
            .O(N__72336),
            .I(N__72328));
    Span4Mux_h I__17778 (
            .O(N__72331),
            .I(N__72325));
    Odrv4 I__17777 (
            .O(N__72328),
            .I(g_9));
    Odrv4 I__17776 (
            .O(N__72325),
            .I(g_9));
    CascadeMux I__17775 (
            .O(N__72320),
            .I(N__72312));
    CascadeMux I__17774 (
            .O(N__72319),
            .I(N__72308));
    InMux I__17773 (
            .O(N__72318),
            .I(N__72301));
    CascadeMux I__17772 (
            .O(N__72317),
            .I(N__72294));
    CascadeMux I__17771 (
            .O(N__72316),
            .I(N__72290));
    CascadeMux I__17770 (
            .O(N__72315),
            .I(N__72285));
    InMux I__17769 (
            .O(N__72312),
            .I(N__72281));
    InMux I__17768 (
            .O(N__72311),
            .I(N__72274));
    InMux I__17767 (
            .O(N__72308),
            .I(N__72274));
    InMux I__17766 (
            .O(N__72307),
            .I(N__72274));
    CascadeMux I__17765 (
            .O(N__72306),
            .I(N__72268));
    CascadeMux I__17764 (
            .O(N__72305),
            .I(N__72265));
    InMux I__17763 (
            .O(N__72304),
            .I(N__72257));
    LocalMux I__17762 (
            .O(N__72301),
            .I(N__72253));
    InMux I__17761 (
            .O(N__72300),
            .I(N__72244));
    InMux I__17760 (
            .O(N__72299),
            .I(N__72239));
    InMux I__17759 (
            .O(N__72298),
            .I(N__72239));
    InMux I__17758 (
            .O(N__72297),
            .I(N__72236));
    InMux I__17757 (
            .O(N__72294),
            .I(N__72231));
    InMux I__17756 (
            .O(N__72293),
            .I(N__72231));
    InMux I__17755 (
            .O(N__72290),
            .I(N__72228));
    CascadeMux I__17754 (
            .O(N__72289),
            .I(N__72217));
    CascadeMux I__17753 (
            .O(N__72288),
            .I(N__72214));
    InMux I__17752 (
            .O(N__72285),
            .I(N__72209));
    CascadeMux I__17751 (
            .O(N__72284),
            .I(N__72206));
    LocalMux I__17750 (
            .O(N__72281),
            .I(N__72201));
    LocalMux I__17749 (
            .O(N__72274),
            .I(N__72201));
    InMux I__17748 (
            .O(N__72273),
            .I(N__72198));
    InMux I__17747 (
            .O(N__72272),
            .I(N__72195));
    InMux I__17746 (
            .O(N__72271),
            .I(N__72185));
    InMux I__17745 (
            .O(N__72268),
            .I(N__72182));
    InMux I__17744 (
            .O(N__72265),
            .I(N__72171));
    InMux I__17743 (
            .O(N__72264),
            .I(N__72171));
    InMux I__17742 (
            .O(N__72263),
            .I(N__72166));
    InMux I__17741 (
            .O(N__72262),
            .I(N__72166));
    InMux I__17740 (
            .O(N__72261),
            .I(N__72161));
    InMux I__17739 (
            .O(N__72260),
            .I(N__72161));
    LocalMux I__17738 (
            .O(N__72257),
            .I(N__72158));
    InMux I__17737 (
            .O(N__72256),
            .I(N__72155));
    Span4Mux_h I__17736 (
            .O(N__72253),
            .I(N__72152));
    InMux I__17735 (
            .O(N__72252),
            .I(N__72149));
    InMux I__17734 (
            .O(N__72251),
            .I(N__72146));
    InMux I__17733 (
            .O(N__72250),
            .I(N__72141));
    InMux I__17732 (
            .O(N__72249),
            .I(N__72141));
    InMux I__17731 (
            .O(N__72248),
            .I(N__72137));
    InMux I__17730 (
            .O(N__72247),
            .I(N__72134));
    LocalMux I__17729 (
            .O(N__72244),
            .I(N__72123));
    LocalMux I__17728 (
            .O(N__72239),
            .I(N__72123));
    LocalMux I__17727 (
            .O(N__72236),
            .I(N__72118));
    LocalMux I__17726 (
            .O(N__72231),
            .I(N__72118));
    LocalMux I__17725 (
            .O(N__72228),
            .I(N__72115));
    InMux I__17724 (
            .O(N__72227),
            .I(N__72110));
    InMux I__17723 (
            .O(N__72226),
            .I(N__72110));
    InMux I__17722 (
            .O(N__72225),
            .I(N__72105));
    InMux I__17721 (
            .O(N__72224),
            .I(N__72105));
    InMux I__17720 (
            .O(N__72223),
            .I(N__72097));
    InMux I__17719 (
            .O(N__72222),
            .I(N__72092));
    InMux I__17718 (
            .O(N__72221),
            .I(N__72092));
    InMux I__17717 (
            .O(N__72220),
            .I(N__72081));
    InMux I__17716 (
            .O(N__72217),
            .I(N__72081));
    InMux I__17715 (
            .O(N__72214),
            .I(N__72081));
    InMux I__17714 (
            .O(N__72213),
            .I(N__72081));
    InMux I__17713 (
            .O(N__72212),
            .I(N__72081));
    LocalMux I__17712 (
            .O(N__72209),
            .I(N__72078));
    InMux I__17711 (
            .O(N__72206),
            .I(N__72075));
    Span4Mux_v I__17710 (
            .O(N__72201),
            .I(N__72068));
    LocalMux I__17709 (
            .O(N__72198),
            .I(N__72068));
    LocalMux I__17708 (
            .O(N__72195),
            .I(N__72068));
    InMux I__17707 (
            .O(N__72194),
            .I(N__72061));
    InMux I__17706 (
            .O(N__72193),
            .I(N__72061));
    InMux I__17705 (
            .O(N__72192),
            .I(N__72061));
    InMux I__17704 (
            .O(N__72191),
            .I(N__72052));
    InMux I__17703 (
            .O(N__72190),
            .I(N__72052));
    InMux I__17702 (
            .O(N__72189),
            .I(N__72052));
    InMux I__17701 (
            .O(N__72188),
            .I(N__72052));
    LocalMux I__17700 (
            .O(N__72185),
            .I(N__72047));
    LocalMux I__17699 (
            .O(N__72182),
            .I(N__72047));
    InMux I__17698 (
            .O(N__72181),
            .I(N__72044));
    InMux I__17697 (
            .O(N__72180),
            .I(N__72033));
    InMux I__17696 (
            .O(N__72179),
            .I(N__72033));
    InMux I__17695 (
            .O(N__72178),
            .I(N__72033));
    InMux I__17694 (
            .O(N__72177),
            .I(N__72033));
    InMux I__17693 (
            .O(N__72176),
            .I(N__72033));
    LocalMux I__17692 (
            .O(N__72171),
            .I(N__72026));
    LocalMux I__17691 (
            .O(N__72166),
            .I(N__72026));
    LocalMux I__17690 (
            .O(N__72161),
            .I(N__72026));
    Span4Mux_h I__17689 (
            .O(N__72158),
            .I(N__72013));
    LocalMux I__17688 (
            .O(N__72155),
            .I(N__72013));
    Span4Mux_h I__17687 (
            .O(N__72152),
            .I(N__72013));
    LocalMux I__17686 (
            .O(N__72149),
            .I(N__72013));
    LocalMux I__17685 (
            .O(N__72146),
            .I(N__72013));
    LocalMux I__17684 (
            .O(N__72141),
            .I(N__72013));
    CascadeMux I__17683 (
            .O(N__72140),
            .I(N__72010));
    LocalMux I__17682 (
            .O(N__72137),
            .I(N__72005));
    LocalMux I__17681 (
            .O(N__72134),
            .I(N__72002));
    InMux I__17680 (
            .O(N__72133),
            .I(N__71997));
    InMux I__17679 (
            .O(N__72132),
            .I(N__71997));
    InMux I__17678 (
            .O(N__72131),
            .I(N__71994));
    InMux I__17677 (
            .O(N__72130),
            .I(N__71987));
    InMux I__17676 (
            .O(N__72129),
            .I(N__71987));
    InMux I__17675 (
            .O(N__72128),
            .I(N__71987));
    Span12Mux_h I__17674 (
            .O(N__72123),
            .I(N__71976));
    Sp12to4 I__17673 (
            .O(N__72118),
            .I(N__71976));
    Sp12to4 I__17672 (
            .O(N__72115),
            .I(N__71976));
    LocalMux I__17671 (
            .O(N__72110),
            .I(N__71976));
    LocalMux I__17670 (
            .O(N__72105),
            .I(N__71976));
    InMux I__17669 (
            .O(N__72104),
            .I(N__71973));
    InMux I__17668 (
            .O(N__72103),
            .I(N__71968));
    InMux I__17667 (
            .O(N__72102),
            .I(N__71968));
    InMux I__17666 (
            .O(N__72101),
            .I(N__71963));
    InMux I__17665 (
            .O(N__72100),
            .I(N__71963));
    LocalMux I__17664 (
            .O(N__72097),
            .I(N__71960));
    LocalMux I__17663 (
            .O(N__72092),
            .I(N__71951));
    LocalMux I__17662 (
            .O(N__72081),
            .I(N__71951));
    Span4Mux_h I__17661 (
            .O(N__72078),
            .I(N__71951));
    LocalMux I__17660 (
            .O(N__72075),
            .I(N__71951));
    Span4Mux_v I__17659 (
            .O(N__72068),
            .I(N__71948));
    LocalMux I__17658 (
            .O(N__72061),
            .I(N__71935));
    LocalMux I__17657 (
            .O(N__72052),
            .I(N__71935));
    Span4Mux_v I__17656 (
            .O(N__72047),
            .I(N__71935));
    LocalMux I__17655 (
            .O(N__72044),
            .I(N__71935));
    LocalMux I__17654 (
            .O(N__72033),
            .I(N__71935));
    Span4Mux_h I__17653 (
            .O(N__72026),
            .I(N__71935));
    Span4Mux_h I__17652 (
            .O(N__72013),
            .I(N__71932));
    InMux I__17651 (
            .O(N__72010),
            .I(N__71925));
    InMux I__17650 (
            .O(N__72009),
            .I(N__71925));
    InMux I__17649 (
            .O(N__72008),
            .I(N__71925));
    Span4Mux_v I__17648 (
            .O(N__72005),
            .I(N__71922));
    Span4Mux_h I__17647 (
            .O(N__72002),
            .I(N__71915));
    LocalMux I__17646 (
            .O(N__71997),
            .I(N__71915));
    LocalMux I__17645 (
            .O(N__71994),
            .I(N__71915));
    LocalMux I__17644 (
            .O(N__71987),
            .I(N__71910));
    Span12Mux_v I__17643 (
            .O(N__71976),
            .I(N__71910));
    LocalMux I__17642 (
            .O(N__71973),
            .I(N__71895));
    LocalMux I__17641 (
            .O(N__71968),
            .I(N__71895));
    LocalMux I__17640 (
            .O(N__71963),
            .I(N__71895));
    Span4Mux_v I__17639 (
            .O(N__71960),
            .I(N__71895));
    Span4Mux_v I__17638 (
            .O(N__71951),
            .I(N__71895));
    Span4Mux_h I__17637 (
            .O(N__71948),
            .I(N__71895));
    Span4Mux_v I__17636 (
            .O(N__71935),
            .I(N__71895));
    Span4Mux_h I__17635 (
            .O(N__71932),
            .I(N__71892));
    LocalMux I__17634 (
            .O(N__71925),
            .I(PROM_ROMDATA_dintern_adflt));
    Odrv4 I__17633 (
            .O(N__71922),
            .I(PROM_ROMDATA_dintern_adflt));
    Odrv4 I__17632 (
            .O(N__71915),
            .I(PROM_ROMDATA_dintern_adflt));
    Odrv12 I__17631 (
            .O(N__71910),
            .I(PROM_ROMDATA_dintern_adflt));
    Odrv4 I__17630 (
            .O(N__71895),
            .I(PROM_ROMDATA_dintern_adflt));
    Odrv4 I__17629 (
            .O(N__71892),
            .I(PROM_ROMDATA_dintern_adflt));
    CascadeMux I__17628 (
            .O(N__71879),
            .I(PROM_ROMDATA_dintern_25ro_cascade_));
    CascadeMux I__17627 (
            .O(N__71876),
            .I(N__71863));
    InMux I__17626 (
            .O(N__71875),
            .I(N__71860));
    InMux I__17625 (
            .O(N__71874),
            .I(N__71855));
    InMux I__17624 (
            .O(N__71873),
            .I(N__71855));
    InMux I__17623 (
            .O(N__71872),
            .I(N__71849));
    InMux I__17622 (
            .O(N__71871),
            .I(N__71842));
    InMux I__17621 (
            .O(N__71870),
            .I(N__71842));
    InMux I__17620 (
            .O(N__71869),
            .I(N__71842));
    InMux I__17619 (
            .O(N__71868),
            .I(N__71835));
    InMux I__17618 (
            .O(N__71867),
            .I(N__71835));
    InMux I__17617 (
            .O(N__71866),
            .I(N__71835));
    InMux I__17616 (
            .O(N__71863),
            .I(N__71832));
    LocalMux I__17615 (
            .O(N__71860),
            .I(N__71816));
    LocalMux I__17614 (
            .O(N__71855),
            .I(N__71813));
    InMux I__17613 (
            .O(N__71854),
            .I(N__71810));
    CascadeMux I__17612 (
            .O(N__71853),
            .I(N__71807));
    CascadeMux I__17611 (
            .O(N__71852),
            .I(N__71799));
    LocalMux I__17610 (
            .O(N__71849),
            .I(N__71792));
    LocalMux I__17609 (
            .O(N__71842),
            .I(N__71792));
    LocalMux I__17608 (
            .O(N__71835),
            .I(N__71792));
    LocalMux I__17607 (
            .O(N__71832),
            .I(N__71789));
    InMux I__17606 (
            .O(N__71831),
            .I(N__71786));
    InMux I__17605 (
            .O(N__71830),
            .I(N__71783));
    InMux I__17604 (
            .O(N__71829),
            .I(N__71776));
    InMux I__17603 (
            .O(N__71828),
            .I(N__71776));
    InMux I__17602 (
            .O(N__71827),
            .I(N__71776));
    InMux I__17601 (
            .O(N__71826),
            .I(N__71765));
    InMux I__17600 (
            .O(N__71825),
            .I(N__71765));
    InMux I__17599 (
            .O(N__71824),
            .I(N__71765));
    InMux I__17598 (
            .O(N__71823),
            .I(N__71765));
    InMux I__17597 (
            .O(N__71822),
            .I(N__71765));
    CascadeMux I__17596 (
            .O(N__71821),
            .I(N__71762));
    InMux I__17595 (
            .O(N__71820),
            .I(N__71759));
    CascadeMux I__17594 (
            .O(N__71819),
            .I(N__71755));
    Span4Mux_h I__17593 (
            .O(N__71816),
            .I(N__71752));
    Span4Mux_v I__17592 (
            .O(N__71813),
            .I(N__71749));
    LocalMux I__17591 (
            .O(N__71810),
            .I(N__71746));
    InMux I__17590 (
            .O(N__71807),
            .I(N__71742));
    InMux I__17589 (
            .O(N__71806),
            .I(N__71739));
    InMux I__17588 (
            .O(N__71805),
            .I(N__71730));
    InMux I__17587 (
            .O(N__71804),
            .I(N__71730));
    InMux I__17586 (
            .O(N__71803),
            .I(N__71730));
    InMux I__17585 (
            .O(N__71802),
            .I(N__71730));
    InMux I__17584 (
            .O(N__71799),
            .I(N__71727));
    Span4Mux_v I__17583 (
            .O(N__71792),
            .I(N__71722));
    Span4Mux_v I__17582 (
            .O(N__71789),
            .I(N__71722));
    LocalMux I__17581 (
            .O(N__71786),
            .I(N__71715));
    LocalMux I__17580 (
            .O(N__71783),
            .I(N__71715));
    LocalMux I__17579 (
            .O(N__71776),
            .I(N__71715));
    LocalMux I__17578 (
            .O(N__71765),
            .I(N__71712));
    InMux I__17577 (
            .O(N__71762),
            .I(N__71709));
    LocalMux I__17576 (
            .O(N__71759),
            .I(N__71706));
    InMux I__17575 (
            .O(N__71758),
            .I(N__71701));
    InMux I__17574 (
            .O(N__71755),
            .I(N__71701));
    Span4Mux_h I__17573 (
            .O(N__71752),
            .I(N__71698));
    Span4Mux_h I__17572 (
            .O(N__71749),
            .I(N__71693));
    Span4Mux_v I__17571 (
            .O(N__71746),
            .I(N__71693));
    InMux I__17570 (
            .O(N__71745),
            .I(N__71690));
    LocalMux I__17569 (
            .O(N__71742),
            .I(N__71683));
    LocalMux I__17568 (
            .O(N__71739),
            .I(N__71683));
    LocalMux I__17567 (
            .O(N__71730),
            .I(N__71683));
    LocalMux I__17566 (
            .O(N__71727),
            .I(N__71676));
    Span4Mux_h I__17565 (
            .O(N__71722),
            .I(N__71676));
    Span4Mux_v I__17564 (
            .O(N__71715),
            .I(N__71676));
    Odrv12 I__17563 (
            .O(N__71712),
            .I(PROM_ROMDATA_dintern_3ro));
    LocalMux I__17562 (
            .O(N__71709),
            .I(PROM_ROMDATA_dintern_3ro));
    Odrv4 I__17561 (
            .O(N__71706),
            .I(PROM_ROMDATA_dintern_3ro));
    LocalMux I__17560 (
            .O(N__71701),
            .I(PROM_ROMDATA_dintern_3ro));
    Odrv4 I__17559 (
            .O(N__71698),
            .I(PROM_ROMDATA_dintern_3ro));
    Odrv4 I__17558 (
            .O(N__71693),
            .I(PROM_ROMDATA_dintern_3ro));
    LocalMux I__17557 (
            .O(N__71690),
            .I(PROM_ROMDATA_dintern_3ro));
    Odrv4 I__17556 (
            .O(N__71683),
            .I(PROM_ROMDATA_dintern_3ro));
    Odrv4 I__17555 (
            .O(N__71676),
            .I(PROM_ROMDATA_dintern_3ro));
    CascadeMux I__17554 (
            .O(N__71657),
            .I(N__71654));
    CascadeBuf I__17553 (
            .O(N__71654),
            .I(N__71651));
    CascadeMux I__17552 (
            .O(N__71651),
            .I(N__71648));
    CascadeBuf I__17551 (
            .O(N__71648),
            .I(N__71645));
    CascadeMux I__17550 (
            .O(N__71645),
            .I(N__71642));
    CascadeBuf I__17549 (
            .O(N__71642),
            .I(N__71639));
    CascadeMux I__17548 (
            .O(N__71639),
            .I(N__71636));
    InMux I__17547 (
            .O(N__71636),
            .I(N__71633));
    LocalMux I__17546 (
            .O(N__71633),
            .I(N__71630));
    Span4Mux_v I__17545 (
            .O(N__71630),
            .I(N__71627));
    Sp12to4 I__17544 (
            .O(N__71627),
            .I(N__71624));
    Span12Mux_v I__17543 (
            .O(N__71624),
            .I(N__71621));
    Span12Mux_h I__17542 (
            .O(N__71621),
            .I(N__71618));
    Odrv12 I__17541 (
            .O(N__71618),
            .I(CONTROL_romAddReg_7_9));
    InMux I__17540 (
            .O(N__71615),
            .I(N__71612));
    LocalMux I__17539 (
            .O(N__71612),
            .I(N__71609));
    Span4Mux_h I__17538 (
            .O(N__71609),
            .I(N__71606));
    Odrv4 I__17537 (
            .O(N__71606),
            .I(\PROM.ROMDATA.m446_bm ));
    InMux I__17536 (
            .O(N__71603),
            .I(N__71600));
    LocalMux I__17535 (
            .O(N__71600),
            .I(N__71597));
    Span4Mux_h I__17534 (
            .O(N__71597),
            .I(N__71594));
    Span4Mux_h I__17533 (
            .O(N__71594),
            .I(N__71591));
    Odrv4 I__17532 (
            .O(N__71591),
            .I(\PROM.ROMDATA.m447_ns_1 ));
    CascadeMux I__17531 (
            .O(N__71588),
            .I(N__71585));
    InMux I__17530 (
            .O(N__71585),
            .I(N__71582));
    LocalMux I__17529 (
            .O(N__71582),
            .I(\PROM.ROMDATA.m446_am ));
    InMux I__17528 (
            .O(N__71579),
            .I(N__71573));
    InMux I__17527 (
            .O(N__71578),
            .I(N__71573));
    LocalMux I__17526 (
            .O(N__71573),
            .I(N__71570));
    Span4Mux_v I__17525 (
            .O(N__71570),
            .I(N__71567));
    Sp12to4 I__17524 (
            .O(N__71567),
            .I(N__71564));
    Span12Mux_h I__17523 (
            .O(N__71564),
            .I(N__71561));
    Odrv12 I__17522 (
            .O(N__71561),
            .I(\PROM.ROMDATA.m447_ns ));
    CEMux I__17521 (
            .O(N__71558),
            .I(N__71555));
    LocalMux I__17520 (
            .O(N__71555),
            .I(N__71550));
    CEMux I__17519 (
            .O(N__71554),
            .I(N__71547));
    CEMux I__17518 (
            .O(N__71553),
            .I(N__71544));
    Span4Mux_h I__17517 (
            .O(N__71550),
            .I(N__71539));
    LocalMux I__17516 (
            .O(N__71547),
            .I(N__71539));
    LocalMux I__17515 (
            .O(N__71544),
            .I(N__71536));
    Span4Mux_h I__17514 (
            .O(N__71539),
            .I(N__71533));
    Span4Mux_v I__17513 (
            .O(N__71536),
            .I(N__71530));
    Span4Mux_h I__17512 (
            .O(N__71533),
            .I(N__71527));
    Span4Mux_h I__17511 (
            .O(N__71530),
            .I(N__71522));
    Span4Mux_h I__17510 (
            .O(N__71527),
            .I(N__71522));
    Odrv4 I__17509 (
            .O(N__71522),
            .I(\ALU.un1_a41_7_0 ));
    InMux I__17508 (
            .O(N__71519),
            .I(N__71516));
    LocalMux I__17507 (
            .O(N__71516),
            .I(N__71512));
    InMux I__17506 (
            .O(N__71515),
            .I(N__71509));
    Odrv4 I__17505 (
            .O(N__71512),
            .I(\ALU.un1_operation_13Z0Z_2 ));
    LocalMux I__17504 (
            .O(N__71509),
            .I(\ALU.un1_operation_13Z0Z_2 ));
    CascadeMux I__17503 (
            .O(N__71504),
            .I(N__71501));
    InMux I__17502 (
            .O(N__71501),
            .I(N__71495));
    InMux I__17501 (
            .O(N__71500),
            .I(N__71495));
    LocalMux I__17500 (
            .O(N__71495),
            .I(N__71492));
    Sp12to4 I__17499 (
            .O(N__71492),
            .I(N__71487));
    InMux I__17498 (
            .O(N__71491),
            .I(N__71484));
    InMux I__17497 (
            .O(N__71490),
            .I(N__71481));
    Span12Mux_v I__17496 (
            .O(N__71487),
            .I(N__71478));
    LocalMux I__17495 (
            .O(N__71484),
            .I(\ALU.un1_operation_10_0 ));
    LocalMux I__17494 (
            .O(N__71481),
            .I(\ALU.un1_operation_10_0 ));
    Odrv12 I__17493 (
            .O(N__71478),
            .I(\ALU.un1_operation_10_0 ));
    InMux I__17492 (
            .O(N__71471),
            .I(N__71464));
    InMux I__17491 (
            .O(N__71470),
            .I(N__71460));
    InMux I__17490 (
            .O(N__71469),
            .I(N__71455));
    InMux I__17489 (
            .O(N__71468),
            .I(N__71455));
    InMux I__17488 (
            .O(N__71467),
            .I(N__71445));
    LocalMux I__17487 (
            .O(N__71464),
            .I(N__71442));
    InMux I__17486 (
            .O(N__71463),
            .I(N__71437));
    LocalMux I__17485 (
            .O(N__71460),
            .I(N__71432));
    LocalMux I__17484 (
            .O(N__71455),
            .I(N__71429));
    InMux I__17483 (
            .O(N__71454),
            .I(N__71426));
    InMux I__17482 (
            .O(N__71453),
            .I(N__71418));
    InMux I__17481 (
            .O(N__71452),
            .I(N__71418));
    InMux I__17480 (
            .O(N__71451),
            .I(N__71411));
    InMux I__17479 (
            .O(N__71450),
            .I(N__71411));
    InMux I__17478 (
            .O(N__71449),
            .I(N__71411));
    CascadeMux I__17477 (
            .O(N__71448),
            .I(N__71407));
    LocalMux I__17476 (
            .O(N__71445),
            .I(N__71402));
    Span4Mux_v I__17475 (
            .O(N__71442),
            .I(N__71402));
    InMux I__17474 (
            .O(N__71441),
            .I(N__71396));
    InMux I__17473 (
            .O(N__71440),
            .I(N__71391));
    LocalMux I__17472 (
            .O(N__71437),
            .I(N__71388));
    InMux I__17471 (
            .O(N__71436),
            .I(N__71385));
    CascadeMux I__17470 (
            .O(N__71435),
            .I(N__71381));
    Span4Mux_v I__17469 (
            .O(N__71432),
            .I(N__71377));
    Span4Mux_h I__17468 (
            .O(N__71429),
            .I(N__71372));
    LocalMux I__17467 (
            .O(N__71426),
            .I(N__71372));
    InMux I__17466 (
            .O(N__71425),
            .I(N__71367));
    InMux I__17465 (
            .O(N__71424),
            .I(N__71367));
    InMux I__17464 (
            .O(N__71423),
            .I(N__71364));
    LocalMux I__17463 (
            .O(N__71418),
            .I(N__71361));
    LocalMux I__17462 (
            .O(N__71411),
            .I(N__71358));
    InMux I__17461 (
            .O(N__71410),
            .I(N__71353));
    InMux I__17460 (
            .O(N__71407),
            .I(N__71353));
    Span4Mux_v I__17459 (
            .O(N__71402),
            .I(N__71350));
    InMux I__17458 (
            .O(N__71401),
            .I(N__71347));
    InMux I__17457 (
            .O(N__71400),
            .I(N__71344));
    InMux I__17456 (
            .O(N__71399),
            .I(N__71341));
    LocalMux I__17455 (
            .O(N__71396),
            .I(N__71338));
    InMux I__17454 (
            .O(N__71395),
            .I(N__71333));
    InMux I__17453 (
            .O(N__71394),
            .I(N__71333));
    LocalMux I__17452 (
            .O(N__71391),
            .I(N__71330));
    Span4Mux_v I__17451 (
            .O(N__71388),
            .I(N__71327));
    LocalMux I__17450 (
            .O(N__71385),
            .I(N__71324));
    CascadeMux I__17449 (
            .O(N__71384),
            .I(N__71321));
    InMux I__17448 (
            .O(N__71381),
            .I(N__71315));
    InMux I__17447 (
            .O(N__71380),
            .I(N__71315));
    Span4Mux_h I__17446 (
            .O(N__71377),
            .I(N__71309));
    Span4Mux_v I__17445 (
            .O(N__71372),
            .I(N__71309));
    LocalMux I__17444 (
            .O(N__71367),
            .I(N__71304));
    LocalMux I__17443 (
            .O(N__71364),
            .I(N__71304));
    Span4Mux_v I__17442 (
            .O(N__71361),
            .I(N__71297));
    Span4Mux_h I__17441 (
            .O(N__71358),
            .I(N__71297));
    LocalMux I__17440 (
            .O(N__71353),
            .I(N__71297));
    Span4Mux_v I__17439 (
            .O(N__71350),
            .I(N__71292));
    LocalMux I__17438 (
            .O(N__71347),
            .I(N__71292));
    LocalMux I__17437 (
            .O(N__71344),
            .I(N__71289));
    LocalMux I__17436 (
            .O(N__71341),
            .I(N__71282));
    Span4Mux_h I__17435 (
            .O(N__71338),
            .I(N__71282));
    LocalMux I__17434 (
            .O(N__71333),
            .I(N__71282));
    Span4Mux_v I__17433 (
            .O(N__71330),
            .I(N__71279));
    Span4Mux_h I__17432 (
            .O(N__71327),
            .I(N__71274));
    Span4Mux_v I__17431 (
            .O(N__71324),
            .I(N__71274));
    InMux I__17430 (
            .O(N__71321),
            .I(N__71269));
    InMux I__17429 (
            .O(N__71320),
            .I(N__71269));
    LocalMux I__17428 (
            .O(N__71315),
            .I(N__71266));
    InMux I__17427 (
            .O(N__71314),
            .I(N__71263));
    Span4Mux_h I__17426 (
            .O(N__71309),
            .I(N__71260));
    Span4Mux_v I__17425 (
            .O(N__71304),
            .I(N__71257));
    Span4Mux_h I__17424 (
            .O(N__71297),
            .I(N__71254));
    Span4Mux_h I__17423 (
            .O(N__71292),
            .I(N__71251));
    Span4Mux_h I__17422 (
            .O(N__71289),
            .I(N__71248));
    Span4Mux_v I__17421 (
            .O(N__71282),
            .I(N__71245));
    Span4Mux_v I__17420 (
            .O(N__71279),
            .I(N__71236));
    Span4Mux_h I__17419 (
            .O(N__71274),
            .I(N__71236));
    LocalMux I__17418 (
            .O(N__71269),
            .I(N__71236));
    Span4Mux_v I__17417 (
            .O(N__71266),
            .I(N__71236));
    LocalMux I__17416 (
            .O(N__71263),
            .I(aluReadBus));
    Odrv4 I__17415 (
            .O(N__71260),
            .I(aluReadBus));
    Odrv4 I__17414 (
            .O(N__71257),
            .I(aluReadBus));
    Odrv4 I__17413 (
            .O(N__71254),
            .I(aluReadBus));
    Odrv4 I__17412 (
            .O(N__71251),
            .I(aluReadBus));
    Odrv4 I__17411 (
            .O(N__71248),
            .I(aluReadBus));
    Odrv4 I__17410 (
            .O(N__71245),
            .I(aluReadBus));
    Odrv4 I__17409 (
            .O(N__71236),
            .I(aluReadBus));
    CascadeMux I__17408 (
            .O(N__71219),
            .I(\ALU.un1_operation_13_0_cascade_ ));
    CEMux I__17407 (
            .O(N__71216),
            .I(N__71208));
    CEMux I__17406 (
            .O(N__71215),
            .I(N__71204));
    CEMux I__17405 (
            .O(N__71214),
            .I(N__71201));
    CEMux I__17404 (
            .O(N__71213),
            .I(N__71194));
    CEMux I__17403 (
            .O(N__71212),
            .I(N__71190));
    CEMux I__17402 (
            .O(N__71211),
            .I(N__71186));
    LocalMux I__17401 (
            .O(N__71208),
            .I(N__71183));
    CEMux I__17400 (
            .O(N__71207),
            .I(N__71180));
    LocalMux I__17399 (
            .O(N__71204),
            .I(N__71177));
    LocalMux I__17398 (
            .O(N__71201),
            .I(N__71173));
    CEMux I__17397 (
            .O(N__71200),
            .I(N__71170));
    CEMux I__17396 (
            .O(N__71199),
            .I(N__71167));
    CEMux I__17395 (
            .O(N__71198),
            .I(N__71164));
    CEMux I__17394 (
            .O(N__71197),
            .I(N__71160));
    LocalMux I__17393 (
            .O(N__71194),
            .I(N__71157));
    CEMux I__17392 (
            .O(N__71193),
            .I(N__71154));
    LocalMux I__17391 (
            .O(N__71190),
            .I(N__71151));
    CEMux I__17390 (
            .O(N__71189),
            .I(N__71148));
    LocalMux I__17389 (
            .O(N__71186),
            .I(N__71145));
    Span4Mux_h I__17388 (
            .O(N__71183),
            .I(N__71140));
    LocalMux I__17387 (
            .O(N__71180),
            .I(N__71140));
    Span4Mux_v I__17386 (
            .O(N__71177),
            .I(N__71137));
    CEMux I__17385 (
            .O(N__71176),
            .I(N__71134));
    Span4Mux_v I__17384 (
            .O(N__71173),
            .I(N__71131));
    LocalMux I__17383 (
            .O(N__71170),
            .I(N__71128));
    LocalMux I__17382 (
            .O(N__71167),
            .I(N__71125));
    LocalMux I__17381 (
            .O(N__71164),
            .I(N__71122));
    CEMux I__17380 (
            .O(N__71163),
            .I(N__71119));
    LocalMux I__17379 (
            .O(N__71160),
            .I(N__71116));
    Span4Mux_h I__17378 (
            .O(N__71157),
            .I(N__71113));
    LocalMux I__17377 (
            .O(N__71154),
            .I(N__71110));
    Span4Mux_h I__17376 (
            .O(N__71151),
            .I(N__71105));
    LocalMux I__17375 (
            .O(N__71148),
            .I(N__71105));
    Span4Mux_v I__17374 (
            .O(N__71145),
            .I(N__71102));
    Span4Mux_v I__17373 (
            .O(N__71140),
            .I(N__71097));
    Span4Mux_h I__17372 (
            .O(N__71137),
            .I(N__71097));
    LocalMux I__17371 (
            .O(N__71134),
            .I(N__71094));
    Span4Mux_h I__17370 (
            .O(N__71131),
            .I(N__71089));
    Span4Mux_h I__17369 (
            .O(N__71128),
            .I(N__71089));
    Span4Mux_v I__17368 (
            .O(N__71125),
            .I(N__71084));
    Span4Mux_v I__17367 (
            .O(N__71122),
            .I(N__71084));
    LocalMux I__17366 (
            .O(N__71119),
            .I(N__71081));
    Span4Mux_v I__17365 (
            .O(N__71116),
            .I(N__71076));
    Span4Mux_h I__17364 (
            .O(N__71113),
            .I(N__71076));
    Span4Mux_v I__17363 (
            .O(N__71110),
            .I(N__71071));
    Span4Mux_h I__17362 (
            .O(N__71105),
            .I(N__71071));
    Span4Mux_h I__17361 (
            .O(N__71102),
            .I(N__71066));
    Span4Mux_h I__17360 (
            .O(N__71097),
            .I(N__71066));
    Span4Mux_h I__17359 (
            .O(N__71094),
            .I(N__71063));
    Span4Mux_v I__17358 (
            .O(N__71089),
            .I(N__71060));
    Span4Mux_v I__17357 (
            .O(N__71084),
            .I(N__71057));
    Span4Mux_h I__17356 (
            .O(N__71081),
            .I(N__71052));
    Span4Mux_h I__17355 (
            .O(N__71076),
            .I(N__71052));
    Span4Mux_h I__17354 (
            .O(N__71071),
            .I(N__71049));
    Span4Mux_h I__17353 (
            .O(N__71066),
            .I(N__71046));
    Span4Mux_h I__17352 (
            .O(N__71063),
            .I(N__71043));
    Span4Mux_h I__17351 (
            .O(N__71060),
            .I(N__71038));
    Span4Mux_h I__17350 (
            .O(N__71057),
            .I(N__71038));
    Span4Mux_h I__17349 (
            .O(N__71052),
            .I(N__71035));
    Span4Mux_h I__17348 (
            .O(N__71049),
            .I(N__71030));
    Span4Mux_v I__17347 (
            .O(N__71046),
            .I(N__71030));
    Odrv4 I__17346 (
            .O(N__71043),
            .I(\ALU.un1_a41_9_0 ));
    Odrv4 I__17345 (
            .O(N__71038),
            .I(\ALU.un1_a41_9_0 ));
    Odrv4 I__17344 (
            .O(N__71035),
            .I(\ALU.un1_a41_9_0 ));
    Odrv4 I__17343 (
            .O(N__71030),
            .I(\ALU.un1_a41_9_0 ));
    InMux I__17342 (
            .O(N__71021),
            .I(N__71012));
    InMux I__17341 (
            .O(N__71020),
            .I(N__71012));
    InMux I__17340 (
            .O(N__71019),
            .I(N__71012));
    LocalMux I__17339 (
            .O(N__71012),
            .I(\ALU.un1_a41_3_0_1 ));
    InMux I__17338 (
            .O(N__71009),
            .I(N__70997));
    InMux I__17337 (
            .O(N__71008),
            .I(N__70997));
    InMux I__17336 (
            .O(N__71007),
            .I(N__70997));
    InMux I__17335 (
            .O(N__71006),
            .I(N__70997));
    LocalMux I__17334 (
            .O(N__70997),
            .I(\ALU.un1_operation_13_0 ));
    CEMux I__17333 (
            .O(N__70994),
            .I(N__70990));
    CEMux I__17332 (
            .O(N__70993),
            .I(N__70987));
    LocalMux I__17331 (
            .O(N__70990),
            .I(N__70983));
    LocalMux I__17330 (
            .O(N__70987),
            .I(N__70980));
    CEMux I__17329 (
            .O(N__70986),
            .I(N__70977));
    Span4Mux_h I__17328 (
            .O(N__70983),
            .I(N__70974));
    Span4Mux_v I__17327 (
            .O(N__70980),
            .I(N__70971));
    LocalMux I__17326 (
            .O(N__70977),
            .I(N__70968));
    Span4Mux_h I__17325 (
            .O(N__70974),
            .I(N__70965));
    Span4Mux_v I__17324 (
            .O(N__70971),
            .I(N__70962));
    Span4Mux_h I__17323 (
            .O(N__70968),
            .I(N__70959));
    Span4Mux_h I__17322 (
            .O(N__70965),
            .I(N__70956));
    Sp12to4 I__17321 (
            .O(N__70962),
            .I(N__70953));
    Span4Mux_h I__17320 (
            .O(N__70959),
            .I(N__70948));
    Span4Mux_v I__17319 (
            .O(N__70956),
            .I(N__70948));
    Odrv12 I__17318 (
            .O(N__70953),
            .I(\ALU.un1_a41_3_0 ));
    Odrv4 I__17317 (
            .O(N__70948),
            .I(\ALU.un1_a41_3_0 ));
    CascadeMux I__17316 (
            .O(N__70943),
            .I(N__70937));
    CascadeMux I__17315 (
            .O(N__70942),
            .I(N__70932));
    InMux I__17314 (
            .O(N__70941),
            .I(N__70922));
    InMux I__17313 (
            .O(N__70940),
            .I(N__70922));
    InMux I__17312 (
            .O(N__70937),
            .I(N__70922));
    InMux I__17311 (
            .O(N__70936),
            .I(N__70922));
    InMux I__17310 (
            .O(N__70935),
            .I(N__70915));
    InMux I__17309 (
            .O(N__70932),
            .I(N__70915));
    InMux I__17308 (
            .O(N__70931),
            .I(N__70915));
    LocalMux I__17307 (
            .O(N__70922),
            .I(N__70908));
    LocalMux I__17306 (
            .O(N__70915),
            .I(N__70908));
    InMux I__17305 (
            .O(N__70914),
            .I(N__70905));
    InMux I__17304 (
            .O(N__70913),
            .I(N__70902));
    Span4Mux_v I__17303 (
            .O(N__70908),
            .I(N__70897));
    LocalMux I__17302 (
            .O(N__70905),
            .I(N__70897));
    LocalMux I__17301 (
            .O(N__70902),
            .I(aluResults_2));
    Odrv4 I__17300 (
            .O(N__70897),
            .I(aluResults_2));
    CascadeMux I__17299 (
            .O(N__70892),
            .I(N__70884));
    InMux I__17298 (
            .O(N__70891),
            .I(N__70875));
    InMux I__17297 (
            .O(N__70890),
            .I(N__70875));
    InMux I__17296 (
            .O(N__70889),
            .I(N__70875));
    InMux I__17295 (
            .O(N__70888),
            .I(N__70866));
    InMux I__17294 (
            .O(N__70887),
            .I(N__70866));
    InMux I__17293 (
            .O(N__70884),
            .I(N__70866));
    InMux I__17292 (
            .O(N__70883),
            .I(N__70866));
    InMux I__17291 (
            .O(N__70882),
            .I(N__70862));
    LocalMux I__17290 (
            .O(N__70875),
            .I(N__70859));
    LocalMux I__17289 (
            .O(N__70866),
            .I(N__70856));
    InMux I__17288 (
            .O(N__70865),
            .I(N__70853));
    LocalMux I__17287 (
            .O(N__70862),
            .I(aluResults_1));
    Odrv4 I__17286 (
            .O(N__70859),
            .I(aluResults_1));
    Odrv4 I__17285 (
            .O(N__70856),
            .I(aluResults_1));
    LocalMux I__17284 (
            .O(N__70853),
            .I(aluResults_1));
    CascadeMux I__17283 (
            .O(N__70844),
            .I(N__70841));
    InMux I__17282 (
            .O(N__70841),
            .I(N__70838));
    LocalMux I__17281 (
            .O(N__70838),
            .I(\ALU.un1_a41_2Z0Z_1 ));
    InMux I__17280 (
            .O(N__70835),
            .I(N__70832));
    LocalMux I__17279 (
            .O(N__70832),
            .I(N__70829));
    Span4Mux_v I__17278 (
            .O(N__70829),
            .I(N__70825));
    InMux I__17277 (
            .O(N__70828),
            .I(N__70822));
    Sp12to4 I__17276 (
            .O(N__70825),
            .I(N__70819));
    LocalMux I__17275 (
            .O(N__70822),
            .I(N__70816));
    Span12Mux_h I__17274 (
            .O(N__70819),
            .I(N__70812));
    Span4Mux_h I__17273 (
            .O(N__70816),
            .I(N__70809));
    InMux I__17272 (
            .O(N__70815),
            .I(N__70806));
    Odrv12 I__17271 (
            .O(N__70812),
            .I(controlWord_22));
    Odrv4 I__17270 (
            .O(N__70809),
            .I(controlWord_22));
    LocalMux I__17269 (
            .O(N__70806),
            .I(controlWord_22));
    InMux I__17268 (
            .O(N__70799),
            .I(N__70791));
    CascadeMux I__17267 (
            .O(N__70798),
            .I(N__70782));
    CascadeMux I__17266 (
            .O(N__70797),
            .I(N__70779));
    CascadeMux I__17265 (
            .O(N__70796),
            .I(N__70776));
    InMux I__17264 (
            .O(N__70795),
            .I(N__70773));
    InMux I__17263 (
            .O(N__70794),
            .I(N__70770));
    LocalMux I__17262 (
            .O(N__70791),
            .I(N__70767));
    InMux I__17261 (
            .O(N__70790),
            .I(N__70751));
    InMux I__17260 (
            .O(N__70789),
            .I(N__70746));
    InMux I__17259 (
            .O(N__70788),
            .I(N__70746));
    InMux I__17258 (
            .O(N__70787),
            .I(N__70733));
    InMux I__17257 (
            .O(N__70786),
            .I(N__70733));
    InMux I__17256 (
            .O(N__70785),
            .I(N__70733));
    InMux I__17255 (
            .O(N__70782),
            .I(N__70733));
    InMux I__17254 (
            .O(N__70779),
            .I(N__70733));
    InMux I__17253 (
            .O(N__70776),
            .I(N__70733));
    LocalMux I__17252 (
            .O(N__70773),
            .I(N__70730));
    LocalMux I__17251 (
            .O(N__70770),
            .I(N__70727));
    Span4Mux_v I__17250 (
            .O(N__70767),
            .I(N__70724));
    CascadeMux I__17249 (
            .O(N__70766),
            .I(N__70718));
    CascadeMux I__17248 (
            .O(N__70765),
            .I(N__70715));
    CascadeMux I__17247 (
            .O(N__70764),
            .I(N__70712));
    InMux I__17246 (
            .O(N__70763),
            .I(N__70703));
    InMux I__17245 (
            .O(N__70762),
            .I(N__70703));
    InMux I__17244 (
            .O(N__70761),
            .I(N__70700));
    InMux I__17243 (
            .O(N__70760),
            .I(N__70693));
    InMux I__17242 (
            .O(N__70759),
            .I(N__70693));
    InMux I__17241 (
            .O(N__70758),
            .I(N__70693));
    InMux I__17240 (
            .O(N__70757),
            .I(N__70690));
    InMux I__17239 (
            .O(N__70756),
            .I(N__70683));
    InMux I__17238 (
            .O(N__70755),
            .I(N__70683));
    InMux I__17237 (
            .O(N__70754),
            .I(N__70683));
    LocalMux I__17236 (
            .O(N__70751),
            .I(N__70678));
    LocalMux I__17235 (
            .O(N__70746),
            .I(N__70678));
    LocalMux I__17234 (
            .O(N__70733),
            .I(N__70671));
    Span4Mux_h I__17233 (
            .O(N__70730),
            .I(N__70671));
    Span4Mux_v I__17232 (
            .O(N__70727),
            .I(N__70671));
    Span4Mux_h I__17231 (
            .O(N__70724),
            .I(N__70668));
    InMux I__17230 (
            .O(N__70723),
            .I(N__70661));
    InMux I__17229 (
            .O(N__70722),
            .I(N__70661));
    InMux I__17228 (
            .O(N__70721),
            .I(N__70661));
    InMux I__17227 (
            .O(N__70718),
            .I(N__70646));
    InMux I__17226 (
            .O(N__70715),
            .I(N__70646));
    InMux I__17225 (
            .O(N__70712),
            .I(N__70646));
    InMux I__17224 (
            .O(N__70711),
            .I(N__70646));
    InMux I__17223 (
            .O(N__70710),
            .I(N__70646));
    InMux I__17222 (
            .O(N__70709),
            .I(N__70646));
    InMux I__17221 (
            .O(N__70708),
            .I(N__70646));
    LocalMux I__17220 (
            .O(N__70703),
            .I(N__70643));
    LocalMux I__17219 (
            .O(N__70700),
            .I(N__70640));
    LocalMux I__17218 (
            .O(N__70693),
            .I(N__70631));
    LocalMux I__17217 (
            .O(N__70690),
            .I(N__70631));
    LocalMux I__17216 (
            .O(N__70683),
            .I(N__70631));
    Span12Mux_h I__17215 (
            .O(N__70678),
            .I(N__70631));
    Span4Mux_h I__17214 (
            .O(N__70671),
            .I(N__70626));
    Span4Mux_h I__17213 (
            .O(N__70668),
            .I(N__70626));
    LocalMux I__17212 (
            .O(N__70661),
            .I(\CONTROL.un1_busState101_3_0_0_0 ));
    LocalMux I__17211 (
            .O(N__70646),
            .I(\CONTROL.un1_busState101_3_0_0_0 ));
    Odrv4 I__17210 (
            .O(N__70643),
            .I(\CONTROL.un1_busState101_3_0_0_0 ));
    Odrv12 I__17209 (
            .O(N__70640),
            .I(\CONTROL.un1_busState101_3_0_0_0 ));
    Odrv12 I__17208 (
            .O(N__70631),
            .I(\CONTROL.un1_busState101_3_0_0_0 ));
    Odrv4 I__17207 (
            .O(N__70626),
            .I(\CONTROL.un1_busState101_3_0_0_0 ));
    CascadeMux I__17206 (
            .O(N__70613),
            .I(N__70610));
    InMux I__17205 (
            .O(N__70610),
            .I(N__70607));
    LocalMux I__17204 (
            .O(N__70607),
            .I(N__70604));
    Span4Mux_v I__17203 (
            .O(N__70604),
            .I(N__70600));
    InMux I__17202 (
            .O(N__70603),
            .I(N__70597));
    Span4Mux_h I__17201 (
            .O(N__70600),
            .I(N__70594));
    LocalMux I__17200 (
            .O(N__70597),
            .I(N__70591));
    Span4Mux_h I__17199 (
            .O(N__70594),
            .I(N__70586));
    Span4Mux_h I__17198 (
            .O(N__70591),
            .I(N__70586));
    Span4Mux_v I__17197 (
            .O(N__70586),
            .I(N__70582));
    InMux I__17196 (
            .O(N__70585),
            .I(N__70579));
    Span4Mux_v I__17195 (
            .O(N__70582),
            .I(N__70576));
    LocalMux I__17194 (
            .O(N__70579),
            .I(N__70573));
    Sp12to4 I__17193 (
            .O(N__70576),
            .I(N__70570));
    Span4Mux_h I__17192 (
            .O(N__70573),
            .I(N__70567));
    Span12Mux_s8_v I__17191 (
            .O(N__70570),
            .I(N__70564));
    Span4Mux_h I__17190 (
            .O(N__70567),
            .I(N__70561));
    Odrv12 I__17189 (
            .O(N__70564),
            .I(f_6));
    Odrv4 I__17188 (
            .O(N__70561),
            .I(f_6));
    InMux I__17187 (
            .O(N__70556),
            .I(N__70553));
    LocalMux I__17186 (
            .O(N__70553),
            .I(N__70545));
    InMux I__17185 (
            .O(N__70552),
            .I(N__70536));
    InMux I__17184 (
            .O(N__70551),
            .I(N__70528));
    InMux I__17183 (
            .O(N__70550),
            .I(N__70528));
    InMux I__17182 (
            .O(N__70549),
            .I(N__70528));
    InMux I__17181 (
            .O(N__70548),
            .I(N__70518));
    Span4Mux_h I__17180 (
            .O(N__70545),
            .I(N__70515));
    CascadeMux I__17179 (
            .O(N__70544),
            .I(N__70511));
    InMux I__17178 (
            .O(N__70543),
            .I(N__70500));
    InMux I__17177 (
            .O(N__70542),
            .I(N__70500));
    InMux I__17176 (
            .O(N__70541),
            .I(N__70500));
    InMux I__17175 (
            .O(N__70540),
            .I(N__70500));
    InMux I__17174 (
            .O(N__70539),
            .I(N__70500));
    LocalMux I__17173 (
            .O(N__70536),
            .I(N__70497));
    InMux I__17172 (
            .O(N__70535),
            .I(N__70494));
    LocalMux I__17171 (
            .O(N__70528),
            .I(N__70491));
    InMux I__17170 (
            .O(N__70527),
            .I(N__70478));
    InMux I__17169 (
            .O(N__70526),
            .I(N__70478));
    InMux I__17168 (
            .O(N__70525),
            .I(N__70478));
    InMux I__17167 (
            .O(N__70524),
            .I(N__70478));
    InMux I__17166 (
            .O(N__70523),
            .I(N__70478));
    InMux I__17165 (
            .O(N__70522),
            .I(N__70478));
    InMux I__17164 (
            .O(N__70521),
            .I(N__70475));
    LocalMux I__17163 (
            .O(N__70518),
            .I(N__70472));
    Span4Mux_h I__17162 (
            .O(N__70515),
            .I(N__70469));
    InMux I__17161 (
            .O(N__70514),
            .I(N__70463));
    InMux I__17160 (
            .O(N__70511),
            .I(N__70452));
    LocalMux I__17159 (
            .O(N__70500),
            .I(N__70445));
    Span4Mux_h I__17158 (
            .O(N__70497),
            .I(N__70445));
    LocalMux I__17157 (
            .O(N__70494),
            .I(N__70445));
    Span4Mux_h I__17156 (
            .O(N__70491),
            .I(N__70442));
    LocalMux I__17155 (
            .O(N__70478),
            .I(N__70437));
    LocalMux I__17154 (
            .O(N__70475),
            .I(N__70437));
    Span4Mux_h I__17153 (
            .O(N__70472),
            .I(N__70432));
    Span4Mux_h I__17152 (
            .O(N__70469),
            .I(N__70432));
    InMux I__17151 (
            .O(N__70468),
            .I(N__70425));
    InMux I__17150 (
            .O(N__70467),
            .I(N__70425));
    InMux I__17149 (
            .O(N__70466),
            .I(N__70425));
    LocalMux I__17148 (
            .O(N__70463),
            .I(N__70422));
    InMux I__17147 (
            .O(N__70462),
            .I(N__70417));
    InMux I__17146 (
            .O(N__70461),
            .I(N__70417));
    InMux I__17145 (
            .O(N__70460),
            .I(N__70404));
    InMux I__17144 (
            .O(N__70459),
            .I(N__70404));
    InMux I__17143 (
            .O(N__70458),
            .I(N__70404));
    InMux I__17142 (
            .O(N__70457),
            .I(N__70404));
    InMux I__17141 (
            .O(N__70456),
            .I(N__70404));
    InMux I__17140 (
            .O(N__70455),
            .I(N__70404));
    LocalMux I__17139 (
            .O(N__70452),
            .I(N__70401));
    Span4Mux_h I__17138 (
            .O(N__70445),
            .I(N__70398));
    Span4Mux_h I__17137 (
            .O(N__70442),
            .I(N__70395));
    Span4Mux_v I__17136 (
            .O(N__70437),
            .I(N__70390));
    Span4Mux_h I__17135 (
            .O(N__70432),
            .I(N__70390));
    LocalMux I__17134 (
            .O(N__70425),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    Odrv4 I__17133 (
            .O(N__70422),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    LocalMux I__17132 (
            .O(N__70417),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    LocalMux I__17131 (
            .O(N__70404),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    Odrv4 I__17130 (
            .O(N__70401),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    Odrv4 I__17129 (
            .O(N__70398),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    Odrv4 I__17128 (
            .O(N__70395),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    Odrv4 I__17127 (
            .O(N__70390),
            .I(\CONTROL.un1_busState101_3_0Z0Z_1 ));
    IoInMux I__17126 (
            .O(N__70373),
            .I(N__70370));
    LocalMux I__17125 (
            .O(N__70370),
            .I(N__70366));
    InMux I__17124 (
            .O(N__70369),
            .I(N__70363));
    Span4Mux_s3_h I__17123 (
            .O(N__70366),
            .I(N__70360));
    LocalMux I__17122 (
            .O(N__70363),
            .I(N__70357));
    Sp12to4 I__17121 (
            .O(N__70360),
            .I(N__70354));
    Span12Mux_v I__17120 (
            .O(N__70357),
            .I(N__70351));
    Span12Mux_v I__17119 (
            .O(N__70354),
            .I(N__70348));
    Span12Mux_h I__17118 (
            .O(N__70351),
            .I(N__70345));
    Odrv12 I__17117 (
            .O(N__70348),
            .I(A6_c));
    Odrv12 I__17116 (
            .O(N__70345),
            .I(A6_c));
    CEMux I__17115 (
            .O(N__70340),
            .I(N__70337));
    LocalMux I__17114 (
            .O(N__70337),
            .I(N__70334));
    Span4Mux_v I__17113 (
            .O(N__70334),
            .I(N__70331));
    Span4Mux_h I__17112 (
            .O(N__70331),
            .I(N__70325));
    CEMux I__17111 (
            .O(N__70330),
            .I(N__70322));
    CEMux I__17110 (
            .O(N__70329),
            .I(N__70319));
    CEMux I__17109 (
            .O(N__70328),
            .I(N__70314));
    Span4Mux_v I__17108 (
            .O(N__70325),
            .I(N__70309));
    LocalMux I__17107 (
            .O(N__70322),
            .I(N__70309));
    LocalMux I__17106 (
            .O(N__70319),
            .I(N__70306));
    CEMux I__17105 (
            .O(N__70318),
            .I(N__70303));
    CEMux I__17104 (
            .O(N__70317),
            .I(N__70300));
    LocalMux I__17103 (
            .O(N__70314),
            .I(N__70297));
    Span4Mux_h I__17102 (
            .O(N__70309),
            .I(N__70292));
    Span4Mux_v I__17101 (
            .O(N__70306),
            .I(N__70292));
    LocalMux I__17100 (
            .O(N__70303),
            .I(N__70285));
    LocalMux I__17099 (
            .O(N__70300),
            .I(N__70285));
    Span4Mux_v I__17098 (
            .O(N__70297),
            .I(N__70285));
    Span4Mux_h I__17097 (
            .O(N__70292),
            .I(N__70282));
    Span4Mux_v I__17096 (
            .O(N__70285),
            .I(N__70279));
    Sp12to4 I__17095 (
            .O(N__70282),
            .I(N__70276));
    Odrv4 I__17094 (
            .O(N__70279),
            .I(\CONTROL.N_60 ));
    Odrv12 I__17093 (
            .O(N__70276),
            .I(\CONTROL.N_60 ));
    CascadeMux I__17092 (
            .O(N__70271),
            .I(\PROM.ROMDATA.m281_cascade_ ));
    InMux I__17091 (
            .O(N__70268),
            .I(N__70265));
    LocalMux I__17090 (
            .O(N__70265),
            .I(\ALU.un1_a41_7_0_2 ));
    CascadeMux I__17089 (
            .O(N__70262),
            .I(\ALU.un1_operation_13Z0Z_2_cascade_ ));
    InMux I__17088 (
            .O(N__70259),
            .I(N__70256));
    LocalMux I__17087 (
            .O(N__70256),
            .I(\ALU.un1_a41_4_0_2 ));
    CascadeMux I__17086 (
            .O(N__70253),
            .I(\ALU.un1_a41_4_0_2_cascade_ ));
    CEMux I__17085 (
            .O(N__70250),
            .I(N__70246));
    CEMux I__17084 (
            .O(N__70249),
            .I(N__70243));
    LocalMux I__17083 (
            .O(N__70246),
            .I(N__70240));
    LocalMux I__17082 (
            .O(N__70243),
            .I(N__70236));
    Span4Mux_h I__17081 (
            .O(N__70240),
            .I(N__70233));
    CEMux I__17080 (
            .O(N__70239),
            .I(N__70230));
    Span4Mux_h I__17079 (
            .O(N__70236),
            .I(N__70227));
    Span4Mux_h I__17078 (
            .O(N__70233),
            .I(N__70224));
    LocalMux I__17077 (
            .O(N__70230),
            .I(N__70221));
    Span4Mux_h I__17076 (
            .O(N__70227),
            .I(N__70218));
    Span4Mux_v I__17075 (
            .O(N__70224),
            .I(N__70215));
    Span4Mux_v I__17074 (
            .O(N__70221),
            .I(N__70212));
    Span4Mux_v I__17073 (
            .O(N__70218),
            .I(N__70209));
    Sp12to4 I__17072 (
            .O(N__70215),
            .I(N__70206));
    Odrv4 I__17071 (
            .O(N__70212),
            .I(\ALU.un1_a41_6_0 ));
    Odrv4 I__17070 (
            .O(N__70209),
            .I(\ALU.un1_a41_6_0 ));
    Odrv12 I__17069 (
            .O(N__70206),
            .I(\ALU.un1_a41_6_0 ));
    InMux I__17068 (
            .O(N__70199),
            .I(N__70192));
    InMux I__17067 (
            .O(N__70198),
            .I(N__70192));
    InMux I__17066 (
            .O(N__70197),
            .I(N__70188));
    LocalMux I__17065 (
            .O(N__70192),
            .I(N__70181));
    InMux I__17064 (
            .O(N__70191),
            .I(N__70178));
    LocalMux I__17063 (
            .O(N__70188),
            .I(N__70175));
    InMux I__17062 (
            .O(N__70187),
            .I(N__70172));
    InMux I__17061 (
            .O(N__70186),
            .I(N__70160));
    InMux I__17060 (
            .O(N__70185),
            .I(N__70160));
    InMux I__17059 (
            .O(N__70184),
            .I(N__70160));
    Span4Mux_v I__17058 (
            .O(N__70181),
            .I(N__70154));
    LocalMux I__17057 (
            .O(N__70178),
            .I(N__70147));
    Span4Mux_v I__17056 (
            .O(N__70175),
            .I(N__70147));
    LocalMux I__17055 (
            .O(N__70172),
            .I(N__70147));
    InMux I__17054 (
            .O(N__70171),
            .I(N__70140));
    InMux I__17053 (
            .O(N__70170),
            .I(N__70140));
    InMux I__17052 (
            .O(N__70169),
            .I(N__70140));
    InMux I__17051 (
            .O(N__70168),
            .I(N__70134));
    InMux I__17050 (
            .O(N__70167),
            .I(N__70134));
    LocalMux I__17049 (
            .O(N__70160),
            .I(N__70131));
    InMux I__17048 (
            .O(N__70159),
            .I(N__70128));
    InMux I__17047 (
            .O(N__70158),
            .I(N__70123));
    InMux I__17046 (
            .O(N__70157),
            .I(N__70123));
    Span4Mux_h I__17045 (
            .O(N__70154),
            .I(N__70118));
    Span4Mux_v I__17044 (
            .O(N__70147),
            .I(N__70118));
    LocalMux I__17043 (
            .O(N__70140),
            .I(N__70114));
    InMux I__17042 (
            .O(N__70139),
            .I(N__70111));
    LocalMux I__17041 (
            .O(N__70134),
            .I(N__70106));
    Span4Mux_h I__17040 (
            .O(N__70131),
            .I(N__70106));
    LocalMux I__17039 (
            .O(N__70128),
            .I(N__70103));
    LocalMux I__17038 (
            .O(N__70123),
            .I(N__70100));
    Span4Mux_h I__17037 (
            .O(N__70118),
            .I(N__70097));
    InMux I__17036 (
            .O(N__70117),
            .I(N__70091));
    Span4Mux_v I__17035 (
            .O(N__70114),
            .I(N__70085));
    LocalMux I__17034 (
            .O(N__70111),
            .I(N__70080));
    Span4Mux_v I__17033 (
            .O(N__70106),
            .I(N__70080));
    Span4Mux_v I__17032 (
            .O(N__70103),
            .I(N__70075));
    Span4Mux_v I__17031 (
            .O(N__70100),
            .I(N__70075));
    Sp12to4 I__17030 (
            .O(N__70097),
            .I(N__70072));
    InMux I__17029 (
            .O(N__70096),
            .I(N__70065));
    InMux I__17028 (
            .O(N__70095),
            .I(N__70065));
    InMux I__17027 (
            .O(N__70094),
            .I(N__70065));
    LocalMux I__17026 (
            .O(N__70091),
            .I(N__70062));
    InMux I__17025 (
            .O(N__70090),
            .I(N__70055));
    InMux I__17024 (
            .O(N__70089),
            .I(N__70055));
    InMux I__17023 (
            .O(N__70088),
            .I(N__70055));
    Span4Mux_v I__17022 (
            .O(N__70085),
            .I(N__70047));
    Span4Mux_v I__17021 (
            .O(N__70080),
            .I(N__70047));
    Span4Mux_h I__17020 (
            .O(N__70075),
            .I(N__70047));
    Span12Mux_h I__17019 (
            .O(N__70072),
            .I(N__70042));
    LocalMux I__17018 (
            .O(N__70065),
            .I(N__70042));
    Span4Mux_h I__17017 (
            .O(N__70062),
            .I(N__70037));
    LocalMux I__17016 (
            .O(N__70055),
            .I(N__70037));
    InMux I__17015 (
            .O(N__70054),
            .I(N__70034));
    Span4Mux_h I__17014 (
            .O(N__70047),
            .I(N__70031));
    Span12Mux_v I__17013 (
            .O(N__70042),
            .I(N__70028));
    Sp12to4 I__17012 (
            .O(N__70037),
            .I(N__70025));
    LocalMux I__17011 (
            .O(N__70034),
            .I(aluOperation_2));
    Odrv4 I__17010 (
            .O(N__70031),
            .I(aluOperation_2));
    Odrv12 I__17009 (
            .O(N__70028),
            .I(aluOperation_2));
    Odrv12 I__17008 (
            .O(N__70025),
            .I(aluOperation_2));
    CascadeMux I__17007 (
            .O(N__70016),
            .I(N__70013));
    InMux I__17006 (
            .O(N__70013),
            .I(N__70008));
    CascadeMux I__17005 (
            .O(N__70012),
            .I(N__70004));
    CascadeMux I__17004 (
            .O(N__70011),
            .I(N__70001));
    LocalMux I__17003 (
            .O(N__70008),
            .I(N__69995));
    InMux I__17002 (
            .O(N__70007),
            .I(N__69992));
    InMux I__17001 (
            .O(N__70004),
            .I(N__69989));
    InMux I__17000 (
            .O(N__70001),
            .I(N__69983));
    InMux I__16999 (
            .O(N__70000),
            .I(N__69983));
    InMux I__16998 (
            .O(N__69999),
            .I(N__69978));
    InMux I__16997 (
            .O(N__69998),
            .I(N__69978));
    Span4Mux_v I__16996 (
            .O(N__69995),
            .I(N__69974));
    LocalMux I__16995 (
            .O(N__69992),
            .I(N__69969));
    LocalMux I__16994 (
            .O(N__69989),
            .I(N__69962));
    InMux I__16993 (
            .O(N__69988),
            .I(N__69959));
    LocalMux I__16992 (
            .O(N__69983),
            .I(N__69954));
    LocalMux I__16991 (
            .O(N__69978),
            .I(N__69954));
    InMux I__16990 (
            .O(N__69977),
            .I(N__69951));
    Span4Mux_h I__16989 (
            .O(N__69974),
            .I(N__69948));
    InMux I__16988 (
            .O(N__69973),
            .I(N__69945));
    InMux I__16987 (
            .O(N__69972),
            .I(N__69940));
    Span4Mux_v I__16986 (
            .O(N__69969),
            .I(N__69937));
    InMux I__16985 (
            .O(N__69968),
            .I(N__69932));
    InMux I__16984 (
            .O(N__69967),
            .I(N__69932));
    InMux I__16983 (
            .O(N__69966),
            .I(N__69929));
    CascadeMux I__16982 (
            .O(N__69965),
            .I(N__69925));
    Span4Mux_v I__16981 (
            .O(N__69962),
            .I(N__69922));
    LocalMux I__16980 (
            .O(N__69959),
            .I(N__69919));
    Span4Mux_v I__16979 (
            .O(N__69954),
            .I(N__69914));
    LocalMux I__16978 (
            .O(N__69951),
            .I(N__69914));
    Span4Mux_h I__16977 (
            .O(N__69948),
            .I(N__69909));
    LocalMux I__16976 (
            .O(N__69945),
            .I(N__69909));
    InMux I__16975 (
            .O(N__69944),
            .I(N__69904));
    InMux I__16974 (
            .O(N__69943),
            .I(N__69901));
    LocalMux I__16973 (
            .O(N__69940),
            .I(N__69898));
    Span4Mux_v I__16972 (
            .O(N__69937),
            .I(N__69891));
    LocalMux I__16971 (
            .O(N__69932),
            .I(N__69891));
    LocalMux I__16970 (
            .O(N__69929),
            .I(N__69891));
    InMux I__16969 (
            .O(N__69928),
            .I(N__69886));
    InMux I__16968 (
            .O(N__69925),
            .I(N__69886));
    Span4Mux_v I__16967 (
            .O(N__69922),
            .I(N__69882));
    Span4Mux_v I__16966 (
            .O(N__69919),
            .I(N__69879));
    Sp12to4 I__16965 (
            .O(N__69914),
            .I(N__69876));
    Span4Mux_v I__16964 (
            .O(N__69909),
            .I(N__69873));
    InMux I__16963 (
            .O(N__69908),
            .I(N__69868));
    InMux I__16962 (
            .O(N__69907),
            .I(N__69868));
    LocalMux I__16961 (
            .O(N__69904),
            .I(N__69863));
    LocalMux I__16960 (
            .O(N__69901),
            .I(N__69863));
    Span4Mux_v I__16959 (
            .O(N__69898),
            .I(N__69860));
    Span4Mux_h I__16958 (
            .O(N__69891),
            .I(N__69855));
    LocalMux I__16957 (
            .O(N__69886),
            .I(N__69855));
    CascadeMux I__16956 (
            .O(N__69885),
            .I(N__69852));
    Span4Mux_v I__16955 (
            .O(N__69882),
            .I(N__69849));
    Span4Mux_h I__16954 (
            .O(N__69879),
            .I(N__69846));
    Span12Mux_s9_v I__16953 (
            .O(N__69876),
            .I(N__69839));
    Sp12to4 I__16952 (
            .O(N__69873),
            .I(N__69839));
    LocalMux I__16951 (
            .O(N__69868),
            .I(N__69839));
    Span4Mux_v I__16950 (
            .O(N__69863),
            .I(N__69836));
    Span4Mux_h I__16949 (
            .O(N__69860),
            .I(N__69833));
    Span4Mux_h I__16948 (
            .O(N__69855),
            .I(N__69830));
    InMux I__16947 (
            .O(N__69852),
            .I(N__69827));
    Span4Mux_h I__16946 (
            .O(N__69849),
            .I(N__69822));
    Span4Mux_h I__16945 (
            .O(N__69846),
            .I(N__69822));
    Span12Mux_h I__16944 (
            .O(N__69839),
            .I(N__69819));
    Span4Mux_v I__16943 (
            .O(N__69836),
            .I(N__69812));
    Span4Mux_h I__16942 (
            .O(N__69833),
            .I(N__69812));
    Span4Mux_v I__16941 (
            .O(N__69830),
            .I(N__69812));
    LocalMux I__16940 (
            .O(N__69827),
            .I(aluOperation_4));
    Odrv4 I__16939 (
            .O(N__69822),
            .I(aluOperation_4));
    Odrv12 I__16938 (
            .O(N__69819),
            .I(aluOperation_4));
    Odrv4 I__16937 (
            .O(N__69812),
            .I(aluOperation_4));
    CascadeMux I__16936 (
            .O(N__69803),
            .I(N__69800));
    InMux I__16935 (
            .O(N__69800),
            .I(N__69791));
    InMux I__16934 (
            .O(N__69799),
            .I(N__69791));
    InMux I__16933 (
            .O(N__69798),
            .I(N__69791));
    LocalMux I__16932 (
            .O(N__69791),
            .I(N__69786));
    InMux I__16931 (
            .O(N__69790),
            .I(N__69783));
    InMux I__16930 (
            .O(N__69789),
            .I(N__69780));
    Span4Mux_h I__16929 (
            .O(N__69786),
            .I(N__69773));
    LocalMux I__16928 (
            .O(N__69783),
            .I(N__69773));
    LocalMux I__16927 (
            .O(N__69780),
            .I(N__69773));
    Span4Mux_h I__16926 (
            .O(N__69773),
            .I(N__69770));
    Span4Mux_h I__16925 (
            .O(N__69770),
            .I(N__69767));
    Span4Mux_h I__16924 (
            .O(N__69767),
            .I(N__69763));
    InMux I__16923 (
            .O(N__69766),
            .I(N__69760));
    Span4Mux_h I__16922 (
            .O(N__69763),
            .I(N__69757));
    LocalMux I__16921 (
            .O(N__69760),
            .I(aluOperation_3));
    Odrv4 I__16920 (
            .O(N__69757),
            .I(aluOperation_3));
    CascadeMux I__16919 (
            .O(N__69752),
            .I(N__69749));
    InMux I__16918 (
            .O(N__69749),
            .I(N__69739));
    InMux I__16917 (
            .O(N__69748),
            .I(N__69739));
    CascadeMux I__16916 (
            .O(N__69747),
            .I(N__69736));
    CascadeMux I__16915 (
            .O(N__69746),
            .I(N__69733));
    CascadeMux I__16914 (
            .O(N__69745),
            .I(N__69730));
    CascadeMux I__16913 (
            .O(N__69744),
            .I(N__69726));
    LocalMux I__16912 (
            .O(N__69739),
            .I(N__69723));
    InMux I__16911 (
            .O(N__69736),
            .I(N__69720));
    InMux I__16910 (
            .O(N__69733),
            .I(N__69717));
    InMux I__16909 (
            .O(N__69730),
            .I(N__69712));
    InMux I__16908 (
            .O(N__69729),
            .I(N__69707));
    InMux I__16907 (
            .O(N__69726),
            .I(N__69707));
    Span4Mux_v I__16906 (
            .O(N__69723),
            .I(N__69700));
    LocalMux I__16905 (
            .O(N__69720),
            .I(N__69700));
    LocalMux I__16904 (
            .O(N__69717),
            .I(N__69700));
    CascadeMux I__16903 (
            .O(N__69716),
            .I(N__69694));
    CascadeMux I__16902 (
            .O(N__69715),
            .I(N__69691));
    LocalMux I__16901 (
            .O(N__69712),
            .I(N__69684));
    LocalMux I__16900 (
            .O(N__69707),
            .I(N__69684));
    Span4Mux_v I__16899 (
            .O(N__69700),
            .I(N__69681));
    CascadeMux I__16898 (
            .O(N__69699),
            .I(N__69675));
    CascadeMux I__16897 (
            .O(N__69698),
            .I(N__69672));
    InMux I__16896 (
            .O(N__69697),
            .I(N__69667));
    InMux I__16895 (
            .O(N__69694),
            .I(N__69667));
    InMux I__16894 (
            .O(N__69691),
            .I(N__69661));
    InMux I__16893 (
            .O(N__69690),
            .I(N__69661));
    CascadeMux I__16892 (
            .O(N__69689),
            .I(N__69658));
    Span4Mux_v I__16891 (
            .O(N__69684),
            .I(N__69655));
    Span4Mux_v I__16890 (
            .O(N__69681),
            .I(N__69652));
    CascadeMux I__16889 (
            .O(N__69680),
            .I(N__69648));
    CascadeMux I__16888 (
            .O(N__69679),
            .I(N__69642));
    CascadeMux I__16887 (
            .O(N__69678),
            .I(N__69637));
    InMux I__16886 (
            .O(N__69675),
            .I(N__69634));
    InMux I__16885 (
            .O(N__69672),
            .I(N__69631));
    LocalMux I__16884 (
            .O(N__69667),
            .I(N__69628));
    CascadeMux I__16883 (
            .O(N__69666),
            .I(N__69624));
    LocalMux I__16882 (
            .O(N__69661),
            .I(N__69621));
    InMux I__16881 (
            .O(N__69658),
            .I(N__69618));
    Span4Mux_h I__16880 (
            .O(N__69655),
            .I(N__69613));
    Span4Mux_h I__16879 (
            .O(N__69652),
            .I(N__69613));
    InMux I__16878 (
            .O(N__69651),
            .I(N__69610));
    InMux I__16877 (
            .O(N__69648),
            .I(N__69603));
    InMux I__16876 (
            .O(N__69647),
            .I(N__69603));
    InMux I__16875 (
            .O(N__69646),
            .I(N__69603));
    InMux I__16874 (
            .O(N__69645),
            .I(N__69596));
    InMux I__16873 (
            .O(N__69642),
            .I(N__69596));
    InMux I__16872 (
            .O(N__69641),
            .I(N__69596));
    InMux I__16871 (
            .O(N__69640),
            .I(N__69593));
    InMux I__16870 (
            .O(N__69637),
            .I(N__69590));
    LocalMux I__16869 (
            .O(N__69634),
            .I(N__69583));
    LocalMux I__16868 (
            .O(N__69631),
            .I(N__69583));
    Span4Mux_h I__16867 (
            .O(N__69628),
            .I(N__69583));
    InMux I__16866 (
            .O(N__69627),
            .I(N__69580));
    InMux I__16865 (
            .O(N__69624),
            .I(N__69577));
    Span4Mux_v I__16864 (
            .O(N__69621),
            .I(N__69574));
    LocalMux I__16863 (
            .O(N__69618),
            .I(N__69563));
    Span4Mux_v I__16862 (
            .O(N__69613),
            .I(N__69563));
    LocalMux I__16861 (
            .O(N__69610),
            .I(N__69563));
    LocalMux I__16860 (
            .O(N__69603),
            .I(N__69563));
    LocalMux I__16859 (
            .O(N__69596),
            .I(N__69563));
    LocalMux I__16858 (
            .O(N__69593),
            .I(N__69560));
    LocalMux I__16857 (
            .O(N__69590),
            .I(N__69555));
    Span4Mux_h I__16856 (
            .O(N__69583),
            .I(N__69555));
    LocalMux I__16855 (
            .O(N__69580),
            .I(N__69552));
    LocalMux I__16854 (
            .O(N__69577),
            .I(N__69547));
    Span4Mux_h I__16853 (
            .O(N__69574),
            .I(N__69547));
    Span4Mux_v I__16852 (
            .O(N__69563),
            .I(N__69544));
    Span4Mux_h I__16851 (
            .O(N__69560),
            .I(N__69539));
    Span4Mux_v I__16850 (
            .O(N__69555),
            .I(N__69539));
    Odrv12 I__16849 (
            .O(N__69552),
            .I(\ALU.a32Z0Z_0 ));
    Odrv4 I__16848 (
            .O(N__69547),
            .I(\ALU.a32Z0Z_0 ));
    Odrv4 I__16847 (
            .O(N__69544),
            .I(\ALU.a32Z0Z_0 ));
    Odrv4 I__16846 (
            .O(N__69539),
            .I(\ALU.a32Z0Z_0 ));
    InMux I__16845 (
            .O(N__69530),
            .I(N__69526));
    InMux I__16844 (
            .O(N__69529),
            .I(N__69523));
    LocalMux I__16843 (
            .O(N__69526),
            .I(N__69520));
    LocalMux I__16842 (
            .O(N__69523),
            .I(N__69514));
    Sp12to4 I__16841 (
            .O(N__69520),
            .I(N__69514));
    InMux I__16840 (
            .O(N__69519),
            .I(N__69509));
    Span12Mux_v I__16839 (
            .O(N__69514),
            .I(N__69506));
    InMux I__16838 (
            .O(N__69513),
            .I(N__69503));
    InMux I__16837 (
            .O(N__69512),
            .I(N__69500));
    LocalMux I__16836 (
            .O(N__69509),
            .I(N__69497));
    Span12Mux_h I__16835 (
            .O(N__69506),
            .I(N__69493));
    LocalMux I__16834 (
            .O(N__69503),
            .I(N__69490));
    LocalMux I__16833 (
            .O(N__69500),
            .I(N__69487));
    Span4Mux_h I__16832 (
            .O(N__69497),
            .I(N__69484));
    CascadeMux I__16831 (
            .O(N__69496),
            .I(N__69481));
    Span12Mux_v I__16830 (
            .O(N__69493),
            .I(N__69478));
    Span4Mux_v I__16829 (
            .O(N__69490),
            .I(N__69473));
    Span4Mux_h I__16828 (
            .O(N__69487),
            .I(N__69473));
    Span4Mux_h I__16827 (
            .O(N__69484),
            .I(N__69470));
    InMux I__16826 (
            .O(N__69481),
            .I(N__69467));
    Odrv12 I__16825 (
            .O(N__69478),
            .I(\ALU.un1_operationZ0Z_7 ));
    Odrv4 I__16824 (
            .O(N__69473),
            .I(\ALU.un1_operationZ0Z_7 ));
    Odrv4 I__16823 (
            .O(N__69470),
            .I(\ALU.un1_operationZ0Z_7 ));
    LocalMux I__16822 (
            .O(N__69467),
            .I(\ALU.un1_operationZ0Z_7 ));
    CEMux I__16821 (
            .O(N__69458),
            .I(N__69455));
    LocalMux I__16820 (
            .O(N__69455),
            .I(N__69446));
    CEMux I__16819 (
            .O(N__69454),
            .I(N__69443));
    CEMux I__16818 (
            .O(N__69453),
            .I(N__69440));
    CEMux I__16817 (
            .O(N__69452),
            .I(N__69437));
    CEMux I__16816 (
            .O(N__69451),
            .I(N__69434));
    CEMux I__16815 (
            .O(N__69450),
            .I(N__69431));
    CEMux I__16814 (
            .O(N__69449),
            .I(N__69428));
    Span4Mux_v I__16813 (
            .O(N__69446),
            .I(N__69425));
    LocalMux I__16812 (
            .O(N__69443),
            .I(N__69422));
    LocalMux I__16811 (
            .O(N__69440),
            .I(N__69419));
    LocalMux I__16810 (
            .O(N__69437),
            .I(N__69416));
    LocalMux I__16809 (
            .O(N__69434),
            .I(N__69413));
    LocalMux I__16808 (
            .O(N__69431),
            .I(N__69408));
    LocalMux I__16807 (
            .O(N__69428),
            .I(N__69408));
    Span4Mux_v I__16806 (
            .O(N__69425),
            .I(N__69405));
    Span4Mux_h I__16805 (
            .O(N__69422),
            .I(N__69402));
    Span4Mux_h I__16804 (
            .O(N__69419),
            .I(N__69399));
    Span4Mux_h I__16803 (
            .O(N__69416),
            .I(N__69396));
    Span4Mux_h I__16802 (
            .O(N__69413),
            .I(N__69393));
    Span4Mux_h I__16801 (
            .O(N__69408),
            .I(N__69390));
    Sp12to4 I__16800 (
            .O(N__69405),
            .I(N__69387));
    Span4Mux_h I__16799 (
            .O(N__69402),
            .I(N__69382));
    Span4Mux_h I__16798 (
            .O(N__69399),
            .I(N__69382));
    Span4Mux_h I__16797 (
            .O(N__69396),
            .I(N__69379));
    Span4Mux_h I__16796 (
            .O(N__69393),
            .I(N__69376));
    Sp12to4 I__16795 (
            .O(N__69390),
            .I(N__69373));
    Span12Mux_h I__16794 (
            .O(N__69387),
            .I(N__69370));
    Odrv4 I__16793 (
            .O(N__69382),
            .I(\ALU.un1_a41_2_0 ));
    Odrv4 I__16792 (
            .O(N__69379),
            .I(\ALU.un1_a41_2_0 ));
    Odrv4 I__16791 (
            .O(N__69376),
            .I(\ALU.un1_a41_2_0 ));
    Odrv12 I__16790 (
            .O(N__69373),
            .I(\ALU.un1_a41_2_0 ));
    Odrv12 I__16789 (
            .O(N__69370),
            .I(\ALU.un1_a41_2_0 ));
    CascadeMux I__16788 (
            .O(N__69359),
            .I(N__69356));
    InMux I__16787 (
            .O(N__69356),
            .I(N__69353));
    LocalMux I__16786 (
            .O(N__69353),
            .I(N__69350));
    Span4Mux_h I__16785 (
            .O(N__69350),
            .I(N__69347));
    Span4Mux_h I__16784 (
            .O(N__69347),
            .I(N__69344));
    Span4Mux_v I__16783 (
            .O(N__69344),
            .I(N__69341));
    Odrv4 I__16782 (
            .O(N__69341),
            .I(\PROM.ROMDATA.m160 ));
    CascadeMux I__16781 (
            .O(N__69338),
            .I(N__69334));
    InMux I__16780 (
            .O(N__69337),
            .I(N__69324));
    InMux I__16779 (
            .O(N__69334),
            .I(N__69324));
    InMux I__16778 (
            .O(N__69333),
            .I(N__69324));
    InMux I__16777 (
            .O(N__69332),
            .I(N__69319));
    InMux I__16776 (
            .O(N__69331),
            .I(N__69319));
    LocalMux I__16775 (
            .O(N__69324),
            .I(N__69312));
    LocalMux I__16774 (
            .O(N__69319),
            .I(N__69312));
    InMux I__16773 (
            .O(N__69318),
            .I(N__69309));
    InMux I__16772 (
            .O(N__69317),
            .I(N__69306));
    Span4Mux_v I__16771 (
            .O(N__69312),
            .I(N__69303));
    LocalMux I__16770 (
            .O(N__69309),
            .I(N__69298));
    LocalMux I__16769 (
            .O(N__69306),
            .I(N__69298));
    Span4Mux_h I__16768 (
            .O(N__69303),
            .I(N__69295));
    Span12Mux_v I__16767 (
            .O(N__69298),
            .I(N__69292));
    Span4Mux_h I__16766 (
            .O(N__69295),
            .I(N__69289));
    Odrv12 I__16765 (
            .O(N__69292),
            .I(aluOperation_6));
    Odrv4 I__16764 (
            .O(N__69289),
            .I(aluOperation_6));
    InMux I__16763 (
            .O(N__69284),
            .I(N__69276));
    InMux I__16762 (
            .O(N__69283),
            .I(N__69276));
    InMux I__16761 (
            .O(N__69282),
            .I(N__69271));
    InMux I__16760 (
            .O(N__69281),
            .I(N__69271));
    LocalMux I__16759 (
            .O(N__69276),
            .I(N__69267));
    LocalMux I__16758 (
            .O(N__69271),
            .I(N__69264));
    InMux I__16757 (
            .O(N__69270),
            .I(N__69261));
    Span4Mux_v I__16756 (
            .O(N__69267),
            .I(N__69258));
    Span4Mux_h I__16755 (
            .O(N__69264),
            .I(N__69255));
    LocalMux I__16754 (
            .O(N__69261),
            .I(aluResults_0));
    Odrv4 I__16753 (
            .O(N__69258),
            .I(aluResults_0));
    Odrv4 I__16752 (
            .O(N__69255),
            .I(aluResults_0));
    CascadeMux I__16751 (
            .O(N__69248),
            .I(\ALU.un1_a41_3_0_1_cascade_ ));
    CEMux I__16750 (
            .O(N__69245),
            .I(N__69240));
    CEMux I__16749 (
            .O(N__69244),
            .I(N__69237));
    CEMux I__16748 (
            .O(N__69243),
            .I(N__69234));
    LocalMux I__16747 (
            .O(N__69240),
            .I(N__69231));
    LocalMux I__16746 (
            .O(N__69237),
            .I(N__69228));
    LocalMux I__16745 (
            .O(N__69234),
            .I(N__69225));
    Span4Mux_h I__16744 (
            .O(N__69231),
            .I(N__69222));
    Span4Mux_v I__16743 (
            .O(N__69228),
            .I(N__69219));
    Span4Mux_v I__16742 (
            .O(N__69225),
            .I(N__69216));
    Span4Mux_v I__16741 (
            .O(N__69222),
            .I(N__69213));
    Span4Mux_h I__16740 (
            .O(N__69219),
            .I(N__69210));
    Span4Mux_h I__16739 (
            .O(N__69216),
            .I(N__69207));
    Span4Mux_h I__16738 (
            .O(N__69213),
            .I(N__69204));
    Span4Mux_h I__16737 (
            .O(N__69210),
            .I(N__69201));
    Span4Mux_h I__16736 (
            .O(N__69207),
            .I(N__69198));
    Span4Mux_h I__16735 (
            .O(N__69204),
            .I(N__69195));
    Odrv4 I__16734 (
            .O(N__69201),
            .I(\ALU.un1_a41_5_0 ));
    Odrv4 I__16733 (
            .O(N__69198),
            .I(\ALU.un1_a41_5_0 ));
    Odrv4 I__16732 (
            .O(N__69195),
            .I(\ALU.un1_a41_5_0 ));
    InMux I__16731 (
            .O(N__69188),
            .I(N__69185));
    LocalMux I__16730 (
            .O(N__69185),
            .I(N__69182));
    Span4Mux_v I__16729 (
            .O(N__69182),
            .I(N__69179));
    Odrv4 I__16728 (
            .O(N__69179),
            .I(\ALU.N_863 ));
    CascadeMux I__16727 (
            .O(N__69176),
            .I(\ALU.N_859_cascade_ ));
    CascadeMux I__16726 (
            .O(N__69173),
            .I(\ALU.rshift_15_ns_1_1_cascade_ ));
    InMux I__16725 (
            .O(N__69170),
            .I(N__69165));
    InMux I__16724 (
            .O(N__69169),
            .I(N__69162));
    CascadeMux I__16723 (
            .O(N__69168),
            .I(N__69157));
    LocalMux I__16722 (
            .O(N__69165),
            .I(N__69151));
    LocalMux I__16721 (
            .O(N__69162),
            .I(N__69151));
    InMux I__16720 (
            .O(N__69161),
            .I(N__69146));
    InMux I__16719 (
            .O(N__69160),
            .I(N__69143));
    InMux I__16718 (
            .O(N__69157),
            .I(N__69140));
    InMux I__16717 (
            .O(N__69156),
            .I(N__69137));
    Span4Mux_v I__16716 (
            .O(N__69151),
            .I(N__69134));
    InMux I__16715 (
            .O(N__69150),
            .I(N__69131));
    InMux I__16714 (
            .O(N__69149),
            .I(N__69128));
    LocalMux I__16713 (
            .O(N__69146),
            .I(N__69121));
    LocalMux I__16712 (
            .O(N__69143),
            .I(N__69121));
    LocalMux I__16711 (
            .O(N__69140),
            .I(N__69121));
    LocalMux I__16710 (
            .O(N__69137),
            .I(N__69118));
    Span4Mux_h I__16709 (
            .O(N__69134),
            .I(N__69112));
    LocalMux I__16708 (
            .O(N__69131),
            .I(N__69112));
    LocalMux I__16707 (
            .O(N__69128),
            .I(N__69107));
    Span4Mux_v I__16706 (
            .O(N__69121),
            .I(N__69107));
    Span4Mux_v I__16705 (
            .O(N__69118),
            .I(N__69103));
    InMux I__16704 (
            .O(N__69117),
            .I(N__69100));
    Span4Mux_v I__16703 (
            .O(N__69112),
            .I(N__69095));
    Span4Mux_h I__16702 (
            .O(N__69107),
            .I(N__69095));
    InMux I__16701 (
            .O(N__69106),
            .I(N__69092));
    Span4Mux_h I__16700 (
            .O(N__69103),
            .I(N__69089));
    LocalMux I__16699 (
            .O(N__69100),
            .I(N__69084));
    Span4Mux_h I__16698 (
            .O(N__69095),
            .I(N__69084));
    LocalMux I__16697 (
            .O(N__69092),
            .I(\ALU.a_15_m2_sZ0Z_1 ));
    Odrv4 I__16696 (
            .O(N__69089),
            .I(\ALU.a_15_m2_sZ0Z_1 ));
    Odrv4 I__16695 (
            .O(N__69084),
            .I(\ALU.a_15_m2_sZ0Z_1 ));
    CascadeMux I__16694 (
            .O(N__69077),
            .I(\ALU.rshift_1_cascade_ ));
    IoInMux I__16693 (
            .O(N__69074),
            .I(N__69071));
    LocalMux I__16692 (
            .O(N__69071),
            .I(N__69067));
    IoInMux I__16691 (
            .O(N__69070),
            .I(N__69064));
    IoSpan4Mux I__16690 (
            .O(N__69067),
            .I(N__69061));
    LocalMux I__16689 (
            .O(N__69064),
            .I(N__69058));
    IoSpan4Mux I__16688 (
            .O(N__69061),
            .I(N__69054));
    IoSpan4Mux I__16687 (
            .O(N__69058),
            .I(N__69051));
    InMux I__16686 (
            .O(N__69057),
            .I(N__69048));
    Sp12to4 I__16685 (
            .O(N__69054),
            .I(N__69045));
    Span4Mux_s2_h I__16684 (
            .O(N__69051),
            .I(N__69042));
    LocalMux I__16683 (
            .O(N__69048),
            .I(N__69039));
    Span12Mux_s7_h I__16682 (
            .O(N__69045),
            .I(N__69036));
    Sp12to4 I__16681 (
            .O(N__69042),
            .I(N__69033));
    Span4Mux_v I__16680 (
            .O(N__69039),
            .I(N__69030));
    Span12Mux_h I__16679 (
            .O(N__69036),
            .I(N__69027));
    Span12Mux_v I__16678 (
            .O(N__69033),
            .I(N__69024));
    Sp12to4 I__16677 (
            .O(N__69030),
            .I(N__69021));
    Odrv12 I__16676 (
            .O(N__69027),
            .I(bus_1));
    Odrv12 I__16675 (
            .O(N__69024),
            .I(bus_1));
    Odrv12 I__16674 (
            .O(N__69021),
            .I(bus_1));
    InMux I__16673 (
            .O(N__69014),
            .I(N__69006));
    InMux I__16672 (
            .O(N__69013),
            .I(N__69003));
    InMux I__16671 (
            .O(N__69012),
            .I(N__68999));
    InMux I__16670 (
            .O(N__69011),
            .I(N__68996));
    InMux I__16669 (
            .O(N__69010),
            .I(N__68993));
    InMux I__16668 (
            .O(N__69009),
            .I(N__68990));
    LocalMux I__16667 (
            .O(N__69006),
            .I(N__68986));
    LocalMux I__16666 (
            .O(N__69003),
            .I(N__68983));
    InMux I__16665 (
            .O(N__69002),
            .I(N__68980));
    LocalMux I__16664 (
            .O(N__68999),
            .I(N__68977));
    LocalMux I__16663 (
            .O(N__68996),
            .I(N__68970));
    LocalMux I__16662 (
            .O(N__68993),
            .I(N__68970));
    LocalMux I__16661 (
            .O(N__68990),
            .I(N__68970));
    InMux I__16660 (
            .O(N__68989),
            .I(N__68967));
    Span4Mux_v I__16659 (
            .O(N__68986),
            .I(N__68962));
    Span4Mux_v I__16658 (
            .O(N__68983),
            .I(N__68962));
    LocalMux I__16657 (
            .O(N__68980),
            .I(N__68955));
    Span4Mux_v I__16656 (
            .O(N__68977),
            .I(N__68955));
    Span4Mux_v I__16655 (
            .O(N__68970),
            .I(N__68955));
    LocalMux I__16654 (
            .O(N__68967),
            .I(N__68950));
    Span4Mux_h I__16653 (
            .O(N__68962),
            .I(N__68950));
    Odrv4 I__16652 (
            .O(N__68955),
            .I(\ALU.c_RNI98D92DZ0Z_15 ));
    Odrv4 I__16651 (
            .O(N__68950),
            .I(\ALU.c_RNI98D92DZ0Z_15 ));
    InMux I__16650 (
            .O(N__68945),
            .I(N__68936));
    InMux I__16649 (
            .O(N__68944),
            .I(N__68914));
    InMux I__16648 (
            .O(N__68943),
            .I(N__68911));
    InMux I__16647 (
            .O(N__68942),
            .I(N__68901));
    InMux I__16646 (
            .O(N__68941),
            .I(N__68901));
    InMux I__16645 (
            .O(N__68940),
            .I(N__68901));
    InMux I__16644 (
            .O(N__68939),
            .I(N__68898));
    LocalMux I__16643 (
            .O(N__68936),
            .I(N__68891));
    InMux I__16642 (
            .O(N__68935),
            .I(N__68886));
    InMux I__16641 (
            .O(N__68934),
            .I(N__68886));
    InMux I__16640 (
            .O(N__68933),
            .I(N__68883));
    CascadeMux I__16639 (
            .O(N__68932),
            .I(N__68880));
    InMux I__16638 (
            .O(N__68931),
            .I(N__68875));
    InMux I__16637 (
            .O(N__68930),
            .I(N__68875));
    InMux I__16636 (
            .O(N__68929),
            .I(N__68872));
    InMux I__16635 (
            .O(N__68928),
            .I(N__68867));
    InMux I__16634 (
            .O(N__68927),
            .I(N__68867));
    InMux I__16633 (
            .O(N__68926),
            .I(N__68860));
    InMux I__16632 (
            .O(N__68925),
            .I(N__68860));
    InMux I__16631 (
            .O(N__68924),
            .I(N__68860));
    InMux I__16630 (
            .O(N__68923),
            .I(N__68855));
    InMux I__16629 (
            .O(N__68922),
            .I(N__68855));
    InMux I__16628 (
            .O(N__68921),
            .I(N__68852));
    InMux I__16627 (
            .O(N__68920),
            .I(N__68847));
    InMux I__16626 (
            .O(N__68919),
            .I(N__68847));
    InMux I__16625 (
            .O(N__68918),
            .I(N__68836));
    InMux I__16624 (
            .O(N__68917),
            .I(N__68836));
    LocalMux I__16623 (
            .O(N__68914),
            .I(N__68831));
    LocalMux I__16622 (
            .O(N__68911),
            .I(N__68831));
    InMux I__16621 (
            .O(N__68910),
            .I(N__68826));
    InMux I__16620 (
            .O(N__68909),
            .I(N__68826));
    CascadeMux I__16619 (
            .O(N__68908),
            .I(N__68819));
    LocalMux I__16618 (
            .O(N__68901),
            .I(N__68816));
    LocalMux I__16617 (
            .O(N__68898),
            .I(N__68813));
    InMux I__16616 (
            .O(N__68897),
            .I(N__68804));
    InMux I__16615 (
            .O(N__68896),
            .I(N__68804));
    InMux I__16614 (
            .O(N__68895),
            .I(N__68799));
    InMux I__16613 (
            .O(N__68894),
            .I(N__68799));
    Span4Mux_v I__16612 (
            .O(N__68891),
            .I(N__68796));
    LocalMux I__16611 (
            .O(N__68886),
            .I(N__68791));
    LocalMux I__16610 (
            .O(N__68883),
            .I(N__68791));
    InMux I__16609 (
            .O(N__68880),
            .I(N__68786));
    LocalMux I__16608 (
            .O(N__68875),
            .I(N__68783));
    LocalMux I__16607 (
            .O(N__68872),
            .I(N__68774));
    LocalMux I__16606 (
            .O(N__68867),
            .I(N__68774));
    LocalMux I__16605 (
            .O(N__68860),
            .I(N__68774));
    LocalMux I__16604 (
            .O(N__68855),
            .I(N__68774));
    LocalMux I__16603 (
            .O(N__68852),
            .I(N__68769));
    LocalMux I__16602 (
            .O(N__68847),
            .I(N__68769));
    InMux I__16601 (
            .O(N__68846),
            .I(N__68762));
    InMux I__16600 (
            .O(N__68845),
            .I(N__68762));
    InMux I__16599 (
            .O(N__68844),
            .I(N__68762));
    InMux I__16598 (
            .O(N__68843),
            .I(N__68755));
    InMux I__16597 (
            .O(N__68842),
            .I(N__68755));
    InMux I__16596 (
            .O(N__68841),
            .I(N__68755));
    LocalMux I__16595 (
            .O(N__68836),
            .I(N__68752));
    Span4Mux_h I__16594 (
            .O(N__68831),
            .I(N__68747));
    LocalMux I__16593 (
            .O(N__68826),
            .I(N__68747));
    InMux I__16592 (
            .O(N__68825),
            .I(N__68741));
    InMux I__16591 (
            .O(N__68824),
            .I(N__68734));
    InMux I__16590 (
            .O(N__68823),
            .I(N__68734));
    InMux I__16589 (
            .O(N__68822),
            .I(N__68734));
    InMux I__16588 (
            .O(N__68819),
            .I(N__68730));
    Span4Mux_v I__16587 (
            .O(N__68816),
            .I(N__68722));
    Span4Mux_h I__16586 (
            .O(N__68813),
            .I(N__68722));
    InMux I__16585 (
            .O(N__68812),
            .I(N__68712));
    InMux I__16584 (
            .O(N__68811),
            .I(N__68712));
    InMux I__16583 (
            .O(N__68810),
            .I(N__68712));
    InMux I__16582 (
            .O(N__68809),
            .I(N__68709));
    LocalMux I__16581 (
            .O(N__68804),
            .I(N__68706));
    LocalMux I__16580 (
            .O(N__68799),
            .I(N__68703));
    Span4Mux_v I__16579 (
            .O(N__68796),
            .I(N__68698));
    Span4Mux_v I__16578 (
            .O(N__68791),
            .I(N__68698));
    InMux I__16577 (
            .O(N__68790),
            .I(N__68693));
    InMux I__16576 (
            .O(N__68789),
            .I(N__68693));
    LocalMux I__16575 (
            .O(N__68786),
            .I(N__68690));
    Span4Mux_v I__16574 (
            .O(N__68783),
            .I(N__68679));
    Span4Mux_h I__16573 (
            .O(N__68774),
            .I(N__68679));
    Span4Mux_v I__16572 (
            .O(N__68769),
            .I(N__68679));
    LocalMux I__16571 (
            .O(N__68762),
            .I(N__68679));
    LocalMux I__16570 (
            .O(N__68755),
            .I(N__68679));
    Span4Mux_h I__16569 (
            .O(N__68752),
            .I(N__68674));
    Span4Mux_h I__16568 (
            .O(N__68747),
            .I(N__68674));
    InMux I__16567 (
            .O(N__68746),
            .I(N__68667));
    InMux I__16566 (
            .O(N__68745),
            .I(N__68667));
    InMux I__16565 (
            .O(N__68744),
            .I(N__68667));
    LocalMux I__16564 (
            .O(N__68741),
            .I(N__68662));
    LocalMux I__16563 (
            .O(N__68734),
            .I(N__68662));
    CascadeMux I__16562 (
            .O(N__68733),
            .I(N__68655));
    LocalMux I__16561 (
            .O(N__68730),
            .I(N__68652));
    InMux I__16560 (
            .O(N__68729),
            .I(N__68649));
    InMux I__16559 (
            .O(N__68728),
            .I(N__68646));
    InMux I__16558 (
            .O(N__68727),
            .I(N__68643));
    Span4Mux_v I__16557 (
            .O(N__68722),
            .I(N__68640));
    InMux I__16556 (
            .O(N__68721),
            .I(N__68637));
    InMux I__16555 (
            .O(N__68720),
            .I(N__68632));
    InMux I__16554 (
            .O(N__68719),
            .I(N__68632));
    LocalMux I__16553 (
            .O(N__68712),
            .I(N__68619));
    LocalMux I__16552 (
            .O(N__68709),
            .I(N__68619));
    Span12Mux_s11_h I__16551 (
            .O(N__68706),
            .I(N__68619));
    Span12Mux_v I__16550 (
            .O(N__68703),
            .I(N__68619));
    Sp12to4 I__16549 (
            .O(N__68698),
            .I(N__68619));
    LocalMux I__16548 (
            .O(N__68693),
            .I(N__68619));
    Span4Mux_v I__16547 (
            .O(N__68690),
            .I(N__68614));
    Span4Mux_h I__16546 (
            .O(N__68679),
            .I(N__68614));
    Span4Mux_h I__16545 (
            .O(N__68674),
            .I(N__68607));
    LocalMux I__16544 (
            .O(N__68667),
            .I(N__68607));
    Span4Mux_h I__16543 (
            .O(N__68662),
            .I(N__68607));
    InMux I__16542 (
            .O(N__68661),
            .I(N__68600));
    InMux I__16541 (
            .O(N__68660),
            .I(N__68600));
    InMux I__16540 (
            .O(N__68659),
            .I(N__68600));
    InMux I__16539 (
            .O(N__68658),
            .I(N__68595));
    InMux I__16538 (
            .O(N__68655),
            .I(N__68595));
    Span4Mux_h I__16537 (
            .O(N__68652),
            .I(N__68588));
    LocalMux I__16536 (
            .O(N__68649),
            .I(N__68588));
    LocalMux I__16535 (
            .O(N__68646),
            .I(N__68588));
    LocalMux I__16534 (
            .O(N__68643),
            .I(\ALU.status_19_1 ));
    Odrv4 I__16533 (
            .O(N__68640),
            .I(\ALU.status_19_1 ));
    LocalMux I__16532 (
            .O(N__68637),
            .I(\ALU.status_19_1 ));
    LocalMux I__16531 (
            .O(N__68632),
            .I(\ALU.status_19_1 ));
    Odrv12 I__16530 (
            .O(N__68619),
            .I(\ALU.status_19_1 ));
    Odrv4 I__16529 (
            .O(N__68614),
            .I(\ALU.status_19_1 ));
    Odrv4 I__16528 (
            .O(N__68607),
            .I(\ALU.status_19_1 ));
    LocalMux I__16527 (
            .O(N__68600),
            .I(\ALU.status_19_1 ));
    LocalMux I__16526 (
            .O(N__68595),
            .I(\ALU.status_19_1 ));
    Odrv4 I__16525 (
            .O(N__68588),
            .I(\ALU.status_19_1 ));
    InMux I__16524 (
            .O(N__68567),
            .I(N__68560));
    InMux I__16523 (
            .O(N__68566),
            .I(N__68560));
    InMux I__16522 (
            .O(N__68565),
            .I(N__68557));
    LocalMux I__16521 (
            .O(N__68560),
            .I(N__68553));
    LocalMux I__16520 (
            .O(N__68557),
            .I(N__68550));
    CascadeMux I__16519 (
            .O(N__68556),
            .I(N__68547));
    Span4Mux_v I__16518 (
            .O(N__68553),
            .I(N__68544));
    Span4Mux_v I__16517 (
            .O(N__68550),
            .I(N__68541));
    InMux I__16516 (
            .O(N__68547),
            .I(N__68538));
    Odrv4 I__16515 (
            .O(N__68544),
            .I(\ALU.N_968 ));
    Odrv4 I__16514 (
            .O(N__68541),
            .I(\ALU.N_968 ));
    LocalMux I__16513 (
            .O(N__68538),
            .I(\ALU.N_968 ));
    CascadeMux I__16512 (
            .O(N__68531),
            .I(N__68518));
    CascadeMux I__16511 (
            .O(N__68530),
            .I(N__68512));
    InMux I__16510 (
            .O(N__68529),
            .I(N__68502));
    InMux I__16509 (
            .O(N__68528),
            .I(N__68499));
    InMux I__16508 (
            .O(N__68527),
            .I(N__68494));
    InMux I__16507 (
            .O(N__68526),
            .I(N__68494));
    InMux I__16506 (
            .O(N__68525),
            .I(N__68491));
    InMux I__16505 (
            .O(N__68524),
            .I(N__68485));
    InMux I__16504 (
            .O(N__68523),
            .I(N__68485));
    InMux I__16503 (
            .O(N__68522),
            .I(N__68472));
    InMux I__16502 (
            .O(N__68521),
            .I(N__68472));
    InMux I__16501 (
            .O(N__68518),
            .I(N__68472));
    CascadeMux I__16500 (
            .O(N__68517),
            .I(N__68469));
    InMux I__16499 (
            .O(N__68516),
            .I(N__68465));
    InMux I__16498 (
            .O(N__68515),
            .I(N__68461));
    InMux I__16497 (
            .O(N__68512),
            .I(N__68455));
    InMux I__16496 (
            .O(N__68511),
            .I(N__68452));
    InMux I__16495 (
            .O(N__68510),
            .I(N__68445));
    InMux I__16494 (
            .O(N__68509),
            .I(N__68445));
    InMux I__16493 (
            .O(N__68508),
            .I(N__68445));
    InMux I__16492 (
            .O(N__68507),
            .I(N__68442));
    CascadeMux I__16491 (
            .O(N__68506),
            .I(N__68435));
    CascadeMux I__16490 (
            .O(N__68505),
            .I(N__68432));
    LocalMux I__16489 (
            .O(N__68502),
            .I(N__68426));
    LocalMux I__16488 (
            .O(N__68499),
            .I(N__68426));
    LocalMux I__16487 (
            .O(N__68494),
            .I(N__68423));
    LocalMux I__16486 (
            .O(N__68491),
            .I(N__68420));
    InMux I__16485 (
            .O(N__68490),
            .I(N__68417));
    LocalMux I__16484 (
            .O(N__68485),
            .I(N__68414));
    InMux I__16483 (
            .O(N__68484),
            .I(N__68411));
    InMux I__16482 (
            .O(N__68483),
            .I(N__68404));
    InMux I__16481 (
            .O(N__68482),
            .I(N__68404));
    InMux I__16480 (
            .O(N__68481),
            .I(N__68404));
    InMux I__16479 (
            .O(N__68480),
            .I(N__68399));
    InMux I__16478 (
            .O(N__68479),
            .I(N__68399));
    LocalMux I__16477 (
            .O(N__68472),
            .I(N__68396));
    InMux I__16476 (
            .O(N__68469),
            .I(N__68391));
    InMux I__16475 (
            .O(N__68468),
            .I(N__68388));
    LocalMux I__16474 (
            .O(N__68465),
            .I(N__68385));
    InMux I__16473 (
            .O(N__68464),
            .I(N__68382));
    LocalMux I__16472 (
            .O(N__68461),
            .I(N__68379));
    CascadeMux I__16471 (
            .O(N__68460),
            .I(N__68375));
    InMux I__16470 (
            .O(N__68459),
            .I(N__68371));
    InMux I__16469 (
            .O(N__68458),
            .I(N__68368));
    LocalMux I__16468 (
            .O(N__68455),
            .I(N__68359));
    LocalMux I__16467 (
            .O(N__68452),
            .I(N__68359));
    LocalMux I__16466 (
            .O(N__68445),
            .I(N__68359));
    LocalMux I__16465 (
            .O(N__68442),
            .I(N__68359));
    InMux I__16464 (
            .O(N__68441),
            .I(N__68352));
    InMux I__16463 (
            .O(N__68440),
            .I(N__68352));
    InMux I__16462 (
            .O(N__68439),
            .I(N__68352));
    InMux I__16461 (
            .O(N__68438),
            .I(N__68349));
    InMux I__16460 (
            .O(N__68435),
            .I(N__68346));
    InMux I__16459 (
            .O(N__68432),
            .I(N__68343));
    InMux I__16458 (
            .O(N__68431),
            .I(N__68340));
    Span4Mux_v I__16457 (
            .O(N__68426),
            .I(N__68329));
    Span4Mux_v I__16456 (
            .O(N__68423),
            .I(N__68329));
    Span4Mux_v I__16455 (
            .O(N__68420),
            .I(N__68329));
    LocalMux I__16454 (
            .O(N__68417),
            .I(N__68329));
    Span4Mux_v I__16453 (
            .O(N__68414),
            .I(N__68329));
    LocalMux I__16452 (
            .O(N__68411),
            .I(N__68322));
    LocalMux I__16451 (
            .O(N__68404),
            .I(N__68322));
    LocalMux I__16450 (
            .O(N__68399),
            .I(N__68322));
    Span4Mux_v I__16449 (
            .O(N__68396),
            .I(N__68319));
    InMux I__16448 (
            .O(N__68395),
            .I(N__68316));
    CascadeMux I__16447 (
            .O(N__68394),
            .I(N__68312));
    LocalMux I__16446 (
            .O(N__68391),
            .I(N__68309));
    LocalMux I__16445 (
            .O(N__68388),
            .I(N__68306));
    Span4Mux_v I__16444 (
            .O(N__68385),
            .I(N__68299));
    LocalMux I__16443 (
            .O(N__68382),
            .I(N__68299));
    Span4Mux_h I__16442 (
            .O(N__68379),
            .I(N__68299));
    InMux I__16441 (
            .O(N__68378),
            .I(N__68292));
    InMux I__16440 (
            .O(N__68375),
            .I(N__68292));
    InMux I__16439 (
            .O(N__68374),
            .I(N__68292));
    LocalMux I__16438 (
            .O(N__68371),
            .I(N__68285));
    LocalMux I__16437 (
            .O(N__68368),
            .I(N__68285));
    Span4Mux_v I__16436 (
            .O(N__68359),
            .I(N__68285));
    LocalMux I__16435 (
            .O(N__68352),
            .I(N__68282));
    LocalMux I__16434 (
            .O(N__68349),
            .I(N__68271));
    LocalMux I__16433 (
            .O(N__68346),
            .I(N__68271));
    LocalMux I__16432 (
            .O(N__68343),
            .I(N__68271));
    LocalMux I__16431 (
            .O(N__68340),
            .I(N__68271));
    Sp12to4 I__16430 (
            .O(N__68329),
            .I(N__68267));
    Span4Mux_v I__16429 (
            .O(N__68322),
            .I(N__68260));
    Span4Mux_h I__16428 (
            .O(N__68319),
            .I(N__68260));
    LocalMux I__16427 (
            .O(N__68316),
            .I(N__68260));
    InMux I__16426 (
            .O(N__68315),
            .I(N__68257));
    InMux I__16425 (
            .O(N__68312),
            .I(N__68253));
    Span4Mux_h I__16424 (
            .O(N__68309),
            .I(N__68240));
    Span4Mux_v I__16423 (
            .O(N__68306),
            .I(N__68240));
    Span4Mux_v I__16422 (
            .O(N__68299),
            .I(N__68240));
    LocalMux I__16421 (
            .O(N__68292),
            .I(N__68240));
    Span4Mux_h I__16420 (
            .O(N__68285),
            .I(N__68240));
    Span4Mux_h I__16419 (
            .O(N__68282),
            .I(N__68240));
    InMux I__16418 (
            .O(N__68281),
            .I(N__68237));
    CascadeMux I__16417 (
            .O(N__68280),
            .I(N__68234));
    Span4Mux_v I__16416 (
            .O(N__68271),
            .I(N__68225));
    InMux I__16415 (
            .O(N__68270),
            .I(N__68222));
    Span12Mux_h I__16414 (
            .O(N__68267),
            .I(N__68215));
    Sp12to4 I__16413 (
            .O(N__68260),
            .I(N__68215));
    LocalMux I__16412 (
            .O(N__68257),
            .I(N__68215));
    InMux I__16411 (
            .O(N__68256),
            .I(N__68212));
    LocalMux I__16410 (
            .O(N__68253),
            .I(N__68205));
    Span4Mux_h I__16409 (
            .O(N__68240),
            .I(N__68205));
    LocalMux I__16408 (
            .O(N__68237),
            .I(N__68205));
    InMux I__16407 (
            .O(N__68234),
            .I(N__68196));
    InMux I__16406 (
            .O(N__68233),
            .I(N__68196));
    InMux I__16405 (
            .O(N__68232),
            .I(N__68196));
    InMux I__16404 (
            .O(N__68231),
            .I(N__68196));
    InMux I__16403 (
            .O(N__68230),
            .I(N__68189));
    InMux I__16402 (
            .O(N__68229),
            .I(N__68189));
    InMux I__16401 (
            .O(N__68228),
            .I(N__68189));
    Odrv4 I__16400 (
            .O(N__68225),
            .I(\ALU.status_19_2 ));
    LocalMux I__16399 (
            .O(N__68222),
            .I(\ALU.status_19_2 ));
    Odrv12 I__16398 (
            .O(N__68215),
            .I(\ALU.status_19_2 ));
    LocalMux I__16397 (
            .O(N__68212),
            .I(\ALU.status_19_2 ));
    Odrv4 I__16396 (
            .O(N__68205),
            .I(\ALU.status_19_2 ));
    LocalMux I__16395 (
            .O(N__68196),
            .I(\ALU.status_19_2 ));
    LocalMux I__16394 (
            .O(N__68189),
            .I(\ALU.status_19_2 ));
    InMux I__16393 (
            .O(N__68174),
            .I(N__68171));
    LocalMux I__16392 (
            .O(N__68171),
            .I(N__68168));
    Span4Mux_v I__16391 (
            .O(N__68168),
            .I(N__68163));
    InMux I__16390 (
            .O(N__68167),
            .I(N__68158));
    InMux I__16389 (
            .O(N__68166),
            .I(N__68158));
    Sp12to4 I__16388 (
            .O(N__68163),
            .I(N__68153));
    LocalMux I__16387 (
            .O(N__68158),
            .I(N__68153));
    Odrv12 I__16386 (
            .O(N__68153),
            .I(\ALU.N_867 ));
    InMux I__16385 (
            .O(N__68150),
            .I(N__68147));
    LocalMux I__16384 (
            .O(N__68147),
            .I(\ALU.c_RNICBIG85Z0Z_15 ));
    InMux I__16383 (
            .O(N__68144),
            .I(N__68141));
    LocalMux I__16382 (
            .O(N__68141),
            .I(N__68133));
    InMux I__16381 (
            .O(N__68140),
            .I(N__68130));
    InMux I__16380 (
            .O(N__68139),
            .I(N__68127));
    InMux I__16379 (
            .O(N__68138),
            .I(N__68124));
    InMux I__16378 (
            .O(N__68137),
            .I(N__68119));
    InMux I__16377 (
            .O(N__68136),
            .I(N__68116));
    Span4Mux_v I__16376 (
            .O(N__68133),
            .I(N__68109));
    LocalMux I__16375 (
            .O(N__68130),
            .I(N__68109));
    LocalMux I__16374 (
            .O(N__68127),
            .I(N__68109));
    LocalMux I__16373 (
            .O(N__68124),
            .I(N__68106));
    InMux I__16372 (
            .O(N__68123),
            .I(N__68103));
    InMux I__16371 (
            .O(N__68122),
            .I(N__68100));
    LocalMux I__16370 (
            .O(N__68119),
            .I(\ALU.a_15_ns_snZ0Z_14 ));
    LocalMux I__16369 (
            .O(N__68116),
            .I(\ALU.a_15_ns_snZ0Z_14 ));
    Odrv4 I__16368 (
            .O(N__68109),
            .I(\ALU.a_15_ns_snZ0Z_14 ));
    Odrv4 I__16367 (
            .O(N__68106),
            .I(\ALU.a_15_ns_snZ0Z_14 ));
    LocalMux I__16366 (
            .O(N__68103),
            .I(\ALU.a_15_ns_snZ0Z_14 ));
    LocalMux I__16365 (
            .O(N__68100),
            .I(\ALU.a_15_ns_snZ0Z_14 ));
    InMux I__16364 (
            .O(N__68087),
            .I(N__68083));
    InMux I__16363 (
            .O(N__68086),
            .I(N__68080));
    LocalMux I__16362 (
            .O(N__68083),
            .I(N__68071));
    LocalMux I__16361 (
            .O(N__68080),
            .I(N__68071));
    InMux I__16360 (
            .O(N__68079),
            .I(N__68068));
    InMux I__16359 (
            .O(N__68078),
            .I(N__68065));
    InMux I__16358 (
            .O(N__68077),
            .I(N__68062));
    InMux I__16357 (
            .O(N__68076),
            .I(N__68059));
    Span4Mux_h I__16356 (
            .O(N__68071),
            .I(N__68054));
    LocalMux I__16355 (
            .O(N__68068),
            .I(N__68049));
    LocalMux I__16354 (
            .O(N__68065),
            .I(N__68049));
    LocalMux I__16353 (
            .O(N__68062),
            .I(N__68046));
    LocalMux I__16352 (
            .O(N__68059),
            .I(N__68043));
    InMux I__16351 (
            .O(N__68058),
            .I(N__68040));
    InMux I__16350 (
            .O(N__68057),
            .I(N__68037));
    Span4Mux_h I__16349 (
            .O(N__68054),
            .I(N__68034));
    Span4Mux_v I__16348 (
            .O(N__68049),
            .I(N__68023));
    Span4Mux_v I__16347 (
            .O(N__68046),
            .I(N__68023));
    Span4Mux_h I__16346 (
            .O(N__68043),
            .I(N__68023));
    LocalMux I__16345 (
            .O(N__68040),
            .I(N__68023));
    LocalMux I__16344 (
            .O(N__68037),
            .I(N__68023));
    Span4Mux_h I__16343 (
            .O(N__68034),
            .I(N__68020));
    Span4Mux_h I__16342 (
            .O(N__68023),
            .I(N__68017));
    Odrv4 I__16341 (
            .O(N__68020),
            .I(\ALU.lshift_14 ));
    Odrv4 I__16340 (
            .O(N__68017),
            .I(\ALU.lshift_14 ));
    InMux I__16339 (
            .O(N__68012),
            .I(N__68008));
    InMux I__16338 (
            .O(N__68011),
            .I(N__68005));
    LocalMux I__16337 (
            .O(N__68008),
            .I(N__67997));
    LocalMux I__16336 (
            .O(N__68005),
            .I(N__67994));
    InMux I__16335 (
            .O(N__68004),
            .I(N__67991));
    InMux I__16334 (
            .O(N__68003),
            .I(N__67988));
    InMux I__16333 (
            .O(N__68002),
            .I(N__67985));
    InMux I__16332 (
            .O(N__68001),
            .I(N__67982));
    InMux I__16331 (
            .O(N__68000),
            .I(N__67979));
    Odrv4 I__16330 (
            .O(N__67997),
            .I(\ALU.a_15_ns_rn_0_14 ));
    Odrv4 I__16329 (
            .O(N__67994),
            .I(\ALU.a_15_ns_rn_0_14 ));
    LocalMux I__16328 (
            .O(N__67991),
            .I(\ALU.a_15_ns_rn_0_14 ));
    LocalMux I__16327 (
            .O(N__67988),
            .I(\ALU.a_15_ns_rn_0_14 ));
    LocalMux I__16326 (
            .O(N__67985),
            .I(\ALU.a_15_ns_rn_0_14 ));
    LocalMux I__16325 (
            .O(N__67982),
            .I(\ALU.a_15_ns_rn_0_14 ));
    LocalMux I__16324 (
            .O(N__67979),
            .I(\ALU.a_15_ns_rn_0_14 ));
    InMux I__16323 (
            .O(N__67964),
            .I(N__67960));
    InMux I__16322 (
            .O(N__67963),
            .I(N__67957));
    LocalMux I__16321 (
            .O(N__67960),
            .I(N__67952));
    LocalMux I__16320 (
            .O(N__67957),
            .I(N__67952));
    Span4Mux_v I__16319 (
            .O(N__67952),
            .I(N__67949));
    Span4Mux_h I__16318 (
            .O(N__67949),
            .I(N__67946));
    Odrv4 I__16317 (
            .O(N__67946),
            .I(\ALU.bZ0Z_14 ));
    CEMux I__16316 (
            .O(N__67943),
            .I(N__67939));
    CEMux I__16315 (
            .O(N__67942),
            .I(N__67935));
    LocalMux I__16314 (
            .O(N__67939),
            .I(N__67932));
    CEMux I__16313 (
            .O(N__67938),
            .I(N__67928));
    LocalMux I__16312 (
            .O(N__67935),
            .I(N__67925));
    Span4Mux_v I__16311 (
            .O(N__67932),
            .I(N__67922));
    CEMux I__16310 (
            .O(N__67931),
            .I(N__67918));
    LocalMux I__16309 (
            .O(N__67928),
            .I(N__67915));
    Span4Mux_v I__16308 (
            .O(N__67925),
            .I(N__67912));
    Span4Mux_h I__16307 (
            .O(N__67922),
            .I(N__67909));
    CEMux I__16306 (
            .O(N__67921),
            .I(N__67906));
    LocalMux I__16305 (
            .O(N__67918),
            .I(N__67903));
    Span4Mux_h I__16304 (
            .O(N__67915),
            .I(N__67900));
    Span4Mux_h I__16303 (
            .O(N__67912),
            .I(N__67897));
    Span4Mux_v I__16302 (
            .O(N__67909),
            .I(N__67894));
    LocalMux I__16301 (
            .O(N__67906),
            .I(N__67891));
    Span4Mux_h I__16300 (
            .O(N__67903),
            .I(N__67888));
    Span4Mux_h I__16299 (
            .O(N__67900),
            .I(N__67885));
    Span4Mux_v I__16298 (
            .O(N__67897),
            .I(N__67880));
    Span4Mux_h I__16297 (
            .O(N__67894),
            .I(N__67880));
    Odrv12 I__16296 (
            .O(N__67891),
            .I(\ALU.un1_a41_8_0 ));
    Odrv4 I__16295 (
            .O(N__67888),
            .I(\ALU.un1_a41_8_0 ));
    Odrv4 I__16294 (
            .O(N__67885),
            .I(\ALU.un1_a41_8_0 ));
    Odrv4 I__16293 (
            .O(N__67880),
            .I(\ALU.un1_a41_8_0 ));
    CEMux I__16292 (
            .O(N__67871),
            .I(N__67868));
    LocalMux I__16291 (
            .O(N__67868),
            .I(N__67865));
    Span4Mux_v I__16290 (
            .O(N__67865),
            .I(N__67861));
    CEMux I__16289 (
            .O(N__67864),
            .I(N__67857));
    Span4Mux_h I__16288 (
            .O(N__67861),
            .I(N__67854));
    CEMux I__16287 (
            .O(N__67860),
            .I(N__67851));
    LocalMux I__16286 (
            .O(N__67857),
            .I(N__67848));
    Span4Mux_h I__16285 (
            .O(N__67854),
            .I(N__67845));
    LocalMux I__16284 (
            .O(N__67851),
            .I(N__67842));
    Sp12to4 I__16283 (
            .O(N__67848),
            .I(N__67839));
    Span4Mux_h I__16282 (
            .O(N__67845),
            .I(N__67836));
    Span4Mux_v I__16281 (
            .O(N__67842),
            .I(N__67833));
    Span12Mux_s11_v I__16280 (
            .O(N__67839),
            .I(N__67830));
    Sp12to4 I__16279 (
            .O(N__67836),
            .I(N__67827));
    Odrv4 I__16278 (
            .O(N__67833),
            .I(\ALU.un1_a41_4_0 ));
    Odrv12 I__16277 (
            .O(N__67830),
            .I(\ALU.un1_a41_4_0 ));
    Odrv12 I__16276 (
            .O(N__67827),
            .I(\ALU.un1_a41_4_0 ));
    InMux I__16275 (
            .O(N__67820),
            .I(N__67817));
    LocalMux I__16274 (
            .O(N__67817),
            .I(N__67814));
    Span12Mux_v I__16273 (
            .O(N__67814),
            .I(N__67811));
    Odrv12 I__16272 (
            .O(N__67811),
            .I(\ALU.un1_operation_5_0 ));
    CascadeMux I__16271 (
            .O(N__67808),
            .I(N__67805));
    InMux I__16270 (
            .O(N__67805),
            .I(N__67802));
    LocalMux I__16269 (
            .O(N__67802),
            .I(N__67799));
    Span4Mux_v I__16268 (
            .O(N__67799),
            .I(N__67796));
    Sp12to4 I__16267 (
            .O(N__67796),
            .I(N__67793));
    Span12Mux_h I__16266 (
            .O(N__67793),
            .I(N__67790));
    Odrv12 I__16265 (
            .O(N__67790),
            .I(aluOperation_5));
    CascadeMux I__16264 (
            .O(N__67787),
            .I(\ALU.un1_operation_10_0_cascade_ ));
    InMux I__16263 (
            .O(N__67784),
            .I(N__67780));
    InMux I__16262 (
            .O(N__67783),
            .I(N__67777));
    LocalMux I__16261 (
            .O(N__67780),
            .I(N__67774));
    LocalMux I__16260 (
            .O(N__67777),
            .I(N__67771));
    Span4Mux_v I__16259 (
            .O(N__67774),
            .I(N__67766));
    Span4Mux_h I__16258 (
            .O(N__67771),
            .I(N__67766));
    Span4Mux_h I__16257 (
            .O(N__67766),
            .I(N__67763));
    Sp12to4 I__16256 (
            .O(N__67763),
            .I(N__67760));
    Odrv12 I__16255 (
            .O(N__67760),
            .I(\ALU.dZ0Z_14 ));
    InMux I__16254 (
            .O(N__67757),
            .I(N__67750));
    InMux I__16253 (
            .O(N__67756),
            .I(N__67747));
    InMux I__16252 (
            .O(N__67755),
            .I(N__67744));
    InMux I__16251 (
            .O(N__67754),
            .I(N__67738));
    InMux I__16250 (
            .O(N__67753),
            .I(N__67735));
    LocalMux I__16249 (
            .O(N__67750),
            .I(N__67732));
    LocalMux I__16248 (
            .O(N__67747),
            .I(N__67729));
    LocalMux I__16247 (
            .O(N__67744),
            .I(N__67726));
    InMux I__16246 (
            .O(N__67743),
            .I(N__67723));
    InMux I__16245 (
            .O(N__67742),
            .I(N__67720));
    InMux I__16244 (
            .O(N__67741),
            .I(N__67717));
    LocalMux I__16243 (
            .O(N__67738),
            .I(N__67712));
    LocalMux I__16242 (
            .O(N__67735),
            .I(N__67712));
    Span4Mux_h I__16241 (
            .O(N__67732),
            .I(N__67707));
    Span4Mux_h I__16240 (
            .O(N__67729),
            .I(N__67707));
    Span12Mux_v I__16239 (
            .O(N__67726),
            .I(N__67704));
    LocalMux I__16238 (
            .O(N__67723),
            .I(\ALU.c_RNIBRG4Q9Z0Z_12 ));
    LocalMux I__16237 (
            .O(N__67720),
            .I(\ALU.c_RNIBRG4Q9Z0Z_12 ));
    LocalMux I__16236 (
            .O(N__67717),
            .I(\ALU.c_RNIBRG4Q9Z0Z_12 ));
    Odrv12 I__16235 (
            .O(N__67712),
            .I(\ALU.c_RNIBRG4Q9Z0Z_12 ));
    Odrv4 I__16234 (
            .O(N__67707),
            .I(\ALU.c_RNIBRG4Q9Z0Z_12 ));
    Odrv12 I__16233 (
            .O(N__67704),
            .I(\ALU.c_RNIBRG4Q9Z0Z_12 ));
    InMux I__16232 (
            .O(N__67691),
            .I(N__67688));
    LocalMux I__16231 (
            .O(N__67688),
            .I(N__67682));
    InMux I__16230 (
            .O(N__67687),
            .I(N__67679));
    InMux I__16229 (
            .O(N__67686),
            .I(N__67676));
    InMux I__16228 (
            .O(N__67685),
            .I(N__67673));
    Span4Mux_v I__16227 (
            .O(N__67682),
            .I(N__67669));
    LocalMux I__16226 (
            .O(N__67679),
            .I(N__67665));
    LocalMux I__16225 (
            .O(N__67676),
            .I(N__67662));
    LocalMux I__16224 (
            .O(N__67673),
            .I(N__67659));
    InMux I__16223 (
            .O(N__67672),
            .I(N__67656));
    Span4Mux_h I__16222 (
            .O(N__67669),
            .I(N__67651));
    InMux I__16221 (
            .O(N__67668),
            .I(N__67648));
    Span4Mux_v I__16220 (
            .O(N__67665),
            .I(N__67639));
    Span4Mux_v I__16219 (
            .O(N__67662),
            .I(N__67639));
    Span4Mux_h I__16218 (
            .O(N__67659),
            .I(N__67639));
    LocalMux I__16217 (
            .O(N__67656),
            .I(N__67639));
    InMux I__16216 (
            .O(N__67655),
            .I(N__67636));
    InMux I__16215 (
            .O(N__67654),
            .I(N__67633));
    Odrv4 I__16214 (
            .O(N__67651),
            .I(\ALU.c_RNIBRG4Q9_0Z0Z_12 ));
    LocalMux I__16213 (
            .O(N__67648),
            .I(\ALU.c_RNIBRG4Q9_0Z0Z_12 ));
    Odrv4 I__16212 (
            .O(N__67639),
            .I(\ALU.c_RNIBRG4Q9_0Z0Z_12 ));
    LocalMux I__16211 (
            .O(N__67636),
            .I(\ALU.c_RNIBRG4Q9_0Z0Z_12 ));
    LocalMux I__16210 (
            .O(N__67633),
            .I(\ALU.c_RNIBRG4Q9_0Z0Z_12 ));
    CascadeMux I__16209 (
            .O(N__67622),
            .I(N__67618));
    InMux I__16208 (
            .O(N__67621),
            .I(N__67614));
    InMux I__16207 (
            .O(N__67618),
            .I(N__67611));
    InMux I__16206 (
            .O(N__67617),
            .I(N__67607));
    LocalMux I__16205 (
            .O(N__67614),
            .I(N__67604));
    LocalMux I__16204 (
            .O(N__67611),
            .I(N__67599));
    InMux I__16203 (
            .O(N__67610),
            .I(N__67596));
    LocalMux I__16202 (
            .O(N__67607),
            .I(N__67590));
    Span4Mux_v I__16201 (
            .O(N__67604),
            .I(N__67590));
    InMux I__16200 (
            .O(N__67603),
            .I(N__67587));
    CascadeMux I__16199 (
            .O(N__67602),
            .I(N__67584));
    Span4Mux_v I__16198 (
            .O(N__67599),
            .I(N__67581));
    LocalMux I__16197 (
            .O(N__67596),
            .I(N__67578));
    InMux I__16196 (
            .O(N__67595),
            .I(N__67575));
    Span4Mux_v I__16195 (
            .O(N__67590),
            .I(N__67570));
    LocalMux I__16194 (
            .O(N__67587),
            .I(N__67570));
    InMux I__16193 (
            .O(N__67584),
            .I(N__67567));
    Odrv4 I__16192 (
            .O(N__67581),
            .I(\ALU.mult_555_c_RNIJF56AMZ0 ));
    Odrv4 I__16191 (
            .O(N__67578),
            .I(\ALU.mult_555_c_RNIJF56AMZ0 ));
    LocalMux I__16190 (
            .O(N__67575),
            .I(\ALU.mult_555_c_RNIJF56AMZ0 ));
    Odrv4 I__16189 (
            .O(N__67570),
            .I(\ALU.mult_555_c_RNIJF56AMZ0 ));
    LocalMux I__16188 (
            .O(N__67567),
            .I(\ALU.mult_555_c_RNIJF56AMZ0 ));
    InMux I__16187 (
            .O(N__67556),
            .I(N__67553));
    LocalMux I__16186 (
            .O(N__67553),
            .I(N__67550));
    Span4Mux_v I__16185 (
            .O(N__67550),
            .I(N__67546));
    InMux I__16184 (
            .O(N__67549),
            .I(N__67543));
    Span4Mux_h I__16183 (
            .O(N__67546),
            .I(N__67538));
    LocalMux I__16182 (
            .O(N__67543),
            .I(N__67538));
    Span4Mux_h I__16181 (
            .O(N__67538),
            .I(N__67535));
    Span4Mux_h I__16180 (
            .O(N__67535),
            .I(N__67532));
    Span4Mux_h I__16179 (
            .O(N__67532),
            .I(N__67529));
    Span4Mux_h I__16178 (
            .O(N__67529),
            .I(N__67526));
    Span4Mux_v I__16177 (
            .O(N__67526),
            .I(N__67523));
    Span4Mux_h I__16176 (
            .O(N__67523),
            .I(N__67520));
    Odrv4 I__16175 (
            .O(N__67520),
            .I(\ALU.cZ0Z_12 ));
    InMux I__16174 (
            .O(N__67517),
            .I(N__67513));
    InMux I__16173 (
            .O(N__67516),
            .I(N__67509));
    LocalMux I__16172 (
            .O(N__67513),
            .I(N__67505));
    InMux I__16171 (
            .O(N__67512),
            .I(N__67501));
    LocalMux I__16170 (
            .O(N__67509),
            .I(N__67498));
    InMux I__16169 (
            .O(N__67508),
            .I(N__67495));
    Span4Mux_v I__16168 (
            .O(N__67505),
            .I(N__67490));
    InMux I__16167 (
            .O(N__67504),
            .I(N__67487));
    LocalMux I__16166 (
            .O(N__67501),
            .I(N__67484));
    Span4Mux_v I__16165 (
            .O(N__67498),
            .I(N__67479));
    LocalMux I__16164 (
            .O(N__67495),
            .I(N__67479));
    InMux I__16163 (
            .O(N__67494),
            .I(N__67476));
    InMux I__16162 (
            .O(N__67493),
            .I(N__67473));
    Odrv4 I__16161 (
            .O(N__67490),
            .I(\ALU.c_RNIO5N04A_0Z0Z_13 ));
    LocalMux I__16160 (
            .O(N__67487),
            .I(\ALU.c_RNIO5N04A_0Z0Z_13 ));
    Odrv4 I__16159 (
            .O(N__67484),
            .I(\ALU.c_RNIO5N04A_0Z0Z_13 ));
    Odrv4 I__16158 (
            .O(N__67479),
            .I(\ALU.c_RNIO5N04A_0Z0Z_13 ));
    LocalMux I__16157 (
            .O(N__67476),
            .I(\ALU.c_RNIO5N04A_0Z0Z_13 ));
    LocalMux I__16156 (
            .O(N__67473),
            .I(\ALU.c_RNIO5N04A_0Z0Z_13 ));
    InMux I__16155 (
            .O(N__67460),
            .I(N__67456));
    InMux I__16154 (
            .O(N__67459),
            .I(N__67452));
    LocalMux I__16153 (
            .O(N__67456),
            .I(N__67446));
    InMux I__16152 (
            .O(N__67455),
            .I(N__67443));
    LocalMux I__16151 (
            .O(N__67452),
            .I(N__67439));
    InMux I__16150 (
            .O(N__67451),
            .I(N__67436));
    InMux I__16149 (
            .O(N__67450),
            .I(N__67433));
    InMux I__16148 (
            .O(N__67449),
            .I(N__67429));
    Span4Mux_h I__16147 (
            .O(N__67446),
            .I(N__67424));
    LocalMux I__16146 (
            .O(N__67443),
            .I(N__67424));
    InMux I__16145 (
            .O(N__67442),
            .I(N__67421));
    Span4Mux_v I__16144 (
            .O(N__67439),
            .I(N__67414));
    LocalMux I__16143 (
            .O(N__67436),
            .I(N__67414));
    LocalMux I__16142 (
            .O(N__67433),
            .I(N__67414));
    InMux I__16141 (
            .O(N__67432),
            .I(N__67411));
    LocalMux I__16140 (
            .O(N__67429),
            .I(\ALU.c_RNIO5N04AZ0Z_13 ));
    Odrv4 I__16139 (
            .O(N__67424),
            .I(\ALU.c_RNIO5N04AZ0Z_13 ));
    LocalMux I__16138 (
            .O(N__67421),
            .I(\ALU.c_RNIO5N04AZ0Z_13 ));
    Odrv4 I__16137 (
            .O(N__67414),
            .I(\ALU.c_RNIO5N04AZ0Z_13 ));
    LocalMux I__16136 (
            .O(N__67411),
            .I(\ALU.c_RNIO5N04AZ0Z_13 ));
    InMux I__16135 (
            .O(N__67400),
            .I(N__67396));
    InMux I__16134 (
            .O(N__67399),
            .I(N__67393));
    LocalMux I__16133 (
            .O(N__67396),
            .I(N__67385));
    LocalMux I__16132 (
            .O(N__67393),
            .I(N__67382));
    InMux I__16131 (
            .O(N__67392),
            .I(N__67379));
    InMux I__16130 (
            .O(N__67391),
            .I(N__67376));
    InMux I__16129 (
            .O(N__67390),
            .I(N__67373));
    InMux I__16128 (
            .O(N__67389),
            .I(N__67370));
    InMux I__16127 (
            .O(N__67388),
            .I(N__67367));
    Odrv4 I__16126 (
            .O(N__67385),
            .I(\ALU.mult_558_c_RNIB75F9GZ0 ));
    Odrv4 I__16125 (
            .O(N__67382),
            .I(\ALU.mult_558_c_RNIB75F9GZ0 ));
    LocalMux I__16124 (
            .O(N__67379),
            .I(\ALU.mult_558_c_RNIB75F9GZ0 ));
    LocalMux I__16123 (
            .O(N__67376),
            .I(\ALU.mult_558_c_RNIB75F9GZ0 ));
    LocalMux I__16122 (
            .O(N__67373),
            .I(\ALU.mult_558_c_RNIB75F9GZ0 ));
    LocalMux I__16121 (
            .O(N__67370),
            .I(\ALU.mult_558_c_RNIB75F9GZ0 ));
    LocalMux I__16120 (
            .O(N__67367),
            .I(\ALU.mult_558_c_RNIB75F9GZ0 ));
    InMux I__16119 (
            .O(N__67352),
            .I(N__67349));
    LocalMux I__16118 (
            .O(N__67349),
            .I(N__67345));
    InMux I__16117 (
            .O(N__67348),
            .I(N__67342));
    Span4Mux_h I__16116 (
            .O(N__67345),
            .I(N__67339));
    LocalMux I__16115 (
            .O(N__67342),
            .I(N__67336));
    Span4Mux_v I__16114 (
            .O(N__67339),
            .I(N__67333));
    Span4Mux_v I__16113 (
            .O(N__67336),
            .I(N__67330));
    Span4Mux_h I__16112 (
            .O(N__67333),
            .I(N__67327));
    Span4Mux_v I__16111 (
            .O(N__67330),
            .I(N__67324));
    Span4Mux_h I__16110 (
            .O(N__67327),
            .I(N__67321));
    Span4Mux_h I__16109 (
            .O(N__67324),
            .I(N__67316));
    Span4Mux_v I__16108 (
            .O(N__67321),
            .I(N__67316));
    Odrv4 I__16107 (
            .O(N__67316),
            .I(\ALU.cZ0Z_13 ));
    InMux I__16106 (
            .O(N__67313),
            .I(N__67309));
    InMux I__16105 (
            .O(N__67312),
            .I(N__67306));
    LocalMux I__16104 (
            .O(N__67309),
            .I(N__67303));
    LocalMux I__16103 (
            .O(N__67306),
            .I(N__67300));
    Span4Mux_v I__16102 (
            .O(N__67303),
            .I(N__67297));
    Span4Mux_v I__16101 (
            .O(N__67300),
            .I(N__67294));
    Span4Mux_h I__16100 (
            .O(N__67297),
            .I(N__67289));
    Span4Mux_h I__16099 (
            .O(N__67294),
            .I(N__67289));
    Odrv4 I__16098 (
            .O(N__67289),
            .I(\ALU.cZ0Z_14 ));
    CascadeMux I__16097 (
            .O(N__67286),
            .I(N__67283));
    InMux I__16096 (
            .O(N__67283),
            .I(N__67277));
    InMux I__16095 (
            .O(N__67282),
            .I(N__67277));
    LocalMux I__16094 (
            .O(N__67277),
            .I(N__67274));
    Span4Mux_v I__16093 (
            .O(N__67274),
            .I(N__67263));
    InMux I__16092 (
            .O(N__67273),
            .I(N__67256));
    InMux I__16091 (
            .O(N__67272),
            .I(N__67256));
    InMux I__16090 (
            .O(N__67271),
            .I(N__67256));
    CascadeMux I__16089 (
            .O(N__67270),
            .I(N__67245));
    InMux I__16088 (
            .O(N__67269),
            .I(N__67239));
    CascadeMux I__16087 (
            .O(N__67268),
            .I(N__67236));
    CascadeMux I__16086 (
            .O(N__67267),
            .I(N__67233));
    CascadeMux I__16085 (
            .O(N__67266),
            .I(N__67227));
    Span4Mux_h I__16084 (
            .O(N__67263),
            .I(N__67220));
    LocalMux I__16083 (
            .O(N__67256),
            .I(N__67220));
    CascadeMux I__16082 (
            .O(N__67255),
            .I(N__67209));
    InMux I__16081 (
            .O(N__67254),
            .I(N__67197));
    InMux I__16080 (
            .O(N__67253),
            .I(N__67197));
    InMux I__16079 (
            .O(N__67252),
            .I(N__67197));
    InMux I__16078 (
            .O(N__67251),
            .I(N__67184));
    InMux I__16077 (
            .O(N__67250),
            .I(N__67184));
    InMux I__16076 (
            .O(N__67249),
            .I(N__67184));
    InMux I__16075 (
            .O(N__67248),
            .I(N__67184));
    InMux I__16074 (
            .O(N__67245),
            .I(N__67184));
    InMux I__16073 (
            .O(N__67244),
            .I(N__67184));
    CascadeMux I__16072 (
            .O(N__67243),
            .I(N__67180));
    CascadeMux I__16071 (
            .O(N__67242),
            .I(N__67176));
    LocalMux I__16070 (
            .O(N__67239),
            .I(N__67173));
    InMux I__16069 (
            .O(N__67236),
            .I(N__67170));
    InMux I__16068 (
            .O(N__67233),
            .I(N__67165));
    InMux I__16067 (
            .O(N__67232),
            .I(N__67165));
    InMux I__16066 (
            .O(N__67231),
            .I(N__67161));
    InMux I__16065 (
            .O(N__67230),
            .I(N__67158));
    InMux I__16064 (
            .O(N__67227),
            .I(N__67151));
    InMux I__16063 (
            .O(N__67226),
            .I(N__67151));
    InMux I__16062 (
            .O(N__67225),
            .I(N__67151));
    Span4Mux_v I__16061 (
            .O(N__67220),
            .I(N__67148));
    InMux I__16060 (
            .O(N__67219),
            .I(N__67145));
    InMux I__16059 (
            .O(N__67218),
            .I(N__67138));
    InMux I__16058 (
            .O(N__67217),
            .I(N__67138));
    InMux I__16057 (
            .O(N__67216),
            .I(N__67138));
    InMux I__16056 (
            .O(N__67215),
            .I(N__67135));
    InMux I__16055 (
            .O(N__67214),
            .I(N__67130));
    InMux I__16054 (
            .O(N__67213),
            .I(N__67130));
    InMux I__16053 (
            .O(N__67212),
            .I(N__67123));
    InMux I__16052 (
            .O(N__67209),
            .I(N__67123));
    InMux I__16051 (
            .O(N__67208),
            .I(N__67123));
    InMux I__16050 (
            .O(N__67207),
            .I(N__67116));
    InMux I__16049 (
            .O(N__67206),
            .I(N__67116));
    InMux I__16048 (
            .O(N__67205),
            .I(N__67116));
    CascadeMux I__16047 (
            .O(N__67204),
            .I(N__67112));
    LocalMux I__16046 (
            .O(N__67197),
            .I(N__67107));
    LocalMux I__16045 (
            .O(N__67184),
            .I(N__67107));
    InMux I__16044 (
            .O(N__67183),
            .I(N__67100));
    InMux I__16043 (
            .O(N__67180),
            .I(N__67100));
    InMux I__16042 (
            .O(N__67179),
            .I(N__67100));
    InMux I__16041 (
            .O(N__67176),
            .I(N__67097));
    Span4Mux_h I__16040 (
            .O(N__67173),
            .I(N__67090));
    LocalMux I__16039 (
            .O(N__67170),
            .I(N__67090));
    LocalMux I__16038 (
            .O(N__67165),
            .I(N__67090));
    InMux I__16037 (
            .O(N__67164),
            .I(N__67087));
    LocalMux I__16036 (
            .O(N__67161),
            .I(N__67066));
    LocalMux I__16035 (
            .O(N__67158),
            .I(N__67066));
    LocalMux I__16034 (
            .O(N__67151),
            .I(N__67066));
    Span4Mux_v I__16033 (
            .O(N__67148),
            .I(N__67066));
    LocalMux I__16032 (
            .O(N__67145),
            .I(N__67066));
    LocalMux I__16031 (
            .O(N__67138),
            .I(N__67066));
    LocalMux I__16030 (
            .O(N__67135),
            .I(N__67066));
    LocalMux I__16029 (
            .O(N__67130),
            .I(N__67066));
    LocalMux I__16028 (
            .O(N__67123),
            .I(N__67066));
    LocalMux I__16027 (
            .O(N__67116),
            .I(N__67066));
    CascadeMux I__16026 (
            .O(N__67115),
            .I(N__67061));
    InMux I__16025 (
            .O(N__67112),
            .I(N__67057));
    Span4Mux_v I__16024 (
            .O(N__67107),
            .I(N__67054));
    LocalMux I__16023 (
            .O(N__67100),
            .I(N__67048));
    LocalMux I__16022 (
            .O(N__67097),
            .I(N__67039));
    Span4Mux_v I__16021 (
            .O(N__67090),
            .I(N__67036));
    LocalMux I__16020 (
            .O(N__67087),
            .I(N__67033));
    Span4Mux_v I__16019 (
            .O(N__67066),
            .I(N__67030));
    InMux I__16018 (
            .O(N__67065),
            .I(N__67027));
    InMux I__16017 (
            .O(N__67064),
            .I(N__67020));
    InMux I__16016 (
            .O(N__67061),
            .I(N__67020));
    InMux I__16015 (
            .O(N__67060),
            .I(N__67020));
    LocalMux I__16014 (
            .O(N__67057),
            .I(N__67017));
    Span4Mux_h I__16013 (
            .O(N__67054),
            .I(N__67014));
    InMux I__16012 (
            .O(N__67053),
            .I(N__67007));
    InMux I__16011 (
            .O(N__67052),
            .I(N__67007));
    InMux I__16010 (
            .O(N__67051),
            .I(N__67007));
    Span4Mux_v I__16009 (
            .O(N__67048),
            .I(N__67004));
    InMux I__16008 (
            .O(N__67047),
            .I(N__66997));
    InMux I__16007 (
            .O(N__67046),
            .I(N__66997));
    InMux I__16006 (
            .O(N__67045),
            .I(N__66997));
    InMux I__16005 (
            .O(N__67044),
            .I(N__66994));
    InMux I__16004 (
            .O(N__67043),
            .I(N__66991));
    InMux I__16003 (
            .O(N__67042),
            .I(N__66988));
    Span4Mux_v I__16002 (
            .O(N__67039),
            .I(N__66985));
    Span4Mux_h I__16001 (
            .O(N__67036),
            .I(N__66982));
    Span4Mux_v I__16000 (
            .O(N__67033),
            .I(N__66977));
    Span4Mux_h I__15999 (
            .O(N__67030),
            .I(N__66977));
    LocalMux I__15998 (
            .O(N__67027),
            .I(N__66973));
    LocalMux I__15997 (
            .O(N__67020),
            .I(N__66970));
    Span4Mux_h I__15996 (
            .O(N__67017),
            .I(N__66963));
    Span4Mux_h I__15995 (
            .O(N__67014),
            .I(N__66963));
    LocalMux I__15994 (
            .O(N__67007),
            .I(N__66963));
    Span4Mux_h I__15993 (
            .O(N__67004),
            .I(N__66958));
    LocalMux I__15992 (
            .O(N__66997),
            .I(N__66958));
    LocalMux I__15991 (
            .O(N__66994),
            .I(N__66951));
    LocalMux I__15990 (
            .O(N__66991),
            .I(N__66951));
    LocalMux I__15989 (
            .O(N__66988),
            .I(N__66951));
    Span4Mux_h I__15988 (
            .O(N__66985),
            .I(N__66948));
    Span4Mux_h I__15987 (
            .O(N__66982),
            .I(N__66945));
    Span4Mux_v I__15986 (
            .O(N__66977),
            .I(N__66942));
    InMux I__15985 (
            .O(N__66976),
            .I(N__66939));
    Span4Mux_v I__15984 (
            .O(N__66973),
            .I(N__66930));
    Span4Mux_v I__15983 (
            .O(N__66970),
            .I(N__66930));
    Span4Mux_v I__15982 (
            .O(N__66963),
            .I(N__66930));
    Span4Mux_h I__15981 (
            .O(N__66958),
            .I(N__66930));
    Sp12to4 I__15980 (
            .O(N__66951),
            .I(N__66927));
    Sp12to4 I__15979 (
            .O(N__66948),
            .I(N__66920));
    Sp12to4 I__15978 (
            .O(N__66945),
            .I(N__66920));
    Sp12to4 I__15977 (
            .O(N__66942),
            .I(N__66920));
    LocalMux I__15976 (
            .O(N__66939),
            .I(N__66915));
    Span4Mux_h I__15975 (
            .O(N__66930),
            .I(N__66915));
    Span12Mux_v I__15974 (
            .O(N__66927),
            .I(N__66910));
    Span12Mux_h I__15973 (
            .O(N__66920),
            .I(N__66910));
    Span4Mux_v I__15972 (
            .O(N__66915),
            .I(N__66907));
    Odrv12 I__15971 (
            .O(N__66910),
            .I(aluOperation_0));
    Odrv4 I__15970 (
            .O(N__66907),
            .I(aluOperation_0));
    CascadeMux I__15969 (
            .O(N__66902),
            .I(N__66898));
    InMux I__15968 (
            .O(N__66901),
            .I(N__66891));
    InMux I__15967 (
            .O(N__66898),
            .I(N__66891));
    CascadeMux I__15966 (
            .O(N__66897),
            .I(N__66888));
    InMux I__15965 (
            .O(N__66896),
            .I(N__66885));
    LocalMux I__15964 (
            .O(N__66891),
            .I(N__66882));
    InMux I__15963 (
            .O(N__66888),
            .I(N__66879));
    LocalMux I__15962 (
            .O(N__66885),
            .I(N__66876));
    Span4Mux_v I__15961 (
            .O(N__66882),
            .I(N__66873));
    LocalMux I__15960 (
            .O(N__66879),
            .I(N__66870));
    Span4Mux_v I__15959 (
            .O(N__66876),
            .I(N__66865));
    Span4Mux_h I__15958 (
            .O(N__66873),
            .I(N__66865));
    Odrv4 I__15957 (
            .O(N__66870),
            .I(\ALU.a_15_d_sZ0Z_10 ));
    Odrv4 I__15956 (
            .O(N__66865),
            .I(\ALU.a_15_d_sZ0Z_10 ));
    InMux I__15955 (
            .O(N__66860),
            .I(N__66857));
    LocalMux I__15954 (
            .O(N__66857),
            .I(N__66853));
    InMux I__15953 (
            .O(N__66856),
            .I(N__66850));
    Odrv4 I__15952 (
            .O(N__66853),
            .I(\ALU.addsub_9 ));
    LocalMux I__15951 (
            .O(N__66850),
            .I(\ALU.addsub_9 ));
    InMux I__15950 (
            .O(N__66845),
            .I(N__66840));
    InMux I__15949 (
            .O(N__66844),
            .I(N__66837));
    InMux I__15948 (
            .O(N__66843),
            .I(N__66834));
    LocalMux I__15947 (
            .O(N__66840),
            .I(N__66828));
    LocalMux I__15946 (
            .O(N__66837),
            .I(N__66822));
    LocalMux I__15945 (
            .O(N__66834),
            .I(N__66822));
    InMux I__15944 (
            .O(N__66833),
            .I(N__66819));
    InMux I__15943 (
            .O(N__66832),
            .I(N__66816));
    InMux I__15942 (
            .O(N__66831),
            .I(N__66813));
    Span4Mux_v I__15941 (
            .O(N__66828),
            .I(N__66810));
    InMux I__15940 (
            .O(N__66827),
            .I(N__66807));
    Sp12to4 I__15939 (
            .O(N__66822),
            .I(N__66801));
    LocalMux I__15938 (
            .O(N__66819),
            .I(N__66801));
    LocalMux I__15937 (
            .O(N__66816),
            .I(N__66796));
    LocalMux I__15936 (
            .O(N__66813),
            .I(N__66796));
    Span4Mux_v I__15935 (
            .O(N__66810),
            .I(N__66791));
    LocalMux I__15934 (
            .O(N__66807),
            .I(N__66791));
    InMux I__15933 (
            .O(N__66806),
            .I(N__66788));
    Span12Mux_v I__15932 (
            .O(N__66801),
            .I(N__66785));
    Span4Mux_v I__15931 (
            .O(N__66796),
            .I(N__66778));
    Span4Mux_h I__15930 (
            .O(N__66791),
            .I(N__66778));
    LocalMux I__15929 (
            .O(N__66788),
            .I(N__66778));
    Odrv12 I__15928 (
            .O(N__66785),
            .I(\ALU.a_15_d_ns_sx_9 ));
    Odrv4 I__15927 (
            .O(N__66778),
            .I(\ALU.a_15_d_ns_sx_9 ));
    CascadeMux I__15926 (
            .O(N__66773),
            .I(N__66769));
    InMux I__15925 (
            .O(N__66772),
            .I(N__66758));
    InMux I__15924 (
            .O(N__66769),
            .I(N__66750));
    InMux I__15923 (
            .O(N__66768),
            .I(N__66747));
    CascadeMux I__15922 (
            .O(N__66767),
            .I(N__66743));
    InMux I__15921 (
            .O(N__66766),
            .I(N__66737));
    InMux I__15920 (
            .O(N__66765),
            .I(N__66737));
    InMux I__15919 (
            .O(N__66764),
            .I(N__66730));
    InMux I__15918 (
            .O(N__66763),
            .I(N__66727));
    InMux I__15917 (
            .O(N__66762),
            .I(N__66722));
    InMux I__15916 (
            .O(N__66761),
            .I(N__66722));
    LocalMux I__15915 (
            .O(N__66758),
            .I(N__66710));
    InMux I__15914 (
            .O(N__66757),
            .I(N__66705));
    InMux I__15913 (
            .O(N__66756),
            .I(N__66705));
    CascadeMux I__15912 (
            .O(N__66755),
            .I(N__66693));
    InMux I__15911 (
            .O(N__66754),
            .I(N__66690));
    InMux I__15910 (
            .O(N__66753),
            .I(N__66687));
    LocalMux I__15909 (
            .O(N__66750),
            .I(N__66677));
    LocalMux I__15908 (
            .O(N__66747),
            .I(N__66677));
    InMux I__15907 (
            .O(N__66746),
            .I(N__66672));
    InMux I__15906 (
            .O(N__66743),
            .I(N__66672));
    InMux I__15905 (
            .O(N__66742),
            .I(N__66669));
    LocalMux I__15904 (
            .O(N__66737),
            .I(N__66666));
    InMux I__15903 (
            .O(N__66736),
            .I(N__66663));
    InMux I__15902 (
            .O(N__66735),
            .I(N__66659));
    InMux I__15901 (
            .O(N__66734),
            .I(N__66654));
    InMux I__15900 (
            .O(N__66733),
            .I(N__66654));
    LocalMux I__15899 (
            .O(N__66730),
            .I(N__66647));
    LocalMux I__15898 (
            .O(N__66727),
            .I(N__66647));
    LocalMux I__15897 (
            .O(N__66722),
            .I(N__66644));
    InMux I__15896 (
            .O(N__66721),
            .I(N__66641));
    InMux I__15895 (
            .O(N__66720),
            .I(N__66634));
    InMux I__15894 (
            .O(N__66719),
            .I(N__66634));
    InMux I__15893 (
            .O(N__66718),
            .I(N__66634));
    CascadeMux I__15892 (
            .O(N__66717),
            .I(N__66631));
    InMux I__15891 (
            .O(N__66716),
            .I(N__66626));
    InMux I__15890 (
            .O(N__66715),
            .I(N__66623));
    InMux I__15889 (
            .O(N__66714),
            .I(N__66618));
    InMux I__15888 (
            .O(N__66713),
            .I(N__66618));
    Span4Mux_h I__15887 (
            .O(N__66710),
            .I(N__66615));
    LocalMux I__15886 (
            .O(N__66705),
            .I(N__66612));
    InMux I__15885 (
            .O(N__66704),
            .I(N__66609));
    InMux I__15884 (
            .O(N__66703),
            .I(N__66604));
    InMux I__15883 (
            .O(N__66702),
            .I(N__66604));
    InMux I__15882 (
            .O(N__66701),
            .I(N__66591));
    InMux I__15881 (
            .O(N__66700),
            .I(N__66591));
    InMux I__15880 (
            .O(N__66699),
            .I(N__66586));
    InMux I__15879 (
            .O(N__66698),
            .I(N__66586));
    InMux I__15878 (
            .O(N__66697),
            .I(N__66583));
    CascadeMux I__15877 (
            .O(N__66696),
            .I(N__66574));
    InMux I__15876 (
            .O(N__66693),
            .I(N__66571));
    LocalMux I__15875 (
            .O(N__66690),
            .I(N__66564));
    LocalMux I__15874 (
            .O(N__66687),
            .I(N__66564));
    InMux I__15873 (
            .O(N__66686),
            .I(N__66559));
    InMux I__15872 (
            .O(N__66685),
            .I(N__66559));
    InMux I__15871 (
            .O(N__66684),
            .I(N__66552));
    InMux I__15870 (
            .O(N__66683),
            .I(N__66552));
    InMux I__15869 (
            .O(N__66682),
            .I(N__66552));
    Span4Mux_v I__15868 (
            .O(N__66677),
            .I(N__66547));
    LocalMux I__15867 (
            .O(N__66672),
            .I(N__66547));
    LocalMux I__15866 (
            .O(N__66669),
            .I(N__66540));
    Span4Mux_v I__15865 (
            .O(N__66666),
            .I(N__66540));
    LocalMux I__15864 (
            .O(N__66663),
            .I(N__66540));
    InMux I__15863 (
            .O(N__66662),
            .I(N__66537));
    LocalMux I__15862 (
            .O(N__66659),
            .I(N__66532));
    LocalMux I__15861 (
            .O(N__66654),
            .I(N__66532));
    InMux I__15860 (
            .O(N__66653),
            .I(N__66529));
    InMux I__15859 (
            .O(N__66652),
            .I(N__66526));
    Span4Mux_h I__15858 (
            .O(N__66647),
            .I(N__66523));
    Span4Mux_h I__15857 (
            .O(N__66644),
            .I(N__66516));
    LocalMux I__15856 (
            .O(N__66641),
            .I(N__66516));
    LocalMux I__15855 (
            .O(N__66634),
            .I(N__66516));
    InMux I__15854 (
            .O(N__66631),
            .I(N__66513));
    InMux I__15853 (
            .O(N__66630),
            .I(N__66508));
    InMux I__15852 (
            .O(N__66629),
            .I(N__66508));
    LocalMux I__15851 (
            .O(N__66626),
            .I(N__66501));
    LocalMux I__15850 (
            .O(N__66623),
            .I(N__66501));
    LocalMux I__15849 (
            .O(N__66618),
            .I(N__66501));
    Span4Mux_v I__15848 (
            .O(N__66615),
            .I(N__66492));
    Span4Mux_v I__15847 (
            .O(N__66612),
            .I(N__66492));
    LocalMux I__15846 (
            .O(N__66609),
            .I(N__66492));
    LocalMux I__15845 (
            .O(N__66604),
            .I(N__66492));
    InMux I__15844 (
            .O(N__66603),
            .I(N__66487));
    InMux I__15843 (
            .O(N__66602),
            .I(N__66487));
    InMux I__15842 (
            .O(N__66601),
            .I(N__66482));
    InMux I__15841 (
            .O(N__66600),
            .I(N__66482));
    InMux I__15840 (
            .O(N__66599),
            .I(N__66473));
    InMux I__15839 (
            .O(N__66598),
            .I(N__66473));
    InMux I__15838 (
            .O(N__66597),
            .I(N__66473));
    InMux I__15837 (
            .O(N__66596),
            .I(N__66473));
    LocalMux I__15836 (
            .O(N__66591),
            .I(N__66468));
    LocalMux I__15835 (
            .O(N__66586),
            .I(N__66468));
    LocalMux I__15834 (
            .O(N__66583),
            .I(N__66465));
    InMux I__15833 (
            .O(N__66582),
            .I(N__66462));
    InMux I__15832 (
            .O(N__66581),
            .I(N__66451));
    InMux I__15831 (
            .O(N__66580),
            .I(N__66451));
    InMux I__15830 (
            .O(N__66579),
            .I(N__66451));
    InMux I__15829 (
            .O(N__66578),
            .I(N__66451));
    InMux I__15828 (
            .O(N__66577),
            .I(N__66451));
    InMux I__15827 (
            .O(N__66574),
            .I(N__66448));
    LocalMux I__15826 (
            .O(N__66571),
            .I(N__66445));
    InMux I__15825 (
            .O(N__66570),
            .I(N__66442));
    InMux I__15824 (
            .O(N__66569),
            .I(N__66438));
    Span4Mux_v I__15823 (
            .O(N__66564),
            .I(N__66435));
    LocalMux I__15822 (
            .O(N__66559),
            .I(N__66426));
    LocalMux I__15821 (
            .O(N__66552),
            .I(N__66426));
    Span4Mux_v I__15820 (
            .O(N__66547),
            .I(N__66426));
    Span4Mux_h I__15819 (
            .O(N__66540),
            .I(N__66426));
    LocalMux I__15818 (
            .O(N__66537),
            .I(N__66421));
    Span4Mux_v I__15817 (
            .O(N__66532),
            .I(N__66421));
    LocalMux I__15816 (
            .O(N__66529),
            .I(N__66418));
    LocalMux I__15815 (
            .O(N__66526),
            .I(N__66415));
    Span4Mux_v I__15814 (
            .O(N__66523),
            .I(N__66410));
    Span4Mux_h I__15813 (
            .O(N__66516),
            .I(N__66410));
    LocalMux I__15812 (
            .O(N__66513),
            .I(N__66401));
    LocalMux I__15811 (
            .O(N__66508),
            .I(N__66401));
    Span4Mux_v I__15810 (
            .O(N__66501),
            .I(N__66401));
    Span4Mux_h I__15809 (
            .O(N__66492),
            .I(N__66401));
    LocalMux I__15808 (
            .O(N__66487),
            .I(N__66394));
    LocalMux I__15807 (
            .O(N__66482),
            .I(N__66394));
    LocalMux I__15806 (
            .O(N__66473),
            .I(N__66394));
    Span4Mux_h I__15805 (
            .O(N__66468),
            .I(N__66385));
    Span4Mux_v I__15804 (
            .O(N__66465),
            .I(N__66385));
    LocalMux I__15803 (
            .O(N__66462),
            .I(N__66385));
    LocalMux I__15802 (
            .O(N__66451),
            .I(N__66385));
    LocalMux I__15801 (
            .O(N__66448),
            .I(N__66378));
    Span4Mux_h I__15800 (
            .O(N__66445),
            .I(N__66378));
    LocalMux I__15799 (
            .O(N__66442),
            .I(N__66378));
    InMux I__15798 (
            .O(N__66441),
            .I(N__66372));
    LocalMux I__15797 (
            .O(N__66438),
            .I(N__66369));
    Span4Mux_v I__15796 (
            .O(N__66435),
            .I(N__66362));
    Span4Mux_h I__15795 (
            .O(N__66426),
            .I(N__66362));
    Span4Mux_v I__15794 (
            .O(N__66421),
            .I(N__66362));
    Span4Mux_v I__15793 (
            .O(N__66418),
            .I(N__66355));
    Span4Mux_v I__15792 (
            .O(N__66415),
            .I(N__66355));
    Span4Mux_h I__15791 (
            .O(N__66410),
            .I(N__66355));
    Span4Mux_h I__15790 (
            .O(N__66401),
            .I(N__66350));
    Span4Mux_v I__15789 (
            .O(N__66394),
            .I(N__66350));
    Span4Mux_h I__15788 (
            .O(N__66385),
            .I(N__66345));
    Span4Mux_v I__15787 (
            .O(N__66378),
            .I(N__66345));
    InMux I__15786 (
            .O(N__66377),
            .I(N__66340));
    InMux I__15785 (
            .O(N__66376),
            .I(N__66340));
    InMux I__15784 (
            .O(N__66375),
            .I(N__66337));
    LocalMux I__15783 (
            .O(N__66372),
            .I(\ALU.status_19 ));
    Odrv4 I__15782 (
            .O(N__66369),
            .I(\ALU.status_19 ));
    Odrv4 I__15781 (
            .O(N__66362),
            .I(\ALU.status_19 ));
    Odrv4 I__15780 (
            .O(N__66355),
            .I(\ALU.status_19 ));
    Odrv4 I__15779 (
            .O(N__66350),
            .I(\ALU.status_19 ));
    Odrv4 I__15778 (
            .O(N__66345),
            .I(\ALU.status_19 ));
    LocalMux I__15777 (
            .O(N__66340),
            .I(\ALU.status_19 ));
    LocalMux I__15776 (
            .O(N__66337),
            .I(\ALU.status_19 ));
    InMux I__15775 (
            .O(N__66320),
            .I(N__66317));
    LocalMux I__15774 (
            .O(N__66317),
            .I(N__66309));
    InMux I__15773 (
            .O(N__66316),
            .I(N__66304));
    InMux I__15772 (
            .O(N__66315),
            .I(N__66304));
    InMux I__15771 (
            .O(N__66314),
            .I(N__66300));
    InMux I__15770 (
            .O(N__66313),
            .I(N__66293));
    InMux I__15769 (
            .O(N__66312),
            .I(N__66289));
    Span4Mux_v I__15768 (
            .O(N__66309),
            .I(N__66284));
    LocalMux I__15767 (
            .O(N__66304),
            .I(N__66281));
    InMux I__15766 (
            .O(N__66303),
            .I(N__66278));
    LocalMux I__15765 (
            .O(N__66300),
            .I(N__66275));
    InMux I__15764 (
            .O(N__66299),
            .I(N__66272));
    InMux I__15763 (
            .O(N__66298),
            .I(N__66266));
    InMux I__15762 (
            .O(N__66297),
            .I(N__66263));
    InMux I__15761 (
            .O(N__66296),
            .I(N__66260));
    LocalMux I__15760 (
            .O(N__66293),
            .I(N__66257));
    InMux I__15759 (
            .O(N__66292),
            .I(N__66254));
    LocalMux I__15758 (
            .O(N__66289),
            .I(N__66245));
    InMux I__15757 (
            .O(N__66288),
            .I(N__66242));
    InMux I__15756 (
            .O(N__66287),
            .I(N__66237));
    Span4Mux_v I__15755 (
            .O(N__66284),
            .I(N__66230));
    Span4Mux_v I__15754 (
            .O(N__66281),
            .I(N__66230));
    LocalMux I__15753 (
            .O(N__66278),
            .I(N__66230));
    Span4Mux_v I__15752 (
            .O(N__66275),
            .I(N__66225));
    LocalMux I__15751 (
            .O(N__66272),
            .I(N__66222));
    InMux I__15750 (
            .O(N__66271),
            .I(N__66215));
    InMux I__15749 (
            .O(N__66270),
            .I(N__66215));
    InMux I__15748 (
            .O(N__66269),
            .I(N__66215));
    LocalMux I__15747 (
            .O(N__66266),
            .I(N__66208));
    LocalMux I__15746 (
            .O(N__66263),
            .I(N__66208));
    LocalMux I__15745 (
            .O(N__66260),
            .I(N__66208));
    Span4Mux_v I__15744 (
            .O(N__66257),
            .I(N__66203));
    LocalMux I__15743 (
            .O(N__66254),
            .I(N__66203));
    InMux I__15742 (
            .O(N__66253),
            .I(N__66198));
    InMux I__15741 (
            .O(N__66252),
            .I(N__66198));
    InMux I__15740 (
            .O(N__66251),
            .I(N__66195));
    InMux I__15739 (
            .O(N__66250),
            .I(N__66188));
    InMux I__15738 (
            .O(N__66249),
            .I(N__66188));
    InMux I__15737 (
            .O(N__66248),
            .I(N__66188));
    Span4Mux_h I__15736 (
            .O(N__66245),
            .I(N__66183));
    LocalMux I__15735 (
            .O(N__66242),
            .I(N__66183));
    InMux I__15734 (
            .O(N__66241),
            .I(N__66180));
    InMux I__15733 (
            .O(N__66240),
            .I(N__66177));
    LocalMux I__15732 (
            .O(N__66237),
            .I(N__66169));
    Span4Mux_h I__15731 (
            .O(N__66230),
            .I(N__66169));
    InMux I__15730 (
            .O(N__66229),
            .I(N__66164));
    InMux I__15729 (
            .O(N__66228),
            .I(N__66164));
    Span4Mux_h I__15728 (
            .O(N__66225),
            .I(N__66161));
    Span4Mux_v I__15727 (
            .O(N__66222),
            .I(N__66154));
    LocalMux I__15726 (
            .O(N__66215),
            .I(N__66154));
    Span4Mux_v I__15725 (
            .O(N__66208),
            .I(N__66154));
    Span4Mux_v I__15724 (
            .O(N__66203),
            .I(N__66151));
    LocalMux I__15723 (
            .O(N__66198),
            .I(N__66140));
    LocalMux I__15722 (
            .O(N__66195),
            .I(N__66140));
    LocalMux I__15721 (
            .O(N__66188),
            .I(N__66140));
    Span4Mux_v I__15720 (
            .O(N__66183),
            .I(N__66140));
    LocalMux I__15719 (
            .O(N__66180),
            .I(N__66140));
    LocalMux I__15718 (
            .O(N__66177),
            .I(N__66137));
    InMux I__15717 (
            .O(N__66176),
            .I(N__66134));
    InMux I__15716 (
            .O(N__66175),
            .I(N__66131));
    InMux I__15715 (
            .O(N__66174),
            .I(N__66128));
    Span4Mux_h I__15714 (
            .O(N__66169),
            .I(N__66124));
    LocalMux I__15713 (
            .O(N__66164),
            .I(N__66117));
    Span4Mux_h I__15712 (
            .O(N__66161),
            .I(N__66117));
    Span4Mux_h I__15711 (
            .O(N__66154),
            .I(N__66117));
    Span4Mux_h I__15710 (
            .O(N__66151),
            .I(N__66112));
    Span4Mux_v I__15709 (
            .O(N__66140),
            .I(N__66112));
    Span12Mux_h I__15708 (
            .O(N__66137),
            .I(N__66103));
    LocalMux I__15707 (
            .O(N__66134),
            .I(N__66103));
    LocalMux I__15706 (
            .O(N__66131),
            .I(N__66103));
    LocalMux I__15705 (
            .O(N__66128),
            .I(N__66103));
    InMux I__15704 (
            .O(N__66127),
            .I(N__66100));
    Odrv4 I__15703 (
            .O(N__66124),
            .I(aluOut_2));
    Odrv4 I__15702 (
            .O(N__66117),
            .I(aluOut_2));
    Odrv4 I__15701 (
            .O(N__66112),
            .I(aluOut_2));
    Odrv12 I__15700 (
            .O(N__66103),
            .I(aluOut_2));
    LocalMux I__15699 (
            .O(N__66100),
            .I(aluOut_2));
    CascadeMux I__15698 (
            .O(N__66089),
            .I(N__66086));
    InMux I__15697 (
            .O(N__66086),
            .I(N__66068));
    InMux I__15696 (
            .O(N__66085),
            .I(N__66068));
    InMux I__15695 (
            .O(N__66084),
            .I(N__66055));
    CascadeMux I__15694 (
            .O(N__66083),
            .I(N__66052));
    InMux I__15693 (
            .O(N__66082),
            .I(N__66040));
    InMux I__15692 (
            .O(N__66081),
            .I(N__66040));
    InMux I__15691 (
            .O(N__66080),
            .I(N__66037));
    InMux I__15690 (
            .O(N__66079),
            .I(N__66030));
    InMux I__15689 (
            .O(N__66078),
            .I(N__66030));
    InMux I__15688 (
            .O(N__66077),
            .I(N__66030));
    InMux I__15687 (
            .O(N__66076),
            .I(N__66023));
    InMux I__15686 (
            .O(N__66075),
            .I(N__66020));
    InMux I__15685 (
            .O(N__66074),
            .I(N__66015));
    InMux I__15684 (
            .O(N__66073),
            .I(N__66015));
    LocalMux I__15683 (
            .O(N__66068),
            .I(N__66007));
    InMux I__15682 (
            .O(N__66067),
            .I(N__66000));
    InMux I__15681 (
            .O(N__66066),
            .I(N__66000));
    InMux I__15680 (
            .O(N__66065),
            .I(N__66000));
    InMux I__15679 (
            .O(N__66064),
            .I(N__65991));
    InMux I__15678 (
            .O(N__66063),
            .I(N__65991));
    InMux I__15677 (
            .O(N__66062),
            .I(N__65991));
    InMux I__15676 (
            .O(N__66061),
            .I(N__65991));
    InMux I__15675 (
            .O(N__66060),
            .I(N__65986));
    InMux I__15674 (
            .O(N__66059),
            .I(N__65981));
    InMux I__15673 (
            .O(N__66058),
            .I(N__65981));
    LocalMux I__15672 (
            .O(N__66055),
            .I(N__65978));
    InMux I__15671 (
            .O(N__66052),
            .I(N__65969));
    InMux I__15670 (
            .O(N__66051),
            .I(N__65969));
    InMux I__15669 (
            .O(N__66050),
            .I(N__65969));
    InMux I__15668 (
            .O(N__66049),
            .I(N__65969));
    InMux I__15667 (
            .O(N__66048),
            .I(N__65959));
    InMux I__15666 (
            .O(N__66047),
            .I(N__65944));
    InMux I__15665 (
            .O(N__66046),
            .I(N__65944));
    InMux I__15664 (
            .O(N__66045),
            .I(N__65944));
    LocalMux I__15663 (
            .O(N__66040),
            .I(N__65937));
    LocalMux I__15662 (
            .O(N__66037),
            .I(N__65937));
    LocalMux I__15661 (
            .O(N__66030),
            .I(N__65937));
    CascadeMux I__15660 (
            .O(N__66029),
            .I(N__65932));
    InMux I__15659 (
            .O(N__66028),
            .I(N__65921));
    InMux I__15658 (
            .O(N__66027),
            .I(N__65921));
    InMux I__15657 (
            .O(N__66026),
            .I(N__65918));
    LocalMux I__15656 (
            .O(N__66023),
            .I(N__65911));
    LocalMux I__15655 (
            .O(N__66020),
            .I(N__65911));
    LocalMux I__15654 (
            .O(N__66015),
            .I(N__65911));
    InMux I__15653 (
            .O(N__66014),
            .I(N__65906));
    InMux I__15652 (
            .O(N__66013),
            .I(N__65906));
    InMux I__15651 (
            .O(N__66012),
            .I(N__65899));
    InMux I__15650 (
            .O(N__66011),
            .I(N__65896));
    InMux I__15649 (
            .O(N__66010),
            .I(N__65893));
    Span4Mux_v I__15648 (
            .O(N__66007),
            .I(N__65890));
    LocalMux I__15647 (
            .O(N__66000),
            .I(N__65887));
    LocalMux I__15646 (
            .O(N__65991),
            .I(N__65884));
    InMux I__15645 (
            .O(N__65990),
            .I(N__65881));
    InMux I__15644 (
            .O(N__65989),
            .I(N__65878));
    LocalMux I__15643 (
            .O(N__65986),
            .I(N__65873));
    LocalMux I__15642 (
            .O(N__65981),
            .I(N__65873));
    Span4Mux_h I__15641 (
            .O(N__65978),
            .I(N__65868));
    LocalMux I__15640 (
            .O(N__65969),
            .I(N__65868));
    InMux I__15639 (
            .O(N__65968),
            .I(N__65861));
    InMux I__15638 (
            .O(N__65967),
            .I(N__65861));
    InMux I__15637 (
            .O(N__65966),
            .I(N__65861));
    InMux I__15636 (
            .O(N__65965),
            .I(N__65852));
    InMux I__15635 (
            .O(N__65964),
            .I(N__65852));
    InMux I__15634 (
            .O(N__65963),
            .I(N__65852));
    InMux I__15633 (
            .O(N__65962),
            .I(N__65852));
    LocalMux I__15632 (
            .O(N__65959),
            .I(N__65849));
    InMux I__15631 (
            .O(N__65958),
            .I(N__65840));
    InMux I__15630 (
            .O(N__65957),
            .I(N__65840));
    InMux I__15629 (
            .O(N__65956),
            .I(N__65840));
    InMux I__15628 (
            .O(N__65955),
            .I(N__65840));
    InMux I__15627 (
            .O(N__65954),
            .I(N__65837));
    InMux I__15626 (
            .O(N__65953),
            .I(N__65834));
    InMux I__15625 (
            .O(N__65952),
            .I(N__65829));
    InMux I__15624 (
            .O(N__65951),
            .I(N__65829));
    LocalMux I__15623 (
            .O(N__65944),
            .I(N__65823));
    Span4Mux_v I__15622 (
            .O(N__65937),
            .I(N__65820));
    InMux I__15621 (
            .O(N__65936),
            .I(N__65817));
    InMux I__15620 (
            .O(N__65935),
            .I(N__65814));
    InMux I__15619 (
            .O(N__65932),
            .I(N__65811));
    InMux I__15618 (
            .O(N__65931),
            .I(N__65808));
    InMux I__15617 (
            .O(N__65930),
            .I(N__65805));
    InMux I__15616 (
            .O(N__65929),
            .I(N__65802));
    CascadeMux I__15615 (
            .O(N__65928),
            .I(N__65799));
    InMux I__15614 (
            .O(N__65927),
            .I(N__65794));
    InMux I__15613 (
            .O(N__65926),
            .I(N__65794));
    LocalMux I__15612 (
            .O(N__65921),
            .I(N__65789));
    LocalMux I__15611 (
            .O(N__65918),
            .I(N__65789));
    Span4Mux_v I__15610 (
            .O(N__65911),
            .I(N__65784));
    LocalMux I__15609 (
            .O(N__65906),
            .I(N__65784));
    InMux I__15608 (
            .O(N__65905),
            .I(N__65779));
    InMux I__15607 (
            .O(N__65904),
            .I(N__65779));
    InMux I__15606 (
            .O(N__65903),
            .I(N__65774));
    InMux I__15605 (
            .O(N__65902),
            .I(N__65774));
    LocalMux I__15604 (
            .O(N__65899),
            .I(N__65771));
    LocalMux I__15603 (
            .O(N__65896),
            .I(N__65766));
    LocalMux I__15602 (
            .O(N__65893),
            .I(N__65766));
    Span4Mux_h I__15601 (
            .O(N__65890),
            .I(N__65759));
    Span4Mux_v I__15600 (
            .O(N__65887),
            .I(N__65759));
    Span4Mux_v I__15599 (
            .O(N__65884),
            .I(N__65759));
    LocalMux I__15598 (
            .O(N__65881),
            .I(N__65756));
    LocalMux I__15597 (
            .O(N__65878),
            .I(N__65750));
    Span4Mux_h I__15596 (
            .O(N__65873),
            .I(N__65743));
    Span4Mux_v I__15595 (
            .O(N__65868),
            .I(N__65743));
    LocalMux I__15594 (
            .O(N__65861),
            .I(N__65743));
    LocalMux I__15593 (
            .O(N__65852),
            .I(N__65740));
    Span4Mux_h I__15592 (
            .O(N__65849),
            .I(N__65737));
    LocalMux I__15591 (
            .O(N__65840),
            .I(N__65734));
    LocalMux I__15590 (
            .O(N__65837),
            .I(N__65727));
    LocalMux I__15589 (
            .O(N__65834),
            .I(N__65727));
    LocalMux I__15588 (
            .O(N__65829),
            .I(N__65727));
    InMux I__15587 (
            .O(N__65828),
            .I(N__65724));
    CascadeMux I__15586 (
            .O(N__65827),
            .I(N__65721));
    CascadeMux I__15585 (
            .O(N__65826),
            .I(N__65712));
    Span4Mux_v I__15584 (
            .O(N__65823),
            .I(N__65701));
    Span4Mux_h I__15583 (
            .O(N__65820),
            .I(N__65701));
    LocalMux I__15582 (
            .O(N__65817),
            .I(N__65701));
    LocalMux I__15581 (
            .O(N__65814),
            .I(N__65701));
    LocalMux I__15580 (
            .O(N__65811),
            .I(N__65698));
    LocalMux I__15579 (
            .O(N__65808),
            .I(N__65695));
    LocalMux I__15578 (
            .O(N__65805),
            .I(N__65690));
    LocalMux I__15577 (
            .O(N__65802),
            .I(N__65690));
    InMux I__15576 (
            .O(N__65799),
            .I(N__65687));
    LocalMux I__15575 (
            .O(N__65794),
            .I(N__65676));
    Span4Mux_v I__15574 (
            .O(N__65789),
            .I(N__65676));
    Span4Mux_h I__15573 (
            .O(N__65784),
            .I(N__65676));
    LocalMux I__15572 (
            .O(N__65779),
            .I(N__65676));
    LocalMux I__15571 (
            .O(N__65774),
            .I(N__65676));
    Span4Mux_v I__15570 (
            .O(N__65771),
            .I(N__65667));
    Span4Mux_v I__15569 (
            .O(N__65766),
            .I(N__65667));
    Span4Mux_h I__15568 (
            .O(N__65759),
            .I(N__65667));
    Span4Mux_v I__15567 (
            .O(N__65756),
            .I(N__65667));
    InMux I__15566 (
            .O(N__65755),
            .I(N__65660));
    InMux I__15565 (
            .O(N__65754),
            .I(N__65660));
    InMux I__15564 (
            .O(N__65753),
            .I(N__65660));
    Span4Mux_v I__15563 (
            .O(N__65750),
            .I(N__65655));
    Span4Mux_h I__15562 (
            .O(N__65743),
            .I(N__65655));
    Span4Mux_v I__15561 (
            .O(N__65740),
            .I(N__65652));
    Span4Mux_h I__15560 (
            .O(N__65737),
            .I(N__65647));
    Span4Mux_h I__15559 (
            .O(N__65734),
            .I(N__65647));
    Span4Mux_h I__15558 (
            .O(N__65727),
            .I(N__65642));
    LocalMux I__15557 (
            .O(N__65724),
            .I(N__65642));
    InMux I__15556 (
            .O(N__65721),
            .I(N__65635));
    InMux I__15555 (
            .O(N__65720),
            .I(N__65635));
    InMux I__15554 (
            .O(N__65719),
            .I(N__65635));
    InMux I__15553 (
            .O(N__65718),
            .I(N__65628));
    InMux I__15552 (
            .O(N__65717),
            .I(N__65628));
    InMux I__15551 (
            .O(N__65716),
            .I(N__65628));
    InMux I__15550 (
            .O(N__65715),
            .I(N__65619));
    InMux I__15549 (
            .O(N__65712),
            .I(N__65619));
    InMux I__15548 (
            .O(N__65711),
            .I(N__65619));
    InMux I__15547 (
            .O(N__65710),
            .I(N__65619));
    Span4Mux_h I__15546 (
            .O(N__65701),
            .I(N__65610));
    Span4Mux_v I__15545 (
            .O(N__65698),
            .I(N__65610));
    Span4Mux_v I__15544 (
            .O(N__65695),
            .I(N__65610));
    Span4Mux_h I__15543 (
            .O(N__65690),
            .I(N__65610));
    LocalMux I__15542 (
            .O(N__65687),
            .I(\ALU.status_19_0 ));
    Odrv4 I__15541 (
            .O(N__65676),
            .I(\ALU.status_19_0 ));
    Odrv4 I__15540 (
            .O(N__65667),
            .I(\ALU.status_19_0 ));
    LocalMux I__15539 (
            .O(N__65660),
            .I(\ALU.status_19_0 ));
    Odrv4 I__15538 (
            .O(N__65655),
            .I(\ALU.status_19_0 ));
    Odrv4 I__15537 (
            .O(N__65652),
            .I(\ALU.status_19_0 ));
    Odrv4 I__15536 (
            .O(N__65647),
            .I(\ALU.status_19_0 ));
    Odrv4 I__15535 (
            .O(N__65642),
            .I(\ALU.status_19_0 ));
    LocalMux I__15534 (
            .O(N__65635),
            .I(\ALU.status_19_0 ));
    LocalMux I__15533 (
            .O(N__65628),
            .I(\ALU.status_19_0 ));
    LocalMux I__15532 (
            .O(N__65619),
            .I(\ALU.status_19_0 ));
    Odrv4 I__15531 (
            .O(N__65610),
            .I(\ALU.status_19_0 ));
    CascadeMux I__15530 (
            .O(N__65585),
            .I(N__65581));
    InMux I__15529 (
            .O(N__65584),
            .I(N__65576));
    InMux I__15528 (
            .O(N__65581),
            .I(N__65576));
    LocalMux I__15527 (
            .O(N__65576),
            .I(N__65571));
    CascadeMux I__15526 (
            .O(N__65575),
            .I(N__65566));
    CascadeMux I__15525 (
            .O(N__65574),
            .I(N__65559));
    Span4Mux_v I__15524 (
            .O(N__65571),
            .I(N__65553));
    InMux I__15523 (
            .O(N__65570),
            .I(N__65547));
    InMux I__15522 (
            .O(N__65569),
            .I(N__65531));
    InMux I__15521 (
            .O(N__65566),
            .I(N__65531));
    InMux I__15520 (
            .O(N__65565),
            .I(N__65528));
    CascadeMux I__15519 (
            .O(N__65564),
            .I(N__65523));
    InMux I__15518 (
            .O(N__65563),
            .I(N__65517));
    InMux I__15517 (
            .O(N__65562),
            .I(N__65514));
    InMux I__15516 (
            .O(N__65559),
            .I(N__65511));
    InMux I__15515 (
            .O(N__65558),
            .I(N__65508));
    InMux I__15514 (
            .O(N__65557),
            .I(N__65505));
    InMux I__15513 (
            .O(N__65556),
            .I(N__65502));
    Span4Mux_h I__15512 (
            .O(N__65553),
            .I(N__65499));
    InMux I__15511 (
            .O(N__65552),
            .I(N__65494));
    InMux I__15510 (
            .O(N__65551),
            .I(N__65494));
    InMux I__15509 (
            .O(N__65550),
            .I(N__65490));
    LocalMux I__15508 (
            .O(N__65547),
            .I(N__65487));
    CascadeMux I__15507 (
            .O(N__65546),
            .I(N__65484));
    InMux I__15506 (
            .O(N__65545),
            .I(N__65474));
    InMux I__15505 (
            .O(N__65544),
            .I(N__65474));
    InMux I__15504 (
            .O(N__65543),
            .I(N__65469));
    InMux I__15503 (
            .O(N__65542),
            .I(N__65469));
    InMux I__15502 (
            .O(N__65541),
            .I(N__65464));
    InMux I__15501 (
            .O(N__65540),
            .I(N__65464));
    InMux I__15500 (
            .O(N__65539),
            .I(N__65461));
    InMux I__15499 (
            .O(N__65538),
            .I(N__65458));
    InMux I__15498 (
            .O(N__65537),
            .I(N__65455));
    InMux I__15497 (
            .O(N__65536),
            .I(N__65452));
    LocalMux I__15496 (
            .O(N__65531),
            .I(N__65447));
    LocalMux I__15495 (
            .O(N__65528),
            .I(N__65447));
    InMux I__15494 (
            .O(N__65527),
            .I(N__65439));
    InMux I__15493 (
            .O(N__65526),
            .I(N__65439));
    InMux I__15492 (
            .O(N__65523),
            .I(N__65434));
    InMux I__15491 (
            .O(N__65522),
            .I(N__65434));
    InMux I__15490 (
            .O(N__65521),
            .I(N__65431));
    InMux I__15489 (
            .O(N__65520),
            .I(N__65428));
    LocalMux I__15488 (
            .O(N__65517),
            .I(N__65423));
    LocalMux I__15487 (
            .O(N__65514),
            .I(N__65423));
    LocalMux I__15486 (
            .O(N__65511),
            .I(N__65418));
    LocalMux I__15485 (
            .O(N__65508),
            .I(N__65418));
    LocalMux I__15484 (
            .O(N__65505),
            .I(N__65409));
    LocalMux I__15483 (
            .O(N__65502),
            .I(N__65409));
    Span4Mux_v I__15482 (
            .O(N__65499),
            .I(N__65409));
    LocalMux I__15481 (
            .O(N__65494),
            .I(N__65409));
    InMux I__15480 (
            .O(N__65493),
            .I(N__65404));
    LocalMux I__15479 (
            .O(N__65490),
            .I(N__65399));
    Span4Mux_h I__15478 (
            .O(N__65487),
            .I(N__65399));
    InMux I__15477 (
            .O(N__65484),
            .I(N__65386));
    InMux I__15476 (
            .O(N__65483),
            .I(N__65386));
    InMux I__15475 (
            .O(N__65482),
            .I(N__65386));
    InMux I__15474 (
            .O(N__65481),
            .I(N__65386));
    InMux I__15473 (
            .O(N__65480),
            .I(N__65386));
    InMux I__15472 (
            .O(N__65479),
            .I(N__65386));
    LocalMux I__15471 (
            .O(N__65474),
            .I(N__65379));
    LocalMux I__15470 (
            .O(N__65469),
            .I(N__65379));
    LocalMux I__15469 (
            .O(N__65464),
            .I(N__65379));
    LocalMux I__15468 (
            .O(N__65461),
            .I(N__65374));
    LocalMux I__15467 (
            .O(N__65458),
            .I(N__65374));
    LocalMux I__15466 (
            .O(N__65455),
            .I(N__65369));
    LocalMux I__15465 (
            .O(N__65452),
            .I(N__65369));
    Span4Mux_v I__15464 (
            .O(N__65447),
            .I(N__65366));
    InMux I__15463 (
            .O(N__65446),
            .I(N__65359));
    InMux I__15462 (
            .O(N__65445),
            .I(N__65359));
    InMux I__15461 (
            .O(N__65444),
            .I(N__65359));
    LocalMux I__15460 (
            .O(N__65439),
            .I(N__65352));
    LocalMux I__15459 (
            .O(N__65434),
            .I(N__65352));
    LocalMux I__15458 (
            .O(N__65431),
            .I(N__65352));
    LocalMux I__15457 (
            .O(N__65428),
            .I(N__65348));
    Span4Mux_v I__15456 (
            .O(N__65423),
            .I(N__65343));
    Span4Mux_v I__15455 (
            .O(N__65418),
            .I(N__65343));
    Span4Mux_h I__15454 (
            .O(N__65409),
            .I(N__65340));
    InMux I__15453 (
            .O(N__65408),
            .I(N__65335));
    InMux I__15452 (
            .O(N__65407),
            .I(N__65335));
    LocalMux I__15451 (
            .O(N__65404),
            .I(N__65326));
    Span4Mux_v I__15450 (
            .O(N__65399),
            .I(N__65326));
    LocalMux I__15449 (
            .O(N__65386),
            .I(N__65326));
    Span4Mux_h I__15448 (
            .O(N__65379),
            .I(N__65326));
    Span12Mux_v I__15447 (
            .O(N__65374),
            .I(N__65319));
    Span12Mux_v I__15446 (
            .O(N__65369),
            .I(N__65319));
    Sp12to4 I__15445 (
            .O(N__65366),
            .I(N__65319));
    LocalMux I__15444 (
            .O(N__65359),
            .I(N__65316));
    Span4Mux_v I__15443 (
            .O(N__65352),
            .I(N__65313));
    InMux I__15442 (
            .O(N__65351),
            .I(N__65310));
    Span4Mux_v I__15441 (
            .O(N__65348),
            .I(N__65305));
    Span4Mux_h I__15440 (
            .O(N__65343),
            .I(N__65305));
    Span4Mux_v I__15439 (
            .O(N__65340),
            .I(N__65298));
    LocalMux I__15438 (
            .O(N__65335),
            .I(N__65298));
    Span4Mux_v I__15437 (
            .O(N__65326),
            .I(N__65298));
    Odrv12 I__15436 (
            .O(N__65319),
            .I(aluOut_1));
    Odrv12 I__15435 (
            .O(N__65316),
            .I(aluOut_1));
    Odrv4 I__15434 (
            .O(N__65313),
            .I(aluOut_1));
    LocalMux I__15433 (
            .O(N__65310),
            .I(aluOut_1));
    Odrv4 I__15432 (
            .O(N__65305),
            .I(aluOut_1));
    Odrv4 I__15431 (
            .O(N__65298),
            .I(aluOut_1));
    InMux I__15430 (
            .O(N__65285),
            .I(N__65282));
    LocalMux I__15429 (
            .O(N__65282),
            .I(\ALU.d_RNIMGKJC1_0Z0Z_2 ));
    CascadeMux I__15428 (
            .O(N__65279),
            .I(\ALU.d_RNIMGKJC1Z0Z_2_cascade_ ));
    InMux I__15427 (
            .O(N__65276),
            .I(N__65273));
    LocalMux I__15426 (
            .O(N__65273),
            .I(N__65269));
    InMux I__15425 (
            .O(N__65272),
            .I(N__65266));
    Span4Mux_v I__15424 (
            .O(N__65269),
            .I(N__65263));
    LocalMux I__15423 (
            .O(N__65266),
            .I(N__65260));
    Sp12to4 I__15422 (
            .O(N__65263),
            .I(N__65255));
    Span12Mux_s9_h I__15421 (
            .O(N__65260),
            .I(N__65255));
    Span12Mux_h I__15420 (
            .O(N__65255),
            .I(N__65252));
    Odrv12 I__15419 (
            .O(N__65252),
            .I(\ALU.N_831 ));
    InMux I__15418 (
            .O(N__65249),
            .I(N__65246));
    LocalMux I__15417 (
            .O(N__65246),
            .I(N__65243));
    Odrv4 I__15416 (
            .O(N__65243),
            .I(\PROM.ROMDATA.m427_bm ));
    CascadeMux I__15415 (
            .O(N__65240),
            .I(\PROM.ROMDATA.m427_am_cascade_ ));
    CascadeMux I__15414 (
            .O(N__65237),
            .I(N__65233));
    InMux I__15413 (
            .O(N__65236),
            .I(N__65228));
    InMux I__15412 (
            .O(N__65233),
            .I(N__65228));
    LocalMux I__15411 (
            .O(N__65228),
            .I(N__65225));
    Span4Mux_v I__15410 (
            .O(N__65225),
            .I(N__65222));
    Sp12to4 I__15409 (
            .O(N__65222),
            .I(N__65219));
    Span12Mux_h I__15408 (
            .O(N__65219),
            .I(N__65216));
    Odrv12 I__15407 (
            .O(N__65216),
            .I(\PROM.ROMDATA.m427_ns ));
    InMux I__15406 (
            .O(N__65213),
            .I(N__65210));
    LocalMux I__15405 (
            .O(N__65210),
            .I(N__65207));
    Span4Mux_h I__15404 (
            .O(N__65207),
            .I(N__65204));
    Odrv4 I__15403 (
            .O(N__65204),
            .I(\PROM.ROMDATA.m492_am ));
    CascadeMux I__15402 (
            .O(N__65201),
            .I(N__65198));
    InMux I__15401 (
            .O(N__65198),
            .I(N__65195));
    LocalMux I__15400 (
            .O(N__65195),
            .I(\PROM.ROMDATA.m492_bm ));
    InMux I__15399 (
            .O(N__65192),
            .I(N__65189));
    LocalMux I__15398 (
            .O(N__65189),
            .I(N__65186));
    Odrv12 I__15397 (
            .O(N__65186),
            .I(\PROM.ROMDATA.m494_ns_1 ));
    InMux I__15396 (
            .O(N__65183),
            .I(N__65180));
    LocalMux I__15395 (
            .O(N__65180),
            .I(N__65177));
    Span4Mux_h I__15394 (
            .O(N__65177),
            .I(N__65174));
    Odrv4 I__15393 (
            .O(N__65174),
            .I(\PROM.ROMDATA.m88 ));
    InMux I__15392 (
            .O(N__65171),
            .I(N__65168));
    LocalMux I__15391 (
            .O(N__65168),
            .I(N__65165));
    Span4Mux_v I__15390 (
            .O(N__65165),
            .I(N__65162));
    Sp12to4 I__15389 (
            .O(N__65162),
            .I(N__65159));
    Span12Mux_h I__15388 (
            .O(N__65159),
            .I(N__65156));
    Odrv12 I__15387 (
            .O(N__65156),
            .I(\PROM.ROMDATA.m514_ns_1 ));
    CascadeMux I__15386 (
            .O(N__65153),
            .I(\PROM.ROMDATA.m181_cascade_ ));
    InMux I__15385 (
            .O(N__65150),
            .I(N__65146));
    CascadeMux I__15384 (
            .O(N__65149),
            .I(N__65143));
    LocalMux I__15383 (
            .O(N__65146),
            .I(N__65140));
    InMux I__15382 (
            .O(N__65143),
            .I(N__65137));
    Span4Mux_v I__15381 (
            .O(N__65140),
            .I(N__65134));
    LocalMux I__15380 (
            .O(N__65137),
            .I(N__65131));
    Span4Mux_v I__15379 (
            .O(N__65134),
            .I(N__65126));
    Span4Mux_h I__15378 (
            .O(N__65131),
            .I(N__65126));
    Span4Mux_h I__15377 (
            .O(N__65126),
            .I(N__65123));
    Span4Mux_v I__15376 (
            .O(N__65123),
            .I(N__65120));
    Span4Mux_h I__15375 (
            .O(N__65120),
            .I(N__65117));
    Odrv4 I__15374 (
            .O(N__65117),
            .I(\PROM.ROMDATA.m514_ns ));
    InMux I__15373 (
            .O(N__65114),
            .I(N__65111));
    LocalMux I__15372 (
            .O(N__65111),
            .I(\PROM.ROMDATA.N_525_mux ));
    InMux I__15371 (
            .O(N__65108),
            .I(N__65105));
    LocalMux I__15370 (
            .O(N__65105),
            .I(\PROM.ROMDATA.m164 ));
    InMux I__15369 (
            .O(N__65102),
            .I(N__65099));
    LocalMux I__15368 (
            .O(N__65099),
            .I(\PROM.ROMDATA.m171_am ));
    InMux I__15367 (
            .O(N__65096),
            .I(N__65093));
    LocalMux I__15366 (
            .O(N__65093),
            .I(N__65090));
    Span4Mux_v I__15365 (
            .O(N__65090),
            .I(N__65086));
    InMux I__15364 (
            .O(N__65089),
            .I(N__65083));
    Span4Mux_h I__15363 (
            .O(N__65086),
            .I(N__65078));
    LocalMux I__15362 (
            .O(N__65083),
            .I(N__65078));
    Span4Mux_v I__15361 (
            .O(N__65078),
            .I(N__65075));
    Span4Mux_h I__15360 (
            .O(N__65075),
            .I(N__65072));
    Span4Mux_h I__15359 (
            .O(N__65072),
            .I(N__65069));
    Span4Mux_h I__15358 (
            .O(N__65069),
            .I(N__65066));
    Span4Mux_v I__15357 (
            .O(N__65066),
            .I(N__65063));
    Odrv4 I__15356 (
            .O(N__65063),
            .I(\ALU.dZ0Z_12 ));
    InMux I__15355 (
            .O(N__65060),
            .I(N__65057));
    LocalMux I__15354 (
            .O(N__65057),
            .I(N__65053));
    InMux I__15353 (
            .O(N__65056),
            .I(N__65050));
    Span4Mux_v I__15352 (
            .O(N__65053),
            .I(N__65047));
    LocalMux I__15351 (
            .O(N__65050),
            .I(N__65044));
    Span4Mux_h I__15350 (
            .O(N__65047),
            .I(N__65041));
    Span12Mux_h I__15349 (
            .O(N__65044),
            .I(N__65038));
    Odrv4 I__15348 (
            .O(N__65041),
            .I(\ALU.dZ0Z_13 ));
    Odrv12 I__15347 (
            .O(N__65038),
            .I(\ALU.dZ0Z_13 ));
    CascadeMux I__15346 (
            .O(N__65033),
            .I(N__65030));
    InMux I__15345 (
            .O(N__65030),
            .I(N__65026));
    CascadeMux I__15344 (
            .O(N__65029),
            .I(N__65023));
    LocalMux I__15343 (
            .O(N__65026),
            .I(N__65020));
    InMux I__15342 (
            .O(N__65023),
            .I(N__65017));
    Span4Mux_v I__15341 (
            .O(N__65020),
            .I(N__65014));
    LocalMux I__15340 (
            .O(N__65017),
            .I(N__65010));
    Span4Mux_h I__15339 (
            .O(N__65014),
            .I(N__65007));
    InMux I__15338 (
            .O(N__65013),
            .I(N__65004));
    Span4Mux_v I__15337 (
            .O(N__65010),
            .I(N__65001));
    Span4Mux_h I__15336 (
            .O(N__65007),
            .I(N__64998));
    LocalMux I__15335 (
            .O(N__65004),
            .I(N__64995));
    Span4Mux_h I__15334 (
            .O(N__65001),
            .I(N__64992));
    Span4Mux_h I__15333 (
            .O(N__64998),
            .I(N__64989));
    Span4Mux_v I__15332 (
            .O(N__64995),
            .I(N__64984));
    Span4Mux_h I__15331 (
            .O(N__64992),
            .I(N__64984));
    Span4Mux_h I__15330 (
            .O(N__64989),
            .I(N__64981));
    Odrv4 I__15329 (
            .O(N__64984),
            .I(\PROM.ROMDATA.m83 ));
    Odrv4 I__15328 (
            .O(N__64981),
            .I(\PROM.ROMDATA.m83 ));
    CascadeMux I__15327 (
            .O(N__64976),
            .I(\PROM.ROMDATA.m83_cascade_ ));
    InMux I__15326 (
            .O(N__64973),
            .I(N__64970));
    LocalMux I__15325 (
            .O(N__64970),
            .I(N__64967));
    Span4Mux_h I__15324 (
            .O(N__64967),
            .I(N__64961));
    InMux I__15323 (
            .O(N__64966),
            .I(N__64958));
    InMux I__15322 (
            .O(N__64965),
            .I(N__64955));
    InMux I__15321 (
            .O(N__64964),
            .I(N__64952));
    Span4Mux_h I__15320 (
            .O(N__64961),
            .I(N__64949));
    LocalMux I__15319 (
            .O(N__64958),
            .I(N__64946));
    LocalMux I__15318 (
            .O(N__64955),
            .I(N__64941));
    LocalMux I__15317 (
            .O(N__64952),
            .I(N__64941));
    Span4Mux_h I__15316 (
            .O(N__64949),
            .I(N__64933));
    Span4Mux_h I__15315 (
            .O(N__64946),
            .I(N__64933));
    Span4Mux_h I__15314 (
            .O(N__64941),
            .I(N__64933));
    InMux I__15313 (
            .O(N__64940),
            .I(N__64930));
    Odrv4 I__15312 (
            .O(N__64933),
            .I(\PROM.ROMDATA.m133 ));
    LocalMux I__15311 (
            .O(N__64930),
            .I(\PROM.ROMDATA.m133 ));
    InMux I__15310 (
            .O(N__64925),
            .I(N__64922));
    LocalMux I__15309 (
            .O(N__64922),
            .I(\PROM.ROMDATA.m161 ));
    InMux I__15308 (
            .O(N__64919),
            .I(N__64916));
    LocalMux I__15307 (
            .O(N__64916),
            .I(\PROM.ROMDATA.m15 ));
    CascadeMux I__15306 (
            .O(N__64913),
            .I(\PROM.ROMDATA.m171_ns_cascade_ ));
    InMux I__15305 (
            .O(N__64910),
            .I(N__64907));
    LocalMux I__15304 (
            .O(N__64907),
            .I(\PROM.ROMDATA.m162 ));
    InMux I__15303 (
            .O(N__64904),
            .I(N__64901));
    LocalMux I__15302 (
            .O(N__64901),
            .I(N__64897));
    InMux I__15301 (
            .O(N__64900),
            .I(N__64894));
    Span4Mux_h I__15300 (
            .O(N__64897),
            .I(N__64891));
    LocalMux I__15299 (
            .O(N__64894),
            .I(N__64888));
    Span4Mux_h I__15298 (
            .O(N__64891),
            .I(N__64885));
    Span4Mux_h I__15297 (
            .O(N__64888),
            .I(N__64882));
    Odrv4 I__15296 (
            .O(N__64885),
            .I(\PROM.ROMDATA.m172 ));
    Odrv4 I__15295 (
            .O(N__64882),
            .I(\PROM.ROMDATA.m172 ));
    InMux I__15294 (
            .O(N__64877),
            .I(N__64872));
    CascadeMux I__15293 (
            .O(N__64876),
            .I(N__64867));
    CascadeMux I__15292 (
            .O(N__64875),
            .I(N__64864));
    LocalMux I__15291 (
            .O(N__64872),
            .I(N__64858));
    CascadeMux I__15290 (
            .O(N__64871),
            .I(N__64855));
    InMux I__15289 (
            .O(N__64870),
            .I(N__64852));
    InMux I__15288 (
            .O(N__64867),
            .I(N__64849));
    InMux I__15287 (
            .O(N__64864),
            .I(N__64844));
    InMux I__15286 (
            .O(N__64863),
            .I(N__64844));
    InMux I__15285 (
            .O(N__64862),
            .I(N__64841));
    CascadeMux I__15284 (
            .O(N__64861),
            .I(N__64838));
    Span4Mux_v I__15283 (
            .O(N__64858),
            .I(N__64834));
    InMux I__15282 (
            .O(N__64855),
            .I(N__64831));
    LocalMux I__15281 (
            .O(N__64852),
            .I(N__64828));
    LocalMux I__15280 (
            .O(N__64849),
            .I(N__64825));
    LocalMux I__15279 (
            .O(N__64844),
            .I(N__64822));
    LocalMux I__15278 (
            .O(N__64841),
            .I(N__64819));
    InMux I__15277 (
            .O(N__64838),
            .I(N__64814));
    InMux I__15276 (
            .O(N__64837),
            .I(N__64814));
    Span4Mux_h I__15275 (
            .O(N__64834),
            .I(N__64809));
    LocalMux I__15274 (
            .O(N__64831),
            .I(N__64809));
    Span4Mux_v I__15273 (
            .O(N__64828),
            .I(N__64804));
    Span4Mux_h I__15272 (
            .O(N__64825),
            .I(N__64804));
    Odrv12 I__15271 (
            .O(N__64822),
            .I(\PROM.ROMDATA.m20 ));
    Odrv12 I__15270 (
            .O(N__64819),
            .I(\PROM.ROMDATA.m20 ));
    LocalMux I__15269 (
            .O(N__64814),
            .I(\PROM.ROMDATA.m20 ));
    Odrv4 I__15268 (
            .O(N__64809),
            .I(\PROM.ROMDATA.m20 ));
    Odrv4 I__15267 (
            .O(N__64804),
            .I(\PROM.ROMDATA.m20 ));
    InMux I__15266 (
            .O(N__64793),
            .I(N__64790));
    LocalMux I__15265 (
            .O(N__64790),
            .I(N__64786));
    InMux I__15264 (
            .O(N__64789),
            .I(N__64783));
    Odrv4 I__15263 (
            .O(N__64786),
            .I(\PROM.ROMDATA.m156 ));
    LocalMux I__15262 (
            .O(N__64783),
            .I(\PROM.ROMDATA.m156 ));
    InMux I__15261 (
            .O(N__64778),
            .I(N__64775));
    LocalMux I__15260 (
            .O(N__64775),
            .I(\PROM.ROMDATA.m171_bm ));
    CascadeMux I__15259 (
            .O(N__64772),
            .I(\PROM.ROMDATA.m383_cascade_ ));
    InMux I__15258 (
            .O(N__64769),
            .I(N__64766));
    LocalMux I__15257 (
            .O(N__64766),
            .I(\PROM.ROMDATA.m140 ));
    CascadeMux I__15256 (
            .O(N__64763),
            .I(\PROM.ROMDATA.m138_cascade_ ));
    CascadeMux I__15255 (
            .O(N__64760),
            .I(\PROM.ROMDATA.m80_bm_1_cascade_ ));
    InMux I__15254 (
            .O(N__64757),
            .I(N__64754));
    LocalMux I__15253 (
            .O(N__64754),
            .I(N__64751));
    Odrv4 I__15252 (
            .O(N__64751),
            .I(\PROM.ROMDATA.m80_bm ));
    InMux I__15251 (
            .O(N__64748),
            .I(N__64742));
    InMux I__15250 (
            .O(N__64747),
            .I(N__64742));
    LocalMux I__15249 (
            .O(N__64742),
            .I(N__64737));
    InMux I__15248 (
            .O(N__64741),
            .I(N__64734));
    InMux I__15247 (
            .O(N__64740),
            .I(N__64731));
    Span4Mux_h I__15246 (
            .O(N__64737),
            .I(N__64728));
    LocalMux I__15245 (
            .O(N__64734),
            .I(N__64725));
    LocalMux I__15244 (
            .O(N__64731),
            .I(N__64722));
    Odrv4 I__15243 (
            .O(N__64728),
            .I(N_417));
    Odrv4 I__15242 (
            .O(N__64725),
            .I(N_417));
    Odrv12 I__15241 (
            .O(N__64722),
            .I(N_417));
    CascadeMux I__15240 (
            .O(N__64715),
            .I(N__64712));
    InMux I__15239 (
            .O(N__64712),
            .I(N__64705));
    InMux I__15238 (
            .O(N__64711),
            .I(N__64705));
    InMux I__15237 (
            .O(N__64710),
            .I(N__64702));
    LocalMux I__15236 (
            .O(N__64705),
            .I(N__64699));
    LocalMux I__15235 (
            .O(N__64702),
            .I(N__64695));
    Span4Mux_h I__15234 (
            .O(N__64699),
            .I(N__64689));
    InMux I__15233 (
            .O(N__64698),
            .I(N__64686));
    Span4Mux_v I__15232 (
            .O(N__64695),
            .I(N__64683));
    InMux I__15231 (
            .O(N__64694),
            .I(N__64680));
    InMux I__15230 (
            .O(N__64693),
            .I(N__64675));
    InMux I__15229 (
            .O(N__64692),
            .I(N__64675));
    Odrv4 I__15228 (
            .O(N__64689),
            .I(CONTROL_addrstack_reto_2));
    LocalMux I__15227 (
            .O(N__64686),
            .I(CONTROL_addrstack_reto_2));
    Odrv4 I__15226 (
            .O(N__64683),
            .I(CONTROL_addrstack_reto_2));
    LocalMux I__15225 (
            .O(N__64680),
            .I(CONTROL_addrstack_reto_2));
    LocalMux I__15224 (
            .O(N__64675),
            .I(CONTROL_addrstack_reto_2));
    InMux I__15223 (
            .O(N__64664),
            .I(N__64659));
    InMux I__15222 (
            .O(N__64663),
            .I(N__64656));
    CascadeMux I__15221 (
            .O(N__64662),
            .I(N__64652));
    LocalMux I__15220 (
            .O(N__64659),
            .I(N__64649));
    LocalMux I__15219 (
            .O(N__64656),
            .I(N__64646));
    InMux I__15218 (
            .O(N__64655),
            .I(N__64643));
    InMux I__15217 (
            .O(N__64652),
            .I(N__64638));
    Span4Mux_v I__15216 (
            .O(N__64649),
            .I(N__64635));
    Span4Mux_v I__15215 (
            .O(N__64646),
            .I(N__64632));
    LocalMux I__15214 (
            .O(N__64643),
            .I(N__64629));
    InMux I__15213 (
            .O(N__64642),
            .I(N__64626));
    CascadeMux I__15212 (
            .O(N__64641),
            .I(N__64623));
    LocalMux I__15211 (
            .O(N__64638),
            .I(N__64620));
    Span4Mux_v I__15210 (
            .O(N__64635),
            .I(N__64616));
    Span4Mux_v I__15209 (
            .O(N__64632),
            .I(N__64611));
    Span4Mux_v I__15208 (
            .O(N__64629),
            .I(N__64611));
    LocalMux I__15207 (
            .O(N__64626),
            .I(N__64608));
    InMux I__15206 (
            .O(N__64623),
            .I(N__64605));
    Span4Mux_h I__15205 (
            .O(N__64620),
            .I(N__64602));
    InMux I__15204 (
            .O(N__64619),
            .I(N__64599));
    Span4Mux_h I__15203 (
            .O(N__64616),
            .I(N__64591));
    Span4Mux_h I__15202 (
            .O(N__64611),
            .I(N__64588));
    Span4Mux_h I__15201 (
            .O(N__64608),
            .I(N__64583));
    LocalMux I__15200 (
            .O(N__64605),
            .I(N__64583));
    Span4Mux_h I__15199 (
            .O(N__64602),
            .I(N__64580));
    LocalMux I__15198 (
            .O(N__64599),
            .I(N__64577));
    InMux I__15197 (
            .O(N__64598),
            .I(N__64574));
    InMux I__15196 (
            .O(N__64597),
            .I(N__64569));
    InMux I__15195 (
            .O(N__64596),
            .I(N__64569));
    InMux I__15194 (
            .O(N__64595),
            .I(N__64566));
    InMux I__15193 (
            .O(N__64594),
            .I(N__64563));
    Odrv4 I__15192 (
            .O(N__64591),
            .I(CONTROL_programCounter11_reto_rep2));
    Odrv4 I__15191 (
            .O(N__64588),
            .I(CONTROL_programCounter11_reto_rep2));
    Odrv4 I__15190 (
            .O(N__64583),
            .I(CONTROL_programCounter11_reto_rep2));
    Odrv4 I__15189 (
            .O(N__64580),
            .I(CONTROL_programCounter11_reto_rep2));
    Odrv12 I__15188 (
            .O(N__64577),
            .I(CONTROL_programCounter11_reto_rep2));
    LocalMux I__15187 (
            .O(N__64574),
            .I(CONTROL_programCounter11_reto_rep2));
    LocalMux I__15186 (
            .O(N__64569),
            .I(CONTROL_programCounter11_reto_rep2));
    LocalMux I__15185 (
            .O(N__64566),
            .I(CONTROL_programCounter11_reto_rep2));
    LocalMux I__15184 (
            .O(N__64563),
            .I(CONTROL_programCounter11_reto_rep2));
    InMux I__15183 (
            .O(N__64544),
            .I(N__64541));
    LocalMux I__15182 (
            .O(N__64541),
            .I(\PROM.ROMDATA.m135 ));
    InMux I__15181 (
            .O(N__64538),
            .I(N__64535));
    LocalMux I__15180 (
            .O(N__64535),
            .I(\PROM.ROMDATA.m132 ));
    InMux I__15179 (
            .O(N__64532),
            .I(N__64528));
    CascadeMux I__15178 (
            .O(N__64531),
            .I(N__64525));
    LocalMux I__15177 (
            .O(N__64528),
            .I(N__64521));
    InMux I__15176 (
            .O(N__64525),
            .I(N__64518));
    InMux I__15175 (
            .O(N__64524),
            .I(N__64515));
    Span4Mux_v I__15174 (
            .O(N__64521),
            .I(N__64512));
    LocalMux I__15173 (
            .O(N__64518),
            .I(N__64509));
    LocalMux I__15172 (
            .O(N__64515),
            .I(N__64506));
    Span4Mux_h I__15171 (
            .O(N__64512),
            .I(N__64503));
    Span4Mux_v I__15170 (
            .O(N__64509),
            .I(N__64500));
    Span4Mux_h I__15169 (
            .O(N__64506),
            .I(N__64497));
    Span4Mux_h I__15168 (
            .O(N__64503),
            .I(N__64492));
    Span4Mux_h I__15167 (
            .O(N__64500),
            .I(N__64492));
    Odrv4 I__15166 (
            .O(N__64497),
            .I(N_418));
    Odrv4 I__15165 (
            .O(N__64492),
            .I(N_418));
    InMux I__15164 (
            .O(N__64487),
            .I(N__64482));
    InMux I__15163 (
            .O(N__64486),
            .I(N__64479));
    InMux I__15162 (
            .O(N__64485),
            .I(N__64476));
    LocalMux I__15161 (
            .O(N__64482),
            .I(N__64473));
    LocalMux I__15160 (
            .O(N__64479),
            .I(N__64470));
    LocalMux I__15159 (
            .O(N__64476),
            .I(N__64467));
    Span12Mux_s11_v I__15158 (
            .O(N__64473),
            .I(N__64462));
    Span4Mux_h I__15157 (
            .O(N__64470),
            .I(N__64459));
    Span4Mux_h I__15156 (
            .O(N__64467),
            .I(N__64456));
    InMux I__15155 (
            .O(N__64466),
            .I(N__64451));
    InMux I__15154 (
            .O(N__64465),
            .I(N__64451));
    Odrv12 I__15153 (
            .O(N__64462),
            .I(CONTROL_addrstack_reto_3));
    Odrv4 I__15152 (
            .O(N__64459),
            .I(CONTROL_addrstack_reto_3));
    Odrv4 I__15151 (
            .O(N__64456),
            .I(CONTROL_addrstack_reto_3));
    LocalMux I__15150 (
            .O(N__64451),
            .I(CONTROL_addrstack_reto_3));
    CascadeMux I__15149 (
            .O(N__64442),
            .I(N__64439));
    InMux I__15148 (
            .O(N__64439),
            .I(N__64436));
    LocalMux I__15147 (
            .O(N__64436),
            .I(\PROM.ROMDATA.m166_e ));
    InMux I__15146 (
            .O(N__64433),
            .I(N__64430));
    LocalMux I__15145 (
            .O(N__64430),
            .I(N__64427));
    Odrv4 I__15144 (
            .O(N__64427),
            .I(\PROM.ROMDATA.m104_ns_1 ));
    InMux I__15143 (
            .O(N__64424),
            .I(N__64421));
    LocalMux I__15142 (
            .O(N__64421),
            .I(\PROM.ROMDATA.m107 ));
    CascadeMux I__15141 (
            .O(N__64418),
            .I(\PROM.ROMDATA.m104_ns_cascade_ ));
    InMux I__15140 (
            .O(N__64415),
            .I(N__64412));
    LocalMux I__15139 (
            .O(N__64412),
            .I(N__64409));
    Span4Mux_v I__15138 (
            .O(N__64409),
            .I(N__64406));
    Span4Mux_h I__15137 (
            .O(N__64406),
            .I(N__64403));
    Odrv4 I__15136 (
            .O(N__64403),
            .I(\PROM.ROMDATA.m109_am ));
    CascadeMux I__15135 (
            .O(N__64400),
            .I(\PROM.ROMDATA.m109_bm_cascade_ ));
    InMux I__15134 (
            .O(N__64397),
            .I(N__64393));
    InMux I__15133 (
            .O(N__64396),
            .I(N__64390));
    LocalMux I__15132 (
            .O(N__64393),
            .I(N__64387));
    LocalMux I__15131 (
            .O(N__64390),
            .I(N__64382));
    Span4Mux_v I__15130 (
            .O(N__64387),
            .I(N__64382));
    Span4Mux_h I__15129 (
            .O(N__64382),
            .I(N__64379));
    Odrv4 I__15128 (
            .O(N__64379),
            .I(\PROM.ROMDATA.m121_ns ));
    InMux I__15127 (
            .O(N__64376),
            .I(N__64373));
    LocalMux I__15126 (
            .O(N__64373),
            .I(\PROM.ROMDATA.m114 ));
    InMux I__15125 (
            .O(N__64370),
            .I(N__64367));
    LocalMux I__15124 (
            .O(N__64367),
            .I(\PROM.ROMDATA.m111 ));
    CascadeMux I__15123 (
            .O(N__64364),
            .I(\PROM.ROMDATA.m120_am_cascade_ ));
    InMux I__15122 (
            .O(N__64361),
            .I(N__64358));
    LocalMux I__15121 (
            .O(N__64358),
            .I(\PROM.ROMDATA.m120_bm ));
    InMux I__15120 (
            .O(N__64355),
            .I(N__64352));
    LocalMux I__15119 (
            .O(N__64352),
            .I(\PROM.ROMDATA.m121_ns_1 ));
    CascadeMux I__15118 (
            .O(N__64349),
            .I(\PROM.ROMDATA.m287_cascade_ ));
    InMux I__15117 (
            .O(N__64346),
            .I(N__64343));
    LocalMux I__15116 (
            .O(N__64343),
            .I(\PROM.ROMDATA.m410_bm ));
    InMux I__15115 (
            .O(N__64340),
            .I(N__64337));
    LocalMux I__15114 (
            .O(N__64337),
            .I(N__64334));
    Span12Mux_v I__15113 (
            .O(N__64334),
            .I(N__64331));
    Odrv12 I__15112 (
            .O(N__64331),
            .I(\PROM.ROMDATA.m66 ));
    CascadeMux I__15111 (
            .O(N__64328),
            .I(N__64325));
    InMux I__15110 (
            .O(N__64325),
            .I(N__64320));
    CascadeMux I__15109 (
            .O(N__64324),
            .I(N__64317));
    InMux I__15108 (
            .O(N__64323),
            .I(N__64314));
    LocalMux I__15107 (
            .O(N__64320),
            .I(N__64311));
    InMux I__15106 (
            .O(N__64317),
            .I(N__64308));
    LocalMux I__15105 (
            .O(N__64314),
            .I(N__64305));
    Odrv4 I__15104 (
            .O(N__64311),
            .I(\PROM.ROMDATA.m163 ));
    LocalMux I__15103 (
            .O(N__64308),
            .I(\PROM.ROMDATA.m163 ));
    Odrv4 I__15102 (
            .O(N__64305),
            .I(\PROM.ROMDATA.m163 ));
    InMux I__15101 (
            .O(N__64298),
            .I(N__64295));
    LocalMux I__15100 (
            .O(N__64295),
            .I(N__64292));
    Span12Mux_v I__15099 (
            .O(N__64292),
            .I(N__64289));
    Odrv12 I__15098 (
            .O(N__64289),
            .I(\PROM.ROMDATA.m490 ));
    CascadeMux I__15097 (
            .O(N__64286),
            .I(N__64283));
    InMux I__15096 (
            .O(N__64283),
            .I(N__64280));
    LocalMux I__15095 (
            .O(N__64280),
            .I(\PROM.ROMDATA.m149 ));
    InMux I__15094 (
            .O(N__64277),
            .I(N__64274));
    LocalMux I__15093 (
            .O(N__64274),
            .I(\PROM.ROMDATA.m118 ));
    InMux I__15092 (
            .O(N__64271),
            .I(N__64268));
    LocalMux I__15091 (
            .O(N__64268),
            .I(\PROM.ROMDATA.m117 ));
    CascadeMux I__15090 (
            .O(N__64265),
            .I(N__64262));
    InMux I__15089 (
            .O(N__64262),
            .I(N__64258));
    InMux I__15088 (
            .O(N__64261),
            .I(N__64255));
    LocalMux I__15087 (
            .O(N__64258),
            .I(N__64251));
    LocalMux I__15086 (
            .O(N__64255),
            .I(N__64247));
    InMux I__15085 (
            .O(N__64254),
            .I(N__64242));
    Span4Mux_v I__15084 (
            .O(N__64251),
            .I(N__64239));
    InMux I__15083 (
            .O(N__64250),
            .I(N__64236));
    Span4Mux_v I__15082 (
            .O(N__64247),
            .I(N__64232));
    InMux I__15081 (
            .O(N__64246),
            .I(N__64229));
    InMux I__15080 (
            .O(N__64245),
            .I(N__64226));
    LocalMux I__15079 (
            .O(N__64242),
            .I(N__64223));
    Sp12to4 I__15078 (
            .O(N__64239),
            .I(N__64218));
    LocalMux I__15077 (
            .O(N__64236),
            .I(N__64218));
    InMux I__15076 (
            .O(N__64235),
            .I(N__64215));
    Odrv4 I__15075 (
            .O(N__64232),
            .I(\PROM.ROMDATA.m157 ));
    LocalMux I__15074 (
            .O(N__64229),
            .I(\PROM.ROMDATA.m157 ));
    LocalMux I__15073 (
            .O(N__64226),
            .I(\PROM.ROMDATA.m157 ));
    Odrv4 I__15072 (
            .O(N__64223),
            .I(\PROM.ROMDATA.m157 ));
    Odrv12 I__15071 (
            .O(N__64218),
            .I(\PROM.ROMDATA.m157 ));
    LocalMux I__15070 (
            .O(N__64215),
            .I(\PROM.ROMDATA.m157 ));
    CascadeMux I__15069 (
            .O(N__64202),
            .I(\PROM.ROMDATA.m456_ns_1_cascade_ ));
    InMux I__15068 (
            .O(N__64199),
            .I(N__64196));
    LocalMux I__15067 (
            .O(N__64196),
            .I(N__64193));
    Span4Mux_v I__15066 (
            .O(N__64193),
            .I(N__64190));
    Odrv4 I__15065 (
            .O(N__64190),
            .I(\PROM.ROMDATA.m456_ns ));
    InMux I__15064 (
            .O(N__64187),
            .I(N__64184));
    LocalMux I__15063 (
            .O(N__64184),
            .I(\PROM.ROMDATA.m414_ns_1 ));
    CascadeMux I__15062 (
            .O(N__64181),
            .I(N__64178));
    InMux I__15061 (
            .O(N__64178),
            .I(N__64175));
    LocalMux I__15060 (
            .O(N__64175),
            .I(N__64172));
    Odrv12 I__15059 (
            .O(N__64172),
            .I(\PROM.ROMDATA.m413_bm ));
    InMux I__15058 (
            .O(N__64169),
            .I(N__64166));
    LocalMux I__15057 (
            .O(N__64166),
            .I(N__64163));
    Span4Mux_h I__15056 (
            .O(N__64163),
            .I(N__64160));
    Odrv4 I__15055 (
            .O(N__64160),
            .I(\PROM.ROMDATA.m414_ns ));
    CascadeMux I__15054 (
            .O(N__64157),
            .I(N__64154));
    InMux I__15053 (
            .O(N__64154),
            .I(N__64151));
    LocalMux I__15052 (
            .O(N__64151),
            .I(N__64148));
    Odrv4 I__15051 (
            .O(N__64148),
            .I(\PROM.ROMDATA.m304 ));
    CascadeMux I__15050 (
            .O(N__64145),
            .I(PROM_ROMDATA_dintern_13ro_cascade_));
    CascadeMux I__15049 (
            .O(N__64142),
            .I(N__64139));
    InMux I__15048 (
            .O(N__64139),
            .I(N__64136));
    LocalMux I__15047 (
            .O(N__64136),
            .I(N__64133));
    Span4Mux_h I__15046 (
            .O(N__64133),
            .I(N__64130));
    Span4Mux_v I__15045 (
            .O(N__64130),
            .I(N__64127));
    Odrv4 I__15044 (
            .O(N__64127),
            .I(\PROM.ROMDATA.m198 ));
    InMux I__15043 (
            .O(N__64124),
            .I(N__64120));
    InMux I__15042 (
            .O(N__64123),
            .I(N__64117));
    LocalMux I__15041 (
            .O(N__64120),
            .I(N__64112));
    LocalMux I__15040 (
            .O(N__64117),
            .I(N__64112));
    Span4Mux_v I__15039 (
            .O(N__64112),
            .I(N__64109));
    Span4Mux_h I__15038 (
            .O(N__64109),
            .I(N__64102));
    InMux I__15037 (
            .O(N__64108),
            .I(N__64099));
    InMux I__15036 (
            .O(N__64107),
            .I(N__64092));
    InMux I__15035 (
            .O(N__64106),
            .I(N__64092));
    InMux I__15034 (
            .O(N__64105),
            .I(N__64092));
    Odrv4 I__15033 (
            .O(N__64102),
            .I(\PROM.ROMDATA.m16 ));
    LocalMux I__15032 (
            .O(N__64099),
            .I(\PROM.ROMDATA.m16 ));
    LocalMux I__15031 (
            .O(N__64092),
            .I(\PROM.ROMDATA.m16 ));
    InMux I__15030 (
            .O(N__64085),
            .I(N__64080));
    InMux I__15029 (
            .O(N__64084),
            .I(N__64075));
    InMux I__15028 (
            .O(N__64083),
            .I(N__64075));
    LocalMux I__15027 (
            .O(N__64080),
            .I(\CONTROL.N_45_0 ));
    LocalMux I__15026 (
            .O(N__64075),
            .I(\CONTROL.N_45_0 ));
    CascadeMux I__15025 (
            .O(N__64070),
            .I(PROM_ROMDATA_dintern_15ro_cascade_));
    CascadeMux I__15024 (
            .O(N__64067),
            .I(N__64064));
    InMux I__15023 (
            .O(N__64064),
            .I(N__64061));
    LocalMux I__15022 (
            .O(N__64061),
            .I(\PROM.ROMDATA.m139 ));
    CascadeMux I__15021 (
            .O(N__64058),
            .I(N__64054));
    InMux I__15020 (
            .O(N__64057),
            .I(N__64049));
    InMux I__15019 (
            .O(N__64054),
            .I(N__64049));
    LocalMux I__15018 (
            .O(N__64049),
            .I(N__64046));
    Span4Mux_v I__15017 (
            .O(N__64046),
            .I(N__64043));
    Span4Mux_h I__15016 (
            .O(N__64043),
            .I(N__64040));
    Span4Mux_h I__15015 (
            .O(N__64040),
            .I(N__64037));
    Span4Mux_v I__15014 (
            .O(N__64037),
            .I(N__64034));
    Odrv4 I__15013 (
            .O(N__64034),
            .I(\PROM.ROMDATA.N_564_mux ));
    InMux I__15012 (
            .O(N__64031),
            .I(N__64028));
    LocalMux I__15011 (
            .O(N__64028),
            .I(N__64025));
    Odrv4 I__15010 (
            .O(N__64025),
            .I(\PROM.ROMDATA.m298_bm ));
    InMux I__15009 (
            .O(N__64022),
            .I(N__64019));
    LocalMux I__15008 (
            .O(N__64019),
            .I(N__64014));
    CascadeMux I__15007 (
            .O(N__64018),
            .I(N__64011));
    InMux I__15006 (
            .O(N__64017),
            .I(N__64008));
    Span4Mux_h I__15005 (
            .O(N__64014),
            .I(N__64004));
    InMux I__15004 (
            .O(N__64011),
            .I(N__64001));
    LocalMux I__15003 (
            .O(N__64008),
            .I(N__63998));
    InMux I__15002 (
            .O(N__64007),
            .I(N__63995));
    Span4Mux_v I__15001 (
            .O(N__64004),
            .I(N__63992));
    LocalMux I__15000 (
            .O(N__64001),
            .I(N__63987));
    Span4Mux_v I__14999 (
            .O(N__63998),
            .I(N__63987));
    LocalMux I__14998 (
            .O(N__63995),
            .I(N__63984));
    Sp12to4 I__14997 (
            .O(N__63992),
            .I(N__63981));
    Span4Mux_v I__14996 (
            .O(N__63987),
            .I(N__63978));
    Span4Mux_h I__14995 (
            .O(N__63984),
            .I(N__63975));
    Odrv12 I__14994 (
            .O(N__63981),
            .I(\PROM.ROMDATA.N_72_i ));
    Odrv4 I__14993 (
            .O(N__63978),
            .I(\PROM.ROMDATA.N_72_i ));
    Odrv4 I__14992 (
            .O(N__63975),
            .I(\PROM.ROMDATA.N_72_i ));
    CascadeMux I__14991 (
            .O(N__63968),
            .I(N__63964));
    InMux I__14990 (
            .O(N__63967),
            .I(N__63959));
    InMux I__14989 (
            .O(N__63964),
            .I(N__63959));
    LocalMux I__14988 (
            .O(N__63959),
            .I(N__63956));
    Span12Mux_v I__14987 (
            .O(N__63956),
            .I(N__63953));
    Odrv12 I__14986 (
            .O(N__63953),
            .I(\PROM.ROMDATA.N_565_mux ));
    InMux I__14985 (
            .O(N__63950),
            .I(N__63947));
    LocalMux I__14984 (
            .O(N__63947),
            .I(N__63944));
    Span4Mux_h I__14983 (
            .O(N__63944),
            .I(N__63941));
    Odrv4 I__14982 (
            .O(N__63941),
            .I(\PROM.ROMDATA.m498_bm ));
    CascadeMux I__14981 (
            .O(N__63938),
            .I(\PROM.ROMDATA.m498_am_cascade_ ));
    CascadeMux I__14980 (
            .O(N__63935),
            .I(N__63932));
    InMux I__14979 (
            .O(N__63932),
            .I(N__63929));
    LocalMux I__14978 (
            .O(N__63929),
            .I(\PROM.ROMDATA.m498_ns ));
    InMux I__14977 (
            .O(N__63926),
            .I(N__63923));
    LocalMux I__14976 (
            .O(N__63923),
            .I(N__63920));
    Span12Mux_v I__14975 (
            .O(N__63920),
            .I(N__63917));
    Odrv12 I__14974 (
            .O(N__63917),
            .I(\PROM.ROMDATA.m317_am ));
    CascadeMux I__14973 (
            .O(N__63914),
            .I(\PROM.ROMDATA.m317_bm_cascade_ ));
    InMux I__14972 (
            .O(N__63911),
            .I(N__63908));
    LocalMux I__14971 (
            .O(N__63908),
            .I(N__63905));
    Span4Mux_v I__14970 (
            .O(N__63905),
            .I(N__63902));
    Odrv4 I__14969 (
            .O(N__63902),
            .I(\PROM.ROMDATA.m312_ns ));
    CascadeMux I__14968 (
            .O(N__63899),
            .I(\PROM.ROMDATA.m317_ns_cascade_ ));
    CascadeMux I__14967 (
            .O(N__63896),
            .I(\PROM.ROMDATA.m325_ns_1_cascade_ ));
    InMux I__14966 (
            .O(N__63893),
            .I(N__63890));
    LocalMux I__14965 (
            .O(N__63890),
            .I(N__63887));
    Odrv4 I__14964 (
            .O(N__63887),
            .I(\PROM.ROMDATA.m320_ns ));
    CascadeMux I__14963 (
            .O(N__63884),
            .I(N__63881));
    InMux I__14962 (
            .O(N__63881),
            .I(N__63878));
    LocalMux I__14961 (
            .O(N__63878),
            .I(N__63875));
    Odrv4 I__14960 (
            .O(N__63875),
            .I(\PROM.ROMDATA.m325_ns ));
    CascadeMux I__14959 (
            .O(N__63872),
            .I(PROM_ROMDATA_dintern_14ro_cascade_));
    InMux I__14958 (
            .O(N__63869),
            .I(N__63866));
    LocalMux I__14957 (
            .O(N__63866),
            .I(\PROM.ROMDATA.m494_ns ));
    InMux I__14956 (
            .O(N__63863),
            .I(\ALU.addsub_cry_12 ));
    InMux I__14955 (
            .O(N__63860),
            .I(N__63857));
    LocalMux I__14954 (
            .O(N__63857),
            .I(\ALU.c_RNIDDGOIZ0Z_14 ));
    CascadeMux I__14953 (
            .O(N__63854),
            .I(N__63849));
    CascadeMux I__14952 (
            .O(N__63853),
            .I(N__63844));
    InMux I__14951 (
            .O(N__63852),
            .I(N__63839));
    InMux I__14950 (
            .O(N__63849),
            .I(N__63836));
    CascadeMux I__14949 (
            .O(N__63848),
            .I(N__63832));
    InMux I__14948 (
            .O(N__63847),
            .I(N__63829));
    InMux I__14947 (
            .O(N__63844),
            .I(N__63826));
    InMux I__14946 (
            .O(N__63843),
            .I(N__63823));
    CascadeMux I__14945 (
            .O(N__63842),
            .I(N__63820));
    LocalMux I__14944 (
            .O(N__63839),
            .I(N__63816));
    LocalMux I__14943 (
            .O(N__63836),
            .I(N__63813));
    InMux I__14942 (
            .O(N__63835),
            .I(N__63810));
    InMux I__14941 (
            .O(N__63832),
            .I(N__63806));
    LocalMux I__14940 (
            .O(N__63829),
            .I(N__63803));
    LocalMux I__14939 (
            .O(N__63826),
            .I(N__63797));
    LocalMux I__14938 (
            .O(N__63823),
            .I(N__63797));
    InMux I__14937 (
            .O(N__63820),
            .I(N__63794));
    CascadeMux I__14936 (
            .O(N__63819),
            .I(N__63791));
    Span4Mux_v I__14935 (
            .O(N__63816),
            .I(N__63788));
    Span4Mux_v I__14934 (
            .O(N__63813),
            .I(N__63783));
    LocalMux I__14933 (
            .O(N__63810),
            .I(N__63783));
    InMux I__14932 (
            .O(N__63809),
            .I(N__63780));
    LocalMux I__14931 (
            .O(N__63806),
            .I(N__63775));
    Span4Mux_v I__14930 (
            .O(N__63803),
            .I(N__63771));
    InMux I__14929 (
            .O(N__63802),
            .I(N__63768));
    Span4Mux_v I__14928 (
            .O(N__63797),
            .I(N__63763));
    LocalMux I__14927 (
            .O(N__63794),
            .I(N__63763));
    InMux I__14926 (
            .O(N__63791),
            .I(N__63760));
    Span4Mux_h I__14925 (
            .O(N__63788),
            .I(N__63753));
    Span4Mux_h I__14924 (
            .O(N__63783),
            .I(N__63753));
    LocalMux I__14923 (
            .O(N__63780),
            .I(N__63753));
    InMux I__14922 (
            .O(N__63779),
            .I(N__63748));
    InMux I__14921 (
            .O(N__63778),
            .I(N__63748));
    Span4Mux_v I__14920 (
            .O(N__63775),
            .I(N__63745));
    InMux I__14919 (
            .O(N__63774),
            .I(N__63742));
    Span4Mux_v I__14918 (
            .O(N__63771),
            .I(N__63739));
    LocalMux I__14917 (
            .O(N__63768),
            .I(N__63734));
    Span4Mux_v I__14916 (
            .O(N__63763),
            .I(N__63734));
    LocalMux I__14915 (
            .O(N__63760),
            .I(N__63731));
    Span4Mux_v I__14914 (
            .O(N__63753),
            .I(N__63728));
    LocalMux I__14913 (
            .O(N__63748),
            .I(N__63721));
    Span4Mux_v I__14912 (
            .O(N__63745),
            .I(N__63721));
    LocalMux I__14911 (
            .O(N__63742),
            .I(N__63721));
    Span4Mux_h I__14910 (
            .O(N__63739),
            .I(N__63716));
    Span4Mux_v I__14909 (
            .O(N__63734),
            .I(N__63716));
    Span4Mux_v I__14908 (
            .O(N__63731),
            .I(N__63711));
    Span4Mux_v I__14907 (
            .O(N__63728),
            .I(N__63711));
    Span4Mux_v I__14906 (
            .O(N__63721),
            .I(N__63706));
    Span4Mux_h I__14905 (
            .O(N__63716),
            .I(N__63706));
    Odrv4 I__14904 (
            .O(N__63711),
            .I(aluOut_14));
    Odrv4 I__14903 (
            .O(N__63706),
            .I(aluOut_14));
    InMux I__14902 (
            .O(N__63701),
            .I(N__63694));
    InMux I__14901 (
            .O(N__63700),
            .I(N__63694));
    InMux I__14900 (
            .O(N__63699),
            .I(N__63691));
    LocalMux I__14899 (
            .O(N__63694),
            .I(N__63688));
    LocalMux I__14898 (
            .O(N__63691),
            .I(\ALU.addsub_14 ));
    Odrv12 I__14897 (
            .O(N__63688),
            .I(\ALU.addsub_14 ));
    InMux I__14896 (
            .O(N__63683),
            .I(\ALU.addsub_cry_13 ));
    InMux I__14895 (
            .O(N__63680),
            .I(N__63677));
    LocalMux I__14894 (
            .O(N__63677),
            .I(\ALU.c_RNI0NMSHZ0Z_15 ));
    InMux I__14893 (
            .O(N__63674),
            .I(N__63671));
    LocalMux I__14892 (
            .O(N__63671),
            .I(N__63665));
    CascadeMux I__14891 (
            .O(N__63670),
            .I(N__63662));
    InMux I__14890 (
            .O(N__63669),
            .I(N__63659));
    InMux I__14889 (
            .O(N__63668),
            .I(N__63655));
    Span4Mux_h I__14888 (
            .O(N__63665),
            .I(N__63652));
    InMux I__14887 (
            .O(N__63662),
            .I(N__63649));
    LocalMux I__14886 (
            .O(N__63659),
            .I(N__63646));
    InMux I__14885 (
            .O(N__63658),
            .I(N__63641));
    LocalMux I__14884 (
            .O(N__63655),
            .I(N__63635));
    Span4Mux_h I__14883 (
            .O(N__63652),
            .I(N__63628));
    LocalMux I__14882 (
            .O(N__63649),
            .I(N__63628));
    Span4Mux_v I__14881 (
            .O(N__63646),
            .I(N__63628));
    InMux I__14880 (
            .O(N__63645),
            .I(N__63625));
    InMux I__14879 (
            .O(N__63644),
            .I(N__63622));
    LocalMux I__14878 (
            .O(N__63641),
            .I(N__63619));
    InMux I__14877 (
            .O(N__63640),
            .I(N__63616));
    InMux I__14876 (
            .O(N__63639),
            .I(N__63607));
    InMux I__14875 (
            .O(N__63638),
            .I(N__63607));
    Span4Mux_v I__14874 (
            .O(N__63635),
            .I(N__63598));
    Span4Mux_h I__14873 (
            .O(N__63628),
            .I(N__63598));
    LocalMux I__14872 (
            .O(N__63625),
            .I(N__63598));
    LocalMux I__14871 (
            .O(N__63622),
            .I(N__63598));
    Span4Mux_h I__14870 (
            .O(N__63619),
            .I(N__63595));
    LocalMux I__14869 (
            .O(N__63616),
            .I(N__63589));
    InMux I__14868 (
            .O(N__63615),
            .I(N__63586));
    CascadeMux I__14867 (
            .O(N__63614),
            .I(N__63583));
    CascadeMux I__14866 (
            .O(N__63613),
            .I(N__63579));
    CascadeMux I__14865 (
            .O(N__63612),
            .I(N__63576));
    LocalMux I__14864 (
            .O(N__63607),
            .I(N__63571));
    Span4Mux_h I__14863 (
            .O(N__63598),
            .I(N__63571));
    Span4Mux_h I__14862 (
            .O(N__63595),
            .I(N__63568));
    InMux I__14861 (
            .O(N__63594),
            .I(N__63561));
    InMux I__14860 (
            .O(N__63593),
            .I(N__63561));
    InMux I__14859 (
            .O(N__63592),
            .I(N__63561));
    Span12Mux_s10_h I__14858 (
            .O(N__63589),
            .I(N__63558));
    LocalMux I__14857 (
            .O(N__63586),
            .I(N__63555));
    InMux I__14856 (
            .O(N__63583),
            .I(N__63548));
    InMux I__14855 (
            .O(N__63582),
            .I(N__63548));
    InMux I__14854 (
            .O(N__63579),
            .I(N__63548));
    InMux I__14853 (
            .O(N__63576),
            .I(N__63545));
    Span4Mux_v I__14852 (
            .O(N__63571),
            .I(N__63542));
    Span4Mux_v I__14851 (
            .O(N__63568),
            .I(N__63537));
    LocalMux I__14850 (
            .O(N__63561),
            .I(N__63537));
    Odrv12 I__14849 (
            .O(N__63558),
            .I(aluOut_15));
    Odrv12 I__14848 (
            .O(N__63555),
            .I(aluOut_15));
    LocalMux I__14847 (
            .O(N__63548),
            .I(aluOut_15));
    LocalMux I__14846 (
            .O(N__63545),
            .I(aluOut_15));
    Odrv4 I__14845 (
            .O(N__63542),
            .I(aluOut_15));
    Odrv4 I__14844 (
            .O(N__63537),
            .I(aluOut_15));
    InMux I__14843 (
            .O(N__63524),
            .I(N__63520));
    InMux I__14842 (
            .O(N__63523),
            .I(N__63517));
    LocalMux I__14841 (
            .O(N__63520),
            .I(N__63513));
    LocalMux I__14840 (
            .O(N__63517),
            .I(N__63509));
    InMux I__14839 (
            .O(N__63516),
            .I(N__63506));
    Span4Mux_h I__14838 (
            .O(N__63513),
            .I(N__63503));
    InMux I__14837 (
            .O(N__63512),
            .I(N__63500));
    Span4Mux_h I__14836 (
            .O(N__63509),
            .I(N__63497));
    LocalMux I__14835 (
            .O(N__63506),
            .I(\ALU.addsub_15 ));
    Odrv4 I__14834 (
            .O(N__63503),
            .I(\ALU.addsub_15 ));
    LocalMux I__14833 (
            .O(N__63500),
            .I(\ALU.addsub_15 ));
    Odrv4 I__14832 (
            .O(N__63497),
            .I(\ALU.addsub_15 ));
    InMux I__14831 (
            .O(N__63488),
            .I(bfn_23_16_0_));
    CascadeMux I__14830 (
            .O(N__63485),
            .I(N__63482));
    InMux I__14829 (
            .O(N__63482),
            .I(N__63478));
    CascadeMux I__14828 (
            .O(N__63481),
            .I(N__63475));
    LocalMux I__14827 (
            .O(N__63478),
            .I(N__63472));
    InMux I__14826 (
            .O(N__63475),
            .I(N__63469));
    Span4Mux_h I__14825 (
            .O(N__63472),
            .I(N__63464));
    LocalMux I__14824 (
            .O(N__63469),
            .I(N__63464));
    Span4Mux_h I__14823 (
            .O(N__63464),
            .I(N__63456));
    InMux I__14822 (
            .O(N__63463),
            .I(N__63453));
    InMux I__14821 (
            .O(N__63462),
            .I(N__63448));
    InMux I__14820 (
            .O(N__63461),
            .I(N__63448));
    InMux I__14819 (
            .O(N__63460),
            .I(N__63443));
    InMux I__14818 (
            .O(N__63459),
            .I(N__63443));
    Span4Mux_v I__14817 (
            .O(N__63456),
            .I(N__63435));
    LocalMux I__14816 (
            .O(N__63453),
            .I(N__63435));
    LocalMux I__14815 (
            .O(N__63448),
            .I(N__63435));
    LocalMux I__14814 (
            .O(N__63443),
            .I(N__63432));
    InMux I__14813 (
            .O(N__63442),
            .I(N__63429));
    Span4Mux_h I__14812 (
            .O(N__63435),
            .I(N__63426));
    Span4Mux_v I__14811 (
            .O(N__63432),
            .I(N__63423));
    LocalMux I__14810 (
            .O(N__63429),
            .I(N__63418));
    Span4Mux_h I__14809 (
            .O(N__63426),
            .I(N__63418));
    Span4Mux_h I__14808 (
            .O(N__63423),
            .I(N__63415));
    Span4Mux_v I__14807 (
            .O(N__63418),
            .I(N__63411));
    Span4Mux_v I__14806 (
            .O(N__63415),
            .I(N__63408));
    InMux I__14805 (
            .O(N__63414),
            .I(N__63405));
    Span4Mux_v I__14804 (
            .O(N__63411),
            .I(N__63402));
    Span4Mux_v I__14803 (
            .O(N__63408),
            .I(N__63399));
    LocalMux I__14802 (
            .O(N__63405),
            .I(aluStatus_1));
    Odrv4 I__14801 (
            .O(N__63402),
            .I(aluStatus_1));
    Odrv4 I__14800 (
            .O(N__63399),
            .I(aluStatus_1));
    InMux I__14799 (
            .O(N__63392),
            .I(\ALU.addsub_cry_15 ));
    InMux I__14798 (
            .O(N__63389),
            .I(N__63386));
    LocalMux I__14797 (
            .O(N__63386),
            .I(N__63383));
    Odrv12 I__14796 (
            .O(N__63383),
            .I(\ALU.N_545 ));
    IoInMux I__14795 (
            .O(N__63380),
            .I(N__63377));
    LocalMux I__14794 (
            .O(N__63377),
            .I(N__63374));
    Span4Mux_s1_h I__14793 (
            .O(N__63374),
            .I(N__63371));
    Span4Mux_v I__14792 (
            .O(N__63371),
            .I(N__63367));
    IoInMux I__14791 (
            .O(N__63370),
            .I(N__63364));
    Span4Mux_v I__14790 (
            .O(N__63367),
            .I(N__63361));
    LocalMux I__14789 (
            .O(N__63364),
            .I(N__63357));
    Span4Mux_h I__14788 (
            .O(N__63361),
            .I(N__63354));
    InMux I__14787 (
            .O(N__63360),
            .I(N__63351));
    IoSpan4Mux I__14786 (
            .O(N__63357),
            .I(N__63348));
    Span4Mux_h I__14785 (
            .O(N__63354),
            .I(N__63343));
    LocalMux I__14784 (
            .O(N__63351),
            .I(N__63343));
    Span4Mux_s3_h I__14783 (
            .O(N__63348),
            .I(N__63340));
    Span4Mux_v I__14782 (
            .O(N__63343),
            .I(N__63337));
    Sp12to4 I__14781 (
            .O(N__63340),
            .I(N__63334));
    Sp12to4 I__14780 (
            .O(N__63337),
            .I(N__63331));
    Span12Mux_v I__14779 (
            .O(N__63334),
            .I(N__63328));
    Span12Mux_h I__14778 (
            .O(N__63331),
            .I(N__63325));
    Odrv12 I__14777 (
            .O(N__63328),
            .I(bus_6));
    Odrv12 I__14776 (
            .O(N__63325),
            .I(bus_6));
    InMux I__14775 (
            .O(N__63320),
            .I(N__63314));
    InMux I__14774 (
            .O(N__63319),
            .I(N__63314));
    LocalMux I__14773 (
            .O(N__63314),
            .I(N__63311));
    Span4Mux_h I__14772 (
            .O(N__63311),
            .I(N__63308));
    Span4Mux_h I__14771 (
            .O(N__63308),
            .I(N__63305));
    Odrv4 I__14770 (
            .O(N__63305),
            .I(\ALU.c_RNIPBAG72Z0Z_14 ));
    CascadeMux I__14769 (
            .O(N__63302),
            .I(N__63294));
    InMux I__14768 (
            .O(N__63301),
            .I(N__63280));
    InMux I__14767 (
            .O(N__63300),
            .I(N__63280));
    InMux I__14766 (
            .O(N__63299),
            .I(N__63280));
    InMux I__14765 (
            .O(N__63298),
            .I(N__63280));
    CascadeMux I__14764 (
            .O(N__63297),
            .I(N__63277));
    InMux I__14763 (
            .O(N__63294),
            .I(N__63270));
    CascadeMux I__14762 (
            .O(N__63293),
            .I(N__63266));
    CascadeMux I__14761 (
            .O(N__63292),
            .I(N__63262));
    InMux I__14760 (
            .O(N__63291),
            .I(N__63257));
    CascadeMux I__14759 (
            .O(N__63290),
            .I(N__63250));
    InMux I__14758 (
            .O(N__63289),
            .I(N__63243));
    LocalMux I__14757 (
            .O(N__63280),
            .I(N__63235));
    InMux I__14756 (
            .O(N__63277),
            .I(N__63232));
    InMux I__14755 (
            .O(N__63276),
            .I(N__63229));
    CascadeMux I__14754 (
            .O(N__63275),
            .I(N__63226));
    CascadeMux I__14753 (
            .O(N__63274),
            .I(N__63222));
    CascadeMux I__14752 (
            .O(N__63273),
            .I(N__63219));
    LocalMux I__14751 (
            .O(N__63270),
            .I(N__63214));
    InMux I__14750 (
            .O(N__63269),
            .I(N__63209));
    InMux I__14749 (
            .O(N__63266),
            .I(N__63209));
    InMux I__14748 (
            .O(N__63265),
            .I(N__63204));
    InMux I__14747 (
            .O(N__63262),
            .I(N__63204));
    InMux I__14746 (
            .O(N__63261),
            .I(N__63199));
    InMux I__14745 (
            .O(N__63260),
            .I(N__63199));
    LocalMux I__14744 (
            .O(N__63257),
            .I(N__63196));
    InMux I__14743 (
            .O(N__63256),
            .I(N__63193));
    InMux I__14742 (
            .O(N__63255),
            .I(N__63188));
    InMux I__14741 (
            .O(N__63254),
            .I(N__63188));
    InMux I__14740 (
            .O(N__63253),
            .I(N__63185));
    InMux I__14739 (
            .O(N__63250),
            .I(N__63178));
    InMux I__14738 (
            .O(N__63249),
            .I(N__63178));
    InMux I__14737 (
            .O(N__63248),
            .I(N__63178));
    InMux I__14736 (
            .O(N__63247),
            .I(N__63173));
    InMux I__14735 (
            .O(N__63246),
            .I(N__63173));
    LocalMux I__14734 (
            .O(N__63243),
            .I(N__63170));
    InMux I__14733 (
            .O(N__63242),
            .I(N__63163));
    InMux I__14732 (
            .O(N__63241),
            .I(N__63163));
    InMux I__14731 (
            .O(N__63240),
            .I(N__63163));
    InMux I__14730 (
            .O(N__63239),
            .I(N__63158));
    InMux I__14729 (
            .O(N__63238),
            .I(N__63158));
    Span4Mux_v I__14728 (
            .O(N__63235),
            .I(N__63151));
    LocalMux I__14727 (
            .O(N__63232),
            .I(N__63151));
    LocalMux I__14726 (
            .O(N__63229),
            .I(N__63151));
    InMux I__14725 (
            .O(N__63226),
            .I(N__63147));
    InMux I__14724 (
            .O(N__63225),
            .I(N__63142));
    InMux I__14723 (
            .O(N__63222),
            .I(N__63142));
    InMux I__14722 (
            .O(N__63219),
            .I(N__63135));
    InMux I__14721 (
            .O(N__63218),
            .I(N__63135));
    InMux I__14720 (
            .O(N__63217),
            .I(N__63135));
    Span4Mux_v I__14719 (
            .O(N__63214),
            .I(N__63132));
    LocalMux I__14718 (
            .O(N__63209),
            .I(N__63125));
    LocalMux I__14717 (
            .O(N__63204),
            .I(N__63125));
    LocalMux I__14716 (
            .O(N__63199),
            .I(N__63125));
    Span4Mux_v I__14715 (
            .O(N__63196),
            .I(N__63122));
    LocalMux I__14714 (
            .O(N__63193),
            .I(N__63117));
    LocalMux I__14713 (
            .O(N__63188),
            .I(N__63117));
    LocalMux I__14712 (
            .O(N__63185),
            .I(N__63109));
    LocalMux I__14711 (
            .O(N__63178),
            .I(N__63106));
    LocalMux I__14710 (
            .O(N__63173),
            .I(N__63103));
    Span4Mux_v I__14709 (
            .O(N__63170),
            .I(N__63100));
    LocalMux I__14708 (
            .O(N__63163),
            .I(N__63093));
    LocalMux I__14707 (
            .O(N__63158),
            .I(N__63093));
    Span4Mux_v I__14706 (
            .O(N__63151),
            .I(N__63093));
    InMux I__14705 (
            .O(N__63150),
            .I(N__63090));
    LocalMux I__14704 (
            .O(N__63147),
            .I(N__63087));
    LocalMux I__14703 (
            .O(N__63142),
            .I(N__63082));
    LocalMux I__14702 (
            .O(N__63135),
            .I(N__63082));
    Span4Mux_v I__14701 (
            .O(N__63132),
            .I(N__63077));
    Span4Mux_v I__14700 (
            .O(N__63125),
            .I(N__63077));
    Span4Mux_v I__14699 (
            .O(N__63122),
            .I(N__63070));
    Span4Mux_v I__14698 (
            .O(N__63117),
            .I(N__63070));
    InMux I__14697 (
            .O(N__63116),
            .I(N__63067));
    InMux I__14696 (
            .O(N__63115),
            .I(N__63062));
    InMux I__14695 (
            .O(N__63114),
            .I(N__63062));
    InMux I__14694 (
            .O(N__63113),
            .I(N__63059));
    InMux I__14693 (
            .O(N__63112),
            .I(N__63056));
    Span4Mux_v I__14692 (
            .O(N__63109),
            .I(N__63053));
    Span4Mux_v I__14691 (
            .O(N__63106),
            .I(N__63050));
    Span4Mux_v I__14690 (
            .O(N__63103),
            .I(N__63047));
    Span4Mux_h I__14689 (
            .O(N__63100),
            .I(N__63044));
    Span4Mux_v I__14688 (
            .O(N__63093),
            .I(N__63041));
    LocalMux I__14687 (
            .O(N__63090),
            .I(N__63036));
    Span4Mux_v I__14686 (
            .O(N__63087),
            .I(N__63036));
    Span4Mux_h I__14685 (
            .O(N__63082),
            .I(N__63031));
    Span4Mux_h I__14684 (
            .O(N__63077),
            .I(N__63031));
    CascadeMux I__14683 (
            .O(N__63076),
            .I(N__63027));
    CascadeMux I__14682 (
            .O(N__63075),
            .I(N__63023));
    Sp12to4 I__14681 (
            .O(N__63070),
            .I(N__63009));
    LocalMux I__14680 (
            .O(N__63067),
            .I(N__63009));
    LocalMux I__14679 (
            .O(N__63062),
            .I(N__63009));
    LocalMux I__14678 (
            .O(N__63059),
            .I(N__63009));
    LocalMux I__14677 (
            .O(N__63056),
            .I(N__63009));
    Sp12to4 I__14676 (
            .O(N__63053),
            .I(N__63009));
    Sp12to4 I__14675 (
            .O(N__63050),
            .I(N__63004));
    Sp12to4 I__14674 (
            .O(N__63047),
            .I(N__63004));
    Sp12to4 I__14673 (
            .O(N__63044),
            .I(N__63001));
    Span4Mux_h I__14672 (
            .O(N__63041),
            .I(N__62998));
    Span4Mux_v I__14671 (
            .O(N__63036),
            .I(N__62993));
    Span4Mux_h I__14670 (
            .O(N__63031),
            .I(N__62993));
    InMux I__14669 (
            .O(N__63030),
            .I(N__62986));
    InMux I__14668 (
            .O(N__63027),
            .I(N__62986));
    InMux I__14667 (
            .O(N__63026),
            .I(N__62986));
    InMux I__14666 (
            .O(N__63023),
            .I(N__62981));
    InMux I__14665 (
            .O(N__63022),
            .I(N__62981));
    Span12Mux_h I__14664 (
            .O(N__63009),
            .I(N__62978));
    Span12Mux_h I__14663 (
            .O(N__63004),
            .I(N__62973));
    Span12Mux_v I__14662 (
            .O(N__63001),
            .I(N__62973));
    Span4Mux_h I__14661 (
            .O(N__62998),
            .I(N__62968));
    Span4Mux_v I__14660 (
            .O(N__62993),
            .I(N__62968));
    LocalMux I__14659 (
            .O(N__62986),
            .I(aluParams_0));
    LocalMux I__14658 (
            .O(N__62981),
            .I(aluParams_0));
    Odrv12 I__14657 (
            .O(N__62978),
            .I(aluParams_0));
    Odrv12 I__14656 (
            .O(N__62973),
            .I(aluParams_0));
    Odrv4 I__14655 (
            .O(N__62968),
            .I(aluParams_0));
    CascadeMux I__14654 (
            .O(N__62957),
            .I(N__62953));
    CascadeMux I__14653 (
            .O(N__62956),
            .I(N__62950));
    InMux I__14652 (
            .O(N__62953),
            .I(N__62946));
    InMux I__14651 (
            .O(N__62950),
            .I(N__62943));
    CascadeMux I__14650 (
            .O(N__62949),
            .I(N__62940));
    LocalMux I__14649 (
            .O(N__62946),
            .I(N__62936));
    LocalMux I__14648 (
            .O(N__62943),
            .I(N__62933));
    InMux I__14647 (
            .O(N__62940),
            .I(N__62928));
    InMux I__14646 (
            .O(N__62939),
            .I(N__62928));
    Span4Mux_h I__14645 (
            .O(N__62936),
            .I(N__62922));
    Span4Mux_v I__14644 (
            .O(N__62933),
            .I(N__62922));
    LocalMux I__14643 (
            .O(N__62928),
            .I(N__62919));
    InMux I__14642 (
            .O(N__62927),
            .I(N__62916));
    Span4Mux_h I__14641 (
            .O(N__62922),
            .I(N__62913));
    Span4Mux_v I__14640 (
            .O(N__62919),
            .I(N__62910));
    LocalMux I__14639 (
            .O(N__62916),
            .I(N__62907));
    Span4Mux_h I__14638 (
            .O(N__62913),
            .I(N__62904));
    Span4Mux_v I__14637 (
            .O(N__62910),
            .I(N__62899));
    Span4Mux_h I__14636 (
            .O(N__62907),
            .I(N__62899));
    Span4Mux_v I__14635 (
            .O(N__62904),
            .I(N__62894));
    Span4Mux_h I__14634 (
            .O(N__62899),
            .I(N__62894));
    Odrv4 I__14633 (
            .O(N__62894),
            .I(\ALU.combOperand2_0_9 ));
    InMux I__14632 (
            .O(N__62891),
            .I(N__62878));
    InMux I__14631 (
            .O(N__62890),
            .I(N__62875));
    InMux I__14630 (
            .O(N__62889),
            .I(N__62868));
    InMux I__14629 (
            .O(N__62888),
            .I(N__62863));
    InMux I__14628 (
            .O(N__62887),
            .I(N__62863));
    CascadeMux I__14627 (
            .O(N__62886),
            .I(N__62860));
    InMux I__14626 (
            .O(N__62885),
            .I(N__62856));
    InMux I__14625 (
            .O(N__62884),
            .I(N__62849));
    InMux I__14624 (
            .O(N__62883),
            .I(N__62849));
    InMux I__14623 (
            .O(N__62882),
            .I(N__62849));
    InMux I__14622 (
            .O(N__62881),
            .I(N__62846));
    LocalMux I__14621 (
            .O(N__62878),
            .I(N__62842));
    LocalMux I__14620 (
            .O(N__62875),
            .I(N__62839));
    InMux I__14619 (
            .O(N__62874),
            .I(N__62836));
    InMux I__14618 (
            .O(N__62873),
            .I(N__62833));
    InMux I__14617 (
            .O(N__62872),
            .I(N__62830));
    InMux I__14616 (
            .O(N__62871),
            .I(N__62826));
    LocalMux I__14615 (
            .O(N__62868),
            .I(N__62821));
    LocalMux I__14614 (
            .O(N__62863),
            .I(N__62821));
    InMux I__14613 (
            .O(N__62860),
            .I(N__62815));
    InMux I__14612 (
            .O(N__62859),
            .I(N__62812));
    LocalMux I__14611 (
            .O(N__62856),
            .I(N__62806));
    LocalMux I__14610 (
            .O(N__62849),
            .I(N__62806));
    LocalMux I__14609 (
            .O(N__62846),
            .I(N__62802));
    InMux I__14608 (
            .O(N__62845),
            .I(N__62798));
    Span4Mux_v I__14607 (
            .O(N__62842),
            .I(N__62793));
    Span4Mux_v I__14606 (
            .O(N__62839),
            .I(N__62793));
    LocalMux I__14605 (
            .O(N__62836),
            .I(N__62786));
    LocalMux I__14604 (
            .O(N__62833),
            .I(N__62786));
    LocalMux I__14603 (
            .O(N__62830),
            .I(N__62786));
    InMux I__14602 (
            .O(N__62829),
            .I(N__62782));
    LocalMux I__14601 (
            .O(N__62826),
            .I(N__62777));
    Span4Mux_v I__14600 (
            .O(N__62821),
            .I(N__62777));
    InMux I__14599 (
            .O(N__62820),
            .I(N__62774));
    InMux I__14598 (
            .O(N__62819),
            .I(N__62769));
    InMux I__14597 (
            .O(N__62818),
            .I(N__62769));
    LocalMux I__14596 (
            .O(N__62815),
            .I(N__62766));
    LocalMux I__14595 (
            .O(N__62812),
            .I(N__62761));
    InMux I__14594 (
            .O(N__62811),
            .I(N__62758));
    Span4Mux_h I__14593 (
            .O(N__62806),
            .I(N__62755));
    InMux I__14592 (
            .O(N__62805),
            .I(N__62752));
    Span4Mux_v I__14591 (
            .O(N__62802),
            .I(N__62749));
    InMux I__14590 (
            .O(N__62801),
            .I(N__62746));
    LocalMux I__14589 (
            .O(N__62798),
            .I(N__62739));
    Span4Mux_h I__14588 (
            .O(N__62793),
            .I(N__62739));
    Span4Mux_v I__14587 (
            .O(N__62786),
            .I(N__62739));
    InMux I__14586 (
            .O(N__62785),
            .I(N__62736));
    LocalMux I__14585 (
            .O(N__62782),
            .I(N__62733));
    Span4Mux_h I__14584 (
            .O(N__62777),
            .I(N__62726));
    LocalMux I__14583 (
            .O(N__62774),
            .I(N__62726));
    LocalMux I__14582 (
            .O(N__62769),
            .I(N__62726));
    Span4Mux_v I__14581 (
            .O(N__62766),
            .I(N__62723));
    InMux I__14580 (
            .O(N__62765),
            .I(N__62718));
    InMux I__14579 (
            .O(N__62764),
            .I(N__62718));
    Span4Mux_v I__14578 (
            .O(N__62761),
            .I(N__62709));
    LocalMux I__14577 (
            .O(N__62758),
            .I(N__62709));
    Span4Mux_v I__14576 (
            .O(N__62755),
            .I(N__62709));
    LocalMux I__14575 (
            .O(N__62752),
            .I(N__62709));
    Sp12to4 I__14574 (
            .O(N__62749),
            .I(N__62704));
    LocalMux I__14573 (
            .O(N__62746),
            .I(N__62704));
    Span4Mux_v I__14572 (
            .O(N__62739),
            .I(N__62701));
    LocalMux I__14571 (
            .O(N__62736),
            .I(N__62698));
    Span4Mux_h I__14570 (
            .O(N__62733),
            .I(N__62693));
    Span4Mux_h I__14569 (
            .O(N__62726),
            .I(N__62693));
    Span4Mux_v I__14568 (
            .O(N__62723),
            .I(N__62688));
    LocalMux I__14567 (
            .O(N__62718),
            .I(N__62688));
    Span4Mux_h I__14566 (
            .O(N__62709),
            .I(N__62685));
    Odrv12 I__14565 (
            .O(N__62704),
            .I(aluOut_9));
    Odrv4 I__14564 (
            .O(N__62701),
            .I(aluOut_9));
    Odrv12 I__14563 (
            .O(N__62698),
            .I(aluOut_9));
    Odrv4 I__14562 (
            .O(N__62693),
            .I(aluOut_9));
    Odrv4 I__14561 (
            .O(N__62688),
            .I(aluOut_9));
    Odrv4 I__14560 (
            .O(N__62685),
            .I(aluOut_9));
    CascadeMux I__14559 (
            .O(N__62672),
            .I(N__62669));
    InMux I__14558 (
            .O(N__62669),
            .I(N__62666));
    LocalMux I__14557 (
            .O(N__62666),
            .I(\ALU.d_RNI70I1IZ0Z_9 ));
    InMux I__14556 (
            .O(N__62663),
            .I(N__62660));
    LocalMux I__14555 (
            .O(N__62660),
            .I(N__62657));
    Span4Mux_h I__14554 (
            .O(N__62657),
            .I(N__62652));
    CascadeMux I__14553 (
            .O(N__62656),
            .I(N__62649));
    InMux I__14552 (
            .O(N__62655),
            .I(N__62645));
    Span4Mux_v I__14551 (
            .O(N__62652),
            .I(N__62642));
    InMux I__14550 (
            .O(N__62649),
            .I(N__62639));
    InMux I__14549 (
            .O(N__62648),
            .I(N__62636));
    LocalMux I__14548 (
            .O(N__62645),
            .I(\ALU.N_980 ));
    Odrv4 I__14547 (
            .O(N__62642),
            .I(\ALU.N_980 ));
    LocalMux I__14546 (
            .O(N__62639),
            .I(\ALU.N_980 ));
    LocalMux I__14545 (
            .O(N__62636),
            .I(\ALU.N_980 ));
    InMux I__14544 (
            .O(N__62627),
            .I(N__62624));
    LocalMux I__14543 (
            .O(N__62624),
            .I(\ALU.N_1029 ));
    InMux I__14542 (
            .O(N__62621),
            .I(N__62618));
    LocalMux I__14541 (
            .O(N__62618),
            .I(N__62615));
    Span4Mux_h I__14540 (
            .O(N__62615),
            .I(N__62612));
    Odrv4 I__14539 (
            .O(N__62612),
            .I(\PROM.ROMDATA.m500_ns_1 ));
    InMux I__14538 (
            .O(N__62609),
            .I(N__62603));
    InMux I__14537 (
            .O(N__62608),
            .I(N__62603));
    LocalMux I__14536 (
            .O(N__62603),
            .I(N__62600));
    Span4Mux_h I__14535 (
            .O(N__62600),
            .I(N__62597));
    Span4Mux_h I__14534 (
            .O(N__62597),
            .I(N__62594));
    Span4Mux_v I__14533 (
            .O(N__62594),
            .I(N__62591));
    Odrv4 I__14532 (
            .O(N__62591),
            .I(\PROM.ROMDATA.m500_ns ));
    CascadeMux I__14531 (
            .O(N__62588),
            .I(N__62580));
    InMux I__14530 (
            .O(N__62587),
            .I(N__62576));
    InMux I__14529 (
            .O(N__62586),
            .I(N__62573));
    CascadeMux I__14528 (
            .O(N__62585),
            .I(N__62567));
    CascadeMux I__14527 (
            .O(N__62584),
            .I(N__62564));
    InMux I__14526 (
            .O(N__62583),
            .I(N__62559));
    InMux I__14525 (
            .O(N__62580),
            .I(N__62559));
    CascadeMux I__14524 (
            .O(N__62579),
            .I(N__62553));
    LocalMux I__14523 (
            .O(N__62576),
            .I(N__62547));
    LocalMux I__14522 (
            .O(N__62573),
            .I(N__62544));
    CascadeMux I__14521 (
            .O(N__62572),
            .I(N__62541));
    InMux I__14520 (
            .O(N__62571),
            .I(N__62538));
    InMux I__14519 (
            .O(N__62570),
            .I(N__62535));
    InMux I__14518 (
            .O(N__62567),
            .I(N__62530));
    InMux I__14517 (
            .O(N__62564),
            .I(N__62530));
    LocalMux I__14516 (
            .O(N__62559),
            .I(N__62527));
    InMux I__14515 (
            .O(N__62558),
            .I(N__62524));
    CascadeMux I__14514 (
            .O(N__62557),
            .I(N__62520));
    InMux I__14513 (
            .O(N__62556),
            .I(N__62515));
    InMux I__14512 (
            .O(N__62553),
            .I(N__62512));
    InMux I__14511 (
            .O(N__62552),
            .I(N__62507));
    InMux I__14510 (
            .O(N__62551),
            .I(N__62507));
    InMux I__14509 (
            .O(N__62550),
            .I(N__62499));
    Span4Mux_v I__14508 (
            .O(N__62547),
            .I(N__62496));
    Span4Mux_v I__14507 (
            .O(N__62544),
            .I(N__62493));
    InMux I__14506 (
            .O(N__62541),
            .I(N__62490));
    LocalMux I__14505 (
            .O(N__62538),
            .I(N__62487));
    LocalMux I__14504 (
            .O(N__62535),
            .I(N__62482));
    LocalMux I__14503 (
            .O(N__62530),
            .I(N__62482));
    Span4Mux_v I__14502 (
            .O(N__62527),
            .I(N__62479));
    LocalMux I__14501 (
            .O(N__62524),
            .I(N__62476));
    InMux I__14500 (
            .O(N__62523),
            .I(N__62473));
    InMux I__14499 (
            .O(N__62520),
            .I(N__62468));
    InMux I__14498 (
            .O(N__62519),
            .I(N__62468));
    InMux I__14497 (
            .O(N__62518),
            .I(N__62465));
    LocalMux I__14496 (
            .O(N__62515),
            .I(N__62462));
    LocalMux I__14495 (
            .O(N__62512),
            .I(N__62459));
    LocalMux I__14494 (
            .O(N__62507),
            .I(N__62456));
    InMux I__14493 (
            .O(N__62506),
            .I(N__62447));
    InMux I__14492 (
            .O(N__62505),
            .I(N__62447));
    InMux I__14491 (
            .O(N__62504),
            .I(N__62447));
    InMux I__14490 (
            .O(N__62503),
            .I(N__62447));
    InMux I__14489 (
            .O(N__62502),
            .I(N__62444));
    LocalMux I__14488 (
            .O(N__62499),
            .I(N__62441));
    Span4Mux_v I__14487 (
            .O(N__62496),
            .I(N__62436));
    Span4Mux_h I__14486 (
            .O(N__62493),
            .I(N__62436));
    LocalMux I__14485 (
            .O(N__62490),
            .I(N__62433));
    Span4Mux_v I__14484 (
            .O(N__62487),
            .I(N__62430));
    Span4Mux_h I__14483 (
            .O(N__62482),
            .I(N__62427));
    Span4Mux_h I__14482 (
            .O(N__62479),
            .I(N__62422));
    Span4Mux_v I__14481 (
            .O(N__62476),
            .I(N__62422));
    LocalMux I__14480 (
            .O(N__62473),
            .I(N__62417));
    LocalMux I__14479 (
            .O(N__62468),
            .I(N__62417));
    LocalMux I__14478 (
            .O(N__62465),
            .I(N__62414));
    Span4Mux_v I__14477 (
            .O(N__62462),
            .I(N__62411));
    Span4Mux_h I__14476 (
            .O(N__62459),
            .I(N__62402));
    Span4Mux_v I__14475 (
            .O(N__62456),
            .I(N__62402));
    LocalMux I__14474 (
            .O(N__62447),
            .I(N__62402));
    LocalMux I__14473 (
            .O(N__62444),
            .I(N__62402));
    Span12Mux_h I__14472 (
            .O(N__62441),
            .I(N__62399));
    Span4Mux_h I__14471 (
            .O(N__62436),
            .I(N__62392));
    Span4Mux_h I__14470 (
            .O(N__62433),
            .I(N__62392));
    Span4Mux_v I__14469 (
            .O(N__62430),
            .I(N__62392));
    Span4Mux_v I__14468 (
            .O(N__62427),
            .I(N__62389));
    Span4Mux_h I__14467 (
            .O(N__62422),
            .I(N__62382));
    Span4Mux_v I__14466 (
            .O(N__62417),
            .I(N__62382));
    Span4Mux_h I__14465 (
            .O(N__62414),
            .I(N__62382));
    Span4Mux_v I__14464 (
            .O(N__62411),
            .I(N__62377));
    Span4Mux_v I__14463 (
            .O(N__62402),
            .I(N__62377));
    Odrv12 I__14462 (
            .O(N__62399),
            .I(aluOut_6));
    Odrv4 I__14461 (
            .O(N__62392),
            .I(aluOut_6));
    Odrv4 I__14460 (
            .O(N__62389),
            .I(aluOut_6));
    Odrv4 I__14459 (
            .O(N__62382),
            .I(aluOut_6));
    Odrv4 I__14458 (
            .O(N__62377),
            .I(aluOut_6));
    CascadeMux I__14457 (
            .O(N__62366),
            .I(N__62363));
    InMux I__14456 (
            .O(N__62363),
            .I(N__62360));
    LocalMux I__14455 (
            .O(N__62360),
            .I(N__62357));
    Span4Mux_v I__14454 (
            .O(N__62357),
            .I(N__62354));
    Span4Mux_h I__14453 (
            .O(N__62354),
            .I(N__62351));
    Sp12to4 I__14452 (
            .O(N__62351),
            .I(N__62348));
    Odrv12 I__14451 (
            .O(N__62348),
            .I(\ALU.d_RNIALE3IZ0Z_6 ));
    InMux I__14450 (
            .O(N__62345),
            .I(N__62342));
    LocalMux I__14449 (
            .O(N__62342),
            .I(N__62339));
    Span4Mux_h I__14448 (
            .O(N__62339),
            .I(N__62335));
    InMux I__14447 (
            .O(N__62338),
            .I(N__62332));
    Odrv4 I__14446 (
            .O(N__62335),
            .I(\ALU.addsub_6 ));
    LocalMux I__14445 (
            .O(N__62332),
            .I(\ALU.addsub_6 ));
    InMux I__14444 (
            .O(N__62327),
            .I(\ALU.addsub_cry_5 ));
    CascadeMux I__14443 (
            .O(N__62324),
            .I(N__62321));
    InMux I__14442 (
            .O(N__62321),
            .I(N__62317));
    CascadeMux I__14441 (
            .O(N__62320),
            .I(N__62311));
    LocalMux I__14440 (
            .O(N__62317),
            .I(N__62308));
    CascadeMux I__14439 (
            .O(N__62316),
            .I(N__62303));
    CascadeMux I__14438 (
            .O(N__62315),
            .I(N__62299));
    InMux I__14437 (
            .O(N__62314),
            .I(N__62295));
    InMux I__14436 (
            .O(N__62311),
            .I(N__62292));
    Span4Mux_v I__14435 (
            .O(N__62308),
            .I(N__62289));
    InMux I__14434 (
            .O(N__62307),
            .I(N__62286));
    CascadeMux I__14433 (
            .O(N__62306),
            .I(N__62282));
    InMux I__14432 (
            .O(N__62303),
            .I(N__62278));
    CascadeMux I__14431 (
            .O(N__62302),
            .I(N__62275));
    InMux I__14430 (
            .O(N__62299),
            .I(N__62266));
    InMux I__14429 (
            .O(N__62298),
            .I(N__62262));
    LocalMux I__14428 (
            .O(N__62295),
            .I(N__62256));
    LocalMux I__14427 (
            .O(N__62292),
            .I(N__62256));
    Span4Mux_h I__14426 (
            .O(N__62289),
            .I(N__62251));
    LocalMux I__14425 (
            .O(N__62286),
            .I(N__62251));
    InMux I__14424 (
            .O(N__62285),
            .I(N__62244));
    InMux I__14423 (
            .O(N__62282),
            .I(N__62244));
    InMux I__14422 (
            .O(N__62281),
            .I(N__62244));
    LocalMux I__14421 (
            .O(N__62278),
            .I(N__62241));
    InMux I__14420 (
            .O(N__62275),
            .I(N__62238));
    InMux I__14419 (
            .O(N__62274),
            .I(N__62235));
    InMux I__14418 (
            .O(N__62273),
            .I(N__62223));
    InMux I__14417 (
            .O(N__62272),
            .I(N__62223));
    InMux I__14416 (
            .O(N__62271),
            .I(N__62223));
    InMux I__14415 (
            .O(N__62270),
            .I(N__62223));
    InMux I__14414 (
            .O(N__62269),
            .I(N__62220));
    LocalMux I__14413 (
            .O(N__62266),
            .I(N__62216));
    InMux I__14412 (
            .O(N__62265),
            .I(N__62213));
    LocalMux I__14411 (
            .O(N__62262),
            .I(N__62210));
    InMux I__14410 (
            .O(N__62261),
            .I(N__62206));
    Span4Mux_v I__14409 (
            .O(N__62256),
            .I(N__62199));
    Span4Mux_h I__14408 (
            .O(N__62251),
            .I(N__62199));
    LocalMux I__14407 (
            .O(N__62244),
            .I(N__62199));
    Span4Mux_v I__14406 (
            .O(N__62241),
            .I(N__62192));
    LocalMux I__14405 (
            .O(N__62238),
            .I(N__62192));
    LocalMux I__14404 (
            .O(N__62235),
            .I(N__62192));
    CascadeMux I__14403 (
            .O(N__62234),
            .I(N__62187));
    InMux I__14402 (
            .O(N__62233),
            .I(N__62182));
    InMux I__14401 (
            .O(N__62232),
            .I(N__62179));
    LocalMux I__14400 (
            .O(N__62223),
            .I(N__62176));
    LocalMux I__14399 (
            .O(N__62220),
            .I(N__62173));
    InMux I__14398 (
            .O(N__62219),
            .I(N__62170));
    Span4Mux_v I__14397 (
            .O(N__62216),
            .I(N__62165));
    LocalMux I__14396 (
            .O(N__62213),
            .I(N__62165));
    Span4Mux_v I__14395 (
            .O(N__62210),
            .I(N__62162));
    InMux I__14394 (
            .O(N__62209),
            .I(N__62159));
    LocalMux I__14393 (
            .O(N__62206),
            .I(N__62151));
    Span4Mux_v I__14392 (
            .O(N__62199),
            .I(N__62151));
    Span4Mux_v I__14391 (
            .O(N__62192),
            .I(N__62148));
    InMux I__14390 (
            .O(N__62191),
            .I(N__62143));
    InMux I__14389 (
            .O(N__62190),
            .I(N__62143));
    InMux I__14388 (
            .O(N__62187),
            .I(N__62138));
    InMux I__14387 (
            .O(N__62186),
            .I(N__62138));
    InMux I__14386 (
            .O(N__62185),
            .I(N__62135));
    LocalMux I__14385 (
            .O(N__62182),
            .I(N__62132));
    LocalMux I__14384 (
            .O(N__62179),
            .I(N__62125));
    Span4Mux_h I__14383 (
            .O(N__62176),
            .I(N__62125));
    Span4Mux_v I__14382 (
            .O(N__62173),
            .I(N__62125));
    LocalMux I__14381 (
            .O(N__62170),
            .I(N__62122));
    Span4Mux_v I__14380 (
            .O(N__62165),
            .I(N__62119));
    Span4Mux_h I__14379 (
            .O(N__62162),
            .I(N__62114));
    LocalMux I__14378 (
            .O(N__62159),
            .I(N__62114));
    InMux I__14377 (
            .O(N__62158),
            .I(N__62107));
    InMux I__14376 (
            .O(N__62157),
            .I(N__62107));
    InMux I__14375 (
            .O(N__62156),
            .I(N__62107));
    Span4Mux_v I__14374 (
            .O(N__62151),
            .I(N__62100));
    Span4Mux_h I__14373 (
            .O(N__62148),
            .I(N__62100));
    LocalMux I__14372 (
            .O(N__62143),
            .I(N__62100));
    LocalMux I__14371 (
            .O(N__62138),
            .I(N__62095));
    LocalMux I__14370 (
            .O(N__62135),
            .I(N__62095));
    Span4Mux_v I__14369 (
            .O(N__62132),
            .I(N__62090));
    Span4Mux_h I__14368 (
            .O(N__62125),
            .I(N__62090));
    Span4Mux_h I__14367 (
            .O(N__62122),
            .I(N__62087));
    Span4Mux_h I__14366 (
            .O(N__62119),
            .I(N__62084));
    Span4Mux_v I__14365 (
            .O(N__62114),
            .I(N__62079));
    LocalMux I__14364 (
            .O(N__62107),
            .I(N__62079));
    Span4Mux_h I__14363 (
            .O(N__62100),
            .I(N__62076));
    Span12Mux_h I__14362 (
            .O(N__62095),
            .I(N__62071));
    Sp12to4 I__14361 (
            .O(N__62090),
            .I(N__62071));
    Odrv4 I__14360 (
            .O(N__62087),
            .I(aluOut_7));
    Odrv4 I__14359 (
            .O(N__62084),
            .I(aluOut_7));
    Odrv4 I__14358 (
            .O(N__62079),
            .I(aluOut_7));
    Odrv4 I__14357 (
            .O(N__62076),
            .I(aluOut_7));
    Odrv12 I__14356 (
            .O(N__62071),
            .I(aluOut_7));
    CascadeMux I__14355 (
            .O(N__62060),
            .I(N__62057));
    InMux I__14354 (
            .O(N__62057),
            .I(N__62054));
    LocalMux I__14353 (
            .O(N__62054),
            .I(N__62051));
    Odrv12 I__14352 (
            .O(N__62051),
            .I(\ALU.d_RNI500DGZ0Z_7 ));
    InMux I__14351 (
            .O(N__62048),
            .I(N__62044));
    InMux I__14350 (
            .O(N__62047),
            .I(N__62041));
    LocalMux I__14349 (
            .O(N__62044),
            .I(N__62038));
    LocalMux I__14348 (
            .O(N__62041),
            .I(N__62035));
    Odrv4 I__14347 (
            .O(N__62038),
            .I(\ALU.addsub_7 ));
    Odrv4 I__14346 (
            .O(N__62035),
            .I(\ALU.addsub_7 ));
    InMux I__14345 (
            .O(N__62030),
            .I(bfn_23_15_0_));
    InMux I__14344 (
            .O(N__62027),
            .I(N__62018));
    CascadeMux I__14343 (
            .O(N__62026),
            .I(N__62014));
    CascadeMux I__14342 (
            .O(N__62025),
            .I(N__62011));
    InMux I__14341 (
            .O(N__62024),
            .I(N__62007));
    InMux I__14340 (
            .O(N__62023),
            .I(N__62004));
    CascadeMux I__14339 (
            .O(N__62022),
            .I(N__62001));
    CascadeMux I__14338 (
            .O(N__62021),
            .I(N__61997));
    LocalMux I__14337 (
            .O(N__62018),
            .I(N__61994));
    InMux I__14336 (
            .O(N__62017),
            .I(N__61991));
    InMux I__14335 (
            .O(N__62014),
            .I(N__61984));
    InMux I__14334 (
            .O(N__62011),
            .I(N__61984));
    InMux I__14333 (
            .O(N__62010),
            .I(N__61984));
    LocalMux I__14332 (
            .O(N__62007),
            .I(N__61979));
    LocalMux I__14331 (
            .O(N__62004),
            .I(N__61972));
    InMux I__14330 (
            .O(N__62001),
            .I(N__61969));
    CascadeMux I__14329 (
            .O(N__62000),
            .I(N__61966));
    InMux I__14328 (
            .O(N__61997),
            .I(N__61963));
    Span4Mux_h I__14327 (
            .O(N__61994),
            .I(N__61960));
    LocalMux I__14326 (
            .O(N__61991),
            .I(N__61955));
    LocalMux I__14325 (
            .O(N__61984),
            .I(N__61955));
    InMux I__14324 (
            .O(N__61983),
            .I(N__61952));
    CascadeMux I__14323 (
            .O(N__61982),
            .I(N__61949));
    Span4Mux_h I__14322 (
            .O(N__61979),
            .I(N__61944));
    InMux I__14321 (
            .O(N__61978),
            .I(N__61939));
    InMux I__14320 (
            .O(N__61977),
            .I(N__61939));
    CascadeMux I__14319 (
            .O(N__61976),
            .I(N__61936));
    CascadeMux I__14318 (
            .O(N__61975),
            .I(N__61932));
    Span4Mux_h I__14317 (
            .O(N__61972),
            .I(N__61925));
    LocalMux I__14316 (
            .O(N__61969),
            .I(N__61925));
    InMux I__14315 (
            .O(N__61966),
            .I(N__61922));
    LocalMux I__14314 (
            .O(N__61963),
            .I(N__61919));
    Span4Mux_v I__14313 (
            .O(N__61960),
            .I(N__61914));
    Span4Mux_v I__14312 (
            .O(N__61955),
            .I(N__61914));
    LocalMux I__14311 (
            .O(N__61952),
            .I(N__61911));
    InMux I__14310 (
            .O(N__61949),
            .I(N__61908));
    CascadeMux I__14309 (
            .O(N__61948),
            .I(N__61905));
    InMux I__14308 (
            .O(N__61947),
            .I(N__61902));
    Span4Mux_h I__14307 (
            .O(N__61944),
            .I(N__61896));
    LocalMux I__14306 (
            .O(N__61939),
            .I(N__61896));
    InMux I__14305 (
            .O(N__61936),
            .I(N__61893));
    InMux I__14304 (
            .O(N__61935),
            .I(N__61890));
    InMux I__14303 (
            .O(N__61932),
            .I(N__61887));
    InMux I__14302 (
            .O(N__61931),
            .I(N__61882));
    InMux I__14301 (
            .O(N__61930),
            .I(N__61882));
    Span4Mux_h I__14300 (
            .O(N__61925),
            .I(N__61878));
    LocalMux I__14299 (
            .O(N__61922),
            .I(N__61869));
    Span4Mux_h I__14298 (
            .O(N__61919),
            .I(N__61869));
    Span4Mux_h I__14297 (
            .O(N__61914),
            .I(N__61869));
    Span4Mux_v I__14296 (
            .O(N__61911),
            .I(N__61869));
    LocalMux I__14295 (
            .O(N__61908),
            .I(N__61866));
    InMux I__14294 (
            .O(N__61905),
            .I(N__61863));
    LocalMux I__14293 (
            .O(N__61902),
            .I(N__61860));
    InMux I__14292 (
            .O(N__61901),
            .I(N__61857));
    Span4Mux_h I__14291 (
            .O(N__61896),
            .I(N__61852));
    LocalMux I__14290 (
            .O(N__61893),
            .I(N__61852));
    LocalMux I__14289 (
            .O(N__61890),
            .I(N__61849));
    LocalMux I__14288 (
            .O(N__61887),
            .I(N__61846));
    LocalMux I__14287 (
            .O(N__61882),
            .I(N__61843));
    InMux I__14286 (
            .O(N__61881),
            .I(N__61840));
    Span4Mux_v I__14285 (
            .O(N__61878),
            .I(N__61837));
    Span4Mux_h I__14284 (
            .O(N__61869),
            .I(N__61833));
    Span4Mux_h I__14283 (
            .O(N__61866),
            .I(N__61830));
    LocalMux I__14282 (
            .O(N__61863),
            .I(N__61827));
    Span4Mux_h I__14281 (
            .O(N__61860),
            .I(N__61820));
    LocalMux I__14280 (
            .O(N__61857),
            .I(N__61820));
    Span4Mux_v I__14279 (
            .O(N__61852),
            .I(N__61820));
    Span12Mux_v I__14278 (
            .O(N__61849),
            .I(N__61817));
    Span4Mux_v I__14277 (
            .O(N__61846),
            .I(N__61812));
    Span4Mux_h I__14276 (
            .O(N__61843),
            .I(N__61812));
    LocalMux I__14275 (
            .O(N__61840),
            .I(N__61807));
    Span4Mux_v I__14274 (
            .O(N__61837),
            .I(N__61807));
    InMux I__14273 (
            .O(N__61836),
            .I(N__61804));
    Span4Mux_v I__14272 (
            .O(N__61833),
            .I(N__61799));
    Span4Mux_h I__14271 (
            .O(N__61830),
            .I(N__61799));
    Span4Mux_h I__14270 (
            .O(N__61827),
            .I(N__61794));
    Span4Mux_v I__14269 (
            .O(N__61820),
            .I(N__61794));
    Odrv12 I__14268 (
            .O(N__61817),
            .I(aluOut_8));
    Odrv4 I__14267 (
            .O(N__61812),
            .I(aluOut_8));
    Odrv4 I__14266 (
            .O(N__61807),
            .I(aluOut_8));
    LocalMux I__14265 (
            .O(N__61804),
            .I(aluOut_8));
    Odrv4 I__14264 (
            .O(N__61799),
            .I(aluOut_8));
    Odrv4 I__14263 (
            .O(N__61794),
            .I(aluOut_8));
    CascadeMux I__14262 (
            .O(N__61781),
            .I(N__61778));
    InMux I__14261 (
            .O(N__61778),
            .I(N__61775));
    LocalMux I__14260 (
            .O(N__61775),
            .I(N__61772));
    Span4Mux_h I__14259 (
            .O(N__61772),
            .I(N__61769));
    Span4Mux_v I__14258 (
            .O(N__61769),
            .I(N__61766));
    Span4Mux_h I__14257 (
            .O(N__61766),
            .I(N__61763));
    Odrv4 I__14256 (
            .O(N__61763),
            .I(\ALU.d_RNIAJ1KHZ0Z_8 ));
    InMux I__14255 (
            .O(N__61760),
            .I(N__61757));
    LocalMux I__14254 (
            .O(N__61757),
            .I(N__61754));
    Span4Mux_v I__14253 (
            .O(N__61754),
            .I(N__61750));
    InMux I__14252 (
            .O(N__61753),
            .I(N__61747));
    Odrv4 I__14251 (
            .O(N__61750),
            .I(\ALU.addsub_8 ));
    LocalMux I__14250 (
            .O(N__61747),
            .I(\ALU.addsub_8 ));
    InMux I__14249 (
            .O(N__61742),
            .I(\ALU.addsub_cry_7 ));
    InMux I__14248 (
            .O(N__61739),
            .I(\ALU.addsub_cry_8 ));
    InMux I__14247 (
            .O(N__61736),
            .I(N__61733));
    LocalMux I__14246 (
            .O(N__61733),
            .I(N__61730));
    Span4Mux_v I__14245 (
            .O(N__61730),
            .I(N__61727));
    Sp12to4 I__14244 (
            .O(N__61727),
            .I(N__61724));
    Span12Mux_h I__14243 (
            .O(N__61724),
            .I(N__61721));
    Odrv12 I__14242 (
            .O(N__61721),
            .I(\ALU.c_RNI1QK5KZ0Z_10 ));
    CascadeMux I__14241 (
            .O(N__61718),
            .I(N__61711));
    CascadeMux I__14240 (
            .O(N__61717),
            .I(N__61707));
    CascadeMux I__14239 (
            .O(N__61716),
            .I(N__61704));
    CascadeMux I__14238 (
            .O(N__61715),
            .I(N__61698));
    InMux I__14237 (
            .O(N__61714),
            .I(N__61692));
    InMux I__14236 (
            .O(N__61711),
            .I(N__61692));
    CascadeMux I__14235 (
            .O(N__61710),
            .I(N__61689));
    InMux I__14234 (
            .O(N__61707),
            .I(N__61686));
    InMux I__14233 (
            .O(N__61704),
            .I(N__61683));
    InMux I__14232 (
            .O(N__61703),
            .I(N__61676));
    InMux I__14231 (
            .O(N__61702),
            .I(N__61676));
    InMux I__14230 (
            .O(N__61701),
            .I(N__61672));
    InMux I__14229 (
            .O(N__61698),
            .I(N__61669));
    InMux I__14228 (
            .O(N__61697),
            .I(N__61663));
    LocalMux I__14227 (
            .O(N__61692),
            .I(N__61658));
    InMux I__14226 (
            .O(N__61689),
            .I(N__61655));
    LocalMux I__14225 (
            .O(N__61686),
            .I(N__61650));
    LocalMux I__14224 (
            .O(N__61683),
            .I(N__61650));
    InMux I__14223 (
            .O(N__61682),
            .I(N__61647));
    InMux I__14222 (
            .O(N__61681),
            .I(N__61644));
    LocalMux I__14221 (
            .O(N__61676),
            .I(N__61641));
    CascadeMux I__14220 (
            .O(N__61675),
            .I(N__61637));
    LocalMux I__14219 (
            .O(N__61672),
            .I(N__61633));
    LocalMux I__14218 (
            .O(N__61669),
            .I(N__61630));
    CascadeMux I__14217 (
            .O(N__61668),
            .I(N__61627));
    InMux I__14216 (
            .O(N__61667),
            .I(N__61624));
    InMux I__14215 (
            .O(N__61666),
            .I(N__61621));
    LocalMux I__14214 (
            .O(N__61663),
            .I(N__61618));
    InMux I__14213 (
            .O(N__61662),
            .I(N__61613));
    InMux I__14212 (
            .O(N__61661),
            .I(N__61613));
    Span4Mux_v I__14211 (
            .O(N__61658),
            .I(N__61610));
    LocalMux I__14210 (
            .O(N__61655),
            .I(N__61607));
    Span4Mux_v I__14209 (
            .O(N__61650),
            .I(N__61604));
    LocalMux I__14208 (
            .O(N__61647),
            .I(N__61599));
    LocalMux I__14207 (
            .O(N__61644),
            .I(N__61599));
    Span4Mux_h I__14206 (
            .O(N__61641),
            .I(N__61596));
    InMux I__14205 (
            .O(N__61640),
            .I(N__61593));
    InMux I__14204 (
            .O(N__61637),
            .I(N__61588));
    InMux I__14203 (
            .O(N__61636),
            .I(N__61588));
    Span4Mux_v I__14202 (
            .O(N__61633),
            .I(N__61583));
    Span4Mux_v I__14201 (
            .O(N__61630),
            .I(N__61583));
    InMux I__14200 (
            .O(N__61627),
            .I(N__61580));
    LocalMux I__14199 (
            .O(N__61624),
            .I(N__61577));
    LocalMux I__14198 (
            .O(N__61621),
            .I(N__61574));
    Span4Mux_h I__14197 (
            .O(N__61618),
            .I(N__61571));
    LocalMux I__14196 (
            .O(N__61613),
            .I(N__61568));
    Sp12to4 I__14195 (
            .O(N__61610),
            .I(N__61565));
    Span4Mux_v I__14194 (
            .O(N__61607),
            .I(N__61562));
    Span4Mux_v I__14193 (
            .O(N__61604),
            .I(N__61559));
    Span4Mux_v I__14192 (
            .O(N__61599),
            .I(N__61556));
    Span4Mux_h I__14191 (
            .O(N__61596),
            .I(N__61553));
    LocalMux I__14190 (
            .O(N__61593),
            .I(N__61546));
    LocalMux I__14189 (
            .O(N__61588),
            .I(N__61546));
    Sp12to4 I__14188 (
            .O(N__61583),
            .I(N__61546));
    LocalMux I__14187 (
            .O(N__61580),
            .I(N__61541));
    Span4Mux_h I__14186 (
            .O(N__61577),
            .I(N__61541));
    Span4Mux_v I__14185 (
            .O(N__61574),
            .I(N__61536));
    Span4Mux_h I__14184 (
            .O(N__61571),
            .I(N__61536));
    Span4Mux_h I__14183 (
            .O(N__61568),
            .I(N__61533));
    Span12Mux_s11_h I__14182 (
            .O(N__61565),
            .I(N__61526));
    Sp12to4 I__14181 (
            .O(N__61562),
            .I(N__61526));
    Sp12to4 I__14180 (
            .O(N__61559),
            .I(N__61526));
    Span4Mux_h I__14179 (
            .O(N__61556),
            .I(N__61521));
    Span4Mux_v I__14178 (
            .O(N__61553),
            .I(N__61521));
    Span12Mux_h I__14177 (
            .O(N__61546),
            .I(N__61516));
    Sp12to4 I__14176 (
            .O(N__61541),
            .I(N__61516));
    Odrv4 I__14175 (
            .O(N__61536),
            .I(aluOut_10));
    Odrv4 I__14174 (
            .O(N__61533),
            .I(aluOut_10));
    Odrv12 I__14173 (
            .O(N__61526),
            .I(aluOut_10));
    Odrv4 I__14172 (
            .O(N__61521),
            .I(aluOut_10));
    Odrv12 I__14171 (
            .O(N__61516),
            .I(aluOut_10));
    InMux I__14170 (
            .O(N__61505),
            .I(N__61502));
    LocalMux I__14169 (
            .O(N__61502),
            .I(N__61499));
    Span4Mux_h I__14168 (
            .O(N__61499),
            .I(N__61496));
    Span4Mux_h I__14167 (
            .O(N__61496),
            .I(N__61493));
    Span4Mux_h I__14166 (
            .O(N__61493),
            .I(N__61489));
    InMux I__14165 (
            .O(N__61492),
            .I(N__61486));
    Span4Mux_v I__14164 (
            .O(N__61489),
            .I(N__61483));
    LocalMux I__14163 (
            .O(N__61486),
            .I(\ALU.addsub_10 ));
    Odrv4 I__14162 (
            .O(N__61483),
            .I(\ALU.addsub_10 ));
    InMux I__14161 (
            .O(N__61478),
            .I(\ALU.addsub_cry_9 ));
    InMux I__14160 (
            .O(N__61475),
            .I(N__61467));
    InMux I__14159 (
            .O(N__61474),
            .I(N__61457));
    InMux I__14158 (
            .O(N__61473),
            .I(N__61454));
    InMux I__14157 (
            .O(N__61472),
            .I(N__61447));
    InMux I__14156 (
            .O(N__61471),
            .I(N__61447));
    InMux I__14155 (
            .O(N__61470),
            .I(N__61447));
    LocalMux I__14154 (
            .O(N__61467),
            .I(N__61443));
    InMux I__14153 (
            .O(N__61466),
            .I(N__61440));
    InMux I__14152 (
            .O(N__61465),
            .I(N__61436));
    InMux I__14151 (
            .O(N__61464),
            .I(N__61428));
    InMux I__14150 (
            .O(N__61463),
            .I(N__61428));
    InMux I__14149 (
            .O(N__61462),
            .I(N__61422));
    InMux I__14148 (
            .O(N__61461),
            .I(N__61417));
    InMux I__14147 (
            .O(N__61460),
            .I(N__61417));
    LocalMux I__14146 (
            .O(N__61457),
            .I(N__61410));
    LocalMux I__14145 (
            .O(N__61454),
            .I(N__61410));
    LocalMux I__14144 (
            .O(N__61447),
            .I(N__61410));
    InMux I__14143 (
            .O(N__61446),
            .I(N__61407));
    Span4Mux_v I__14142 (
            .O(N__61443),
            .I(N__61404));
    LocalMux I__14141 (
            .O(N__61440),
            .I(N__61401));
    InMux I__14140 (
            .O(N__61439),
            .I(N__61398));
    LocalMux I__14139 (
            .O(N__61436),
            .I(N__61395));
    InMux I__14138 (
            .O(N__61435),
            .I(N__61390));
    InMux I__14137 (
            .O(N__61434),
            .I(N__61390));
    InMux I__14136 (
            .O(N__61433),
            .I(N__61387));
    LocalMux I__14135 (
            .O(N__61428),
            .I(N__61384));
    InMux I__14134 (
            .O(N__61427),
            .I(N__61381));
    InMux I__14133 (
            .O(N__61426),
            .I(N__61378));
    InMux I__14132 (
            .O(N__61425),
            .I(N__61375));
    LocalMux I__14131 (
            .O(N__61422),
            .I(N__61372));
    LocalMux I__14130 (
            .O(N__61417),
            .I(N__61365));
    Span4Mux_v I__14129 (
            .O(N__61410),
            .I(N__61365));
    LocalMux I__14128 (
            .O(N__61407),
            .I(N__61365));
    Span4Mux_h I__14127 (
            .O(N__61404),
            .I(N__61353));
    Span4Mux_v I__14126 (
            .O(N__61401),
            .I(N__61353));
    LocalMux I__14125 (
            .O(N__61398),
            .I(N__61353));
    Span4Mux_v I__14124 (
            .O(N__61395),
            .I(N__61353));
    LocalMux I__14123 (
            .O(N__61390),
            .I(N__61353));
    LocalMux I__14122 (
            .O(N__61387),
            .I(N__61350));
    Span4Mux_h I__14121 (
            .O(N__61384),
            .I(N__61347));
    LocalMux I__14120 (
            .O(N__61381),
            .I(N__61344));
    LocalMux I__14119 (
            .O(N__61378),
            .I(N__61341));
    LocalMux I__14118 (
            .O(N__61375),
            .I(N__61334));
    Span4Mux_v I__14117 (
            .O(N__61372),
            .I(N__61334));
    Span4Mux_h I__14116 (
            .O(N__61365),
            .I(N__61334));
    InMux I__14115 (
            .O(N__61364),
            .I(N__61331));
    Span4Mux_v I__14114 (
            .O(N__61353),
            .I(N__61328));
    Span4Mux_v I__14113 (
            .O(N__61350),
            .I(N__61325));
    Span4Mux_h I__14112 (
            .O(N__61347),
            .I(N__61322));
    Span4Mux_h I__14111 (
            .O(N__61344),
            .I(N__61317));
    Span4Mux_v I__14110 (
            .O(N__61341),
            .I(N__61317));
    Span4Mux_h I__14109 (
            .O(N__61334),
            .I(N__61314));
    LocalMux I__14108 (
            .O(N__61331),
            .I(N__61309));
    Sp12to4 I__14107 (
            .O(N__61328),
            .I(N__61309));
    Odrv4 I__14106 (
            .O(N__61325),
            .I(aluOut_11));
    Odrv4 I__14105 (
            .O(N__61322),
            .I(aluOut_11));
    Odrv4 I__14104 (
            .O(N__61317),
            .I(aluOut_11));
    Odrv4 I__14103 (
            .O(N__61314),
            .I(aluOut_11));
    Odrv12 I__14102 (
            .O(N__61309),
            .I(aluOut_11));
    CascadeMux I__14101 (
            .O(N__61298),
            .I(N__61295));
    InMux I__14100 (
            .O(N__61295),
            .I(N__61292));
    LocalMux I__14099 (
            .O(N__61292),
            .I(N__61289));
    Span4Mux_v I__14098 (
            .O(N__61289),
            .I(N__61286));
    Sp12to4 I__14097 (
            .O(N__61286),
            .I(N__61283));
    Span12Mux_h I__14096 (
            .O(N__61283),
            .I(N__61280));
    Odrv12 I__14095 (
            .O(N__61280),
            .I(\ALU.c_RNIRRB4IZ0Z_11 ));
    InMux I__14094 (
            .O(N__61277),
            .I(N__61273));
    InMux I__14093 (
            .O(N__61276),
            .I(N__61270));
    LocalMux I__14092 (
            .O(N__61273),
            .I(N__61267));
    LocalMux I__14091 (
            .O(N__61270),
            .I(N__61264));
    Span4Mux_v I__14090 (
            .O(N__61267),
            .I(N__61261));
    Span4Mux_h I__14089 (
            .O(N__61264),
            .I(N__61258));
    Span4Mux_h I__14088 (
            .O(N__61261),
            .I(N__61255));
    Span4Mux_h I__14087 (
            .O(N__61258),
            .I(N__61252));
    Odrv4 I__14086 (
            .O(N__61255),
            .I(\ALU.addsub_11 ));
    Odrv4 I__14085 (
            .O(N__61252),
            .I(\ALU.addsub_11 ));
    InMux I__14084 (
            .O(N__61247),
            .I(\ALU.addsub_cry_10 ));
    InMux I__14083 (
            .O(N__61244),
            .I(N__61241));
    LocalMux I__14082 (
            .O(N__61241),
            .I(N__61238));
    Span4Mux_h I__14081 (
            .O(N__61238),
            .I(N__61235));
    Span4Mux_v I__14080 (
            .O(N__61235),
            .I(N__61232));
    Span4Mux_h I__14079 (
            .O(N__61232),
            .I(N__61229));
    Odrv4 I__14078 (
            .O(N__61229),
            .I(\ALU.c_RNITVOEKZ0Z_12 ));
    InMux I__14077 (
            .O(N__61226),
            .I(N__61221));
    CascadeMux I__14076 (
            .O(N__61225),
            .I(N__61218));
    CascadeMux I__14075 (
            .O(N__61224),
            .I(N__61213));
    LocalMux I__14074 (
            .O(N__61221),
            .I(N__61207));
    InMux I__14073 (
            .O(N__61218),
            .I(N__61204));
    CascadeMux I__14072 (
            .O(N__61217),
            .I(N__61200));
    CascadeMux I__14071 (
            .O(N__61216),
            .I(N__61196));
    InMux I__14070 (
            .O(N__61213),
            .I(N__61190));
    InMux I__14069 (
            .O(N__61212),
            .I(N__61187));
    InMux I__14068 (
            .O(N__61211),
            .I(N__61184));
    CascadeMux I__14067 (
            .O(N__61210),
            .I(N__61181));
    Span4Mux_v I__14066 (
            .O(N__61207),
            .I(N__61176));
    LocalMux I__14065 (
            .O(N__61204),
            .I(N__61176));
    InMux I__14064 (
            .O(N__61203),
            .I(N__61171));
    InMux I__14063 (
            .O(N__61200),
            .I(N__61171));
    InMux I__14062 (
            .O(N__61199),
            .I(N__61167));
    InMux I__14061 (
            .O(N__61196),
            .I(N__61164));
    InMux I__14060 (
            .O(N__61195),
            .I(N__61161));
    CascadeMux I__14059 (
            .O(N__61194),
            .I(N__61158));
    InMux I__14058 (
            .O(N__61193),
            .I(N__61153));
    LocalMux I__14057 (
            .O(N__61190),
            .I(N__61148));
    LocalMux I__14056 (
            .O(N__61187),
            .I(N__61143));
    LocalMux I__14055 (
            .O(N__61184),
            .I(N__61143));
    InMux I__14054 (
            .O(N__61181),
            .I(N__61140));
    Span4Mux_h I__14053 (
            .O(N__61176),
            .I(N__61135));
    LocalMux I__14052 (
            .O(N__61171),
            .I(N__61135));
    InMux I__14051 (
            .O(N__61170),
            .I(N__61132));
    LocalMux I__14050 (
            .O(N__61167),
            .I(N__61129));
    LocalMux I__14049 (
            .O(N__61164),
            .I(N__61126));
    LocalMux I__14048 (
            .O(N__61161),
            .I(N__61123));
    InMux I__14047 (
            .O(N__61158),
            .I(N__61120));
    InMux I__14046 (
            .O(N__61157),
            .I(N__61115));
    InMux I__14045 (
            .O(N__61156),
            .I(N__61115));
    LocalMux I__14044 (
            .O(N__61153),
            .I(N__61112));
    InMux I__14043 (
            .O(N__61152),
            .I(N__61107));
    InMux I__14042 (
            .O(N__61151),
            .I(N__61107));
    Span4Mux_v I__14041 (
            .O(N__61148),
            .I(N__61104));
    Span4Mux_v I__14040 (
            .O(N__61143),
            .I(N__61101));
    LocalMux I__14039 (
            .O(N__61140),
            .I(N__61094));
    Span4Mux_h I__14038 (
            .O(N__61135),
            .I(N__61094));
    LocalMux I__14037 (
            .O(N__61132),
            .I(N__61094));
    Span4Mux_h I__14036 (
            .O(N__61129),
            .I(N__61091));
    Span4Mux_v I__14035 (
            .O(N__61126),
            .I(N__61082));
    Span4Mux_v I__14034 (
            .O(N__61123),
            .I(N__61082));
    LocalMux I__14033 (
            .O(N__61120),
            .I(N__61082));
    LocalMux I__14032 (
            .O(N__61115),
            .I(N__61082));
    Span4Mux_v I__14031 (
            .O(N__61112),
            .I(N__61079));
    LocalMux I__14030 (
            .O(N__61107),
            .I(N__61076));
    Span4Mux_h I__14029 (
            .O(N__61104),
            .I(N__61071));
    Span4Mux_v I__14028 (
            .O(N__61101),
            .I(N__61071));
    Span4Mux_v I__14027 (
            .O(N__61094),
            .I(N__61068));
    Span4Mux_v I__14026 (
            .O(N__61091),
            .I(N__61063));
    Span4Mux_h I__14025 (
            .O(N__61082),
            .I(N__61063));
    Span4Mux_h I__14024 (
            .O(N__61079),
            .I(N__61058));
    Span4Mux_h I__14023 (
            .O(N__61076),
            .I(N__61058));
    Span4Mux_h I__14022 (
            .O(N__61071),
            .I(N__61053));
    Span4Mux_v I__14021 (
            .O(N__61068),
            .I(N__61053));
    Span4Mux_v I__14020 (
            .O(N__61063),
            .I(N__61050));
    Odrv4 I__14019 (
            .O(N__61058),
            .I(aluOut_12));
    Odrv4 I__14018 (
            .O(N__61053),
            .I(aluOut_12));
    Odrv4 I__14017 (
            .O(N__61050),
            .I(aluOut_12));
    InMux I__14016 (
            .O(N__61043),
            .I(N__61037));
    InMux I__14015 (
            .O(N__61042),
            .I(N__61037));
    LocalMux I__14014 (
            .O(N__61037),
            .I(N__61034));
    Span4Mux_v I__14013 (
            .O(N__61034),
            .I(N__61031));
    Odrv4 I__14012 (
            .O(N__61031),
            .I(\ALU.addsub_12 ));
    InMux I__14011 (
            .O(N__61028),
            .I(\ALU.addsub_cry_11 ));
    InMux I__14010 (
            .O(N__61025),
            .I(N__61022));
    LocalMux I__14009 (
            .O(N__61022),
            .I(\ALU.c_RNIVHVMKZ0Z_13 ));
    CascadeMux I__14008 (
            .O(N__61019),
            .I(N__61015));
    InMux I__14007 (
            .O(N__61018),
            .I(N__61005));
    InMux I__14006 (
            .O(N__61015),
            .I(N__61002));
    InMux I__14005 (
            .O(N__61014),
            .I(N__60999));
    CascadeMux I__14004 (
            .O(N__61013),
            .I(N__60996));
    InMux I__14003 (
            .O(N__61012),
            .I(N__60991));
    InMux I__14002 (
            .O(N__61011),
            .I(N__60987));
    InMux I__14001 (
            .O(N__61010),
            .I(N__60984));
    InMux I__14000 (
            .O(N__61009),
            .I(N__60979));
    InMux I__13999 (
            .O(N__61008),
            .I(N__60979));
    LocalMux I__13998 (
            .O(N__61005),
            .I(N__60972));
    LocalMux I__13997 (
            .O(N__61002),
            .I(N__60972));
    LocalMux I__13996 (
            .O(N__60999),
            .I(N__60972));
    InMux I__13995 (
            .O(N__60996),
            .I(N__60969));
    InMux I__13994 (
            .O(N__60995),
            .I(N__60966));
    InMux I__13993 (
            .O(N__60994),
            .I(N__60961));
    LocalMux I__13992 (
            .O(N__60991),
            .I(N__60958));
    InMux I__13991 (
            .O(N__60990),
            .I(N__60955));
    LocalMux I__13990 (
            .O(N__60987),
            .I(N__60950));
    LocalMux I__13989 (
            .O(N__60984),
            .I(N__60947));
    LocalMux I__13988 (
            .O(N__60979),
            .I(N__60944));
    Span4Mux_h I__13987 (
            .O(N__60972),
            .I(N__60941));
    LocalMux I__13986 (
            .O(N__60969),
            .I(N__60933));
    LocalMux I__13985 (
            .O(N__60966),
            .I(N__60933));
    InMux I__13984 (
            .O(N__60965),
            .I(N__60928));
    InMux I__13983 (
            .O(N__60964),
            .I(N__60928));
    LocalMux I__13982 (
            .O(N__60961),
            .I(N__60925));
    Span4Mux_v I__13981 (
            .O(N__60958),
            .I(N__60920));
    LocalMux I__13980 (
            .O(N__60955),
            .I(N__60920));
    InMux I__13979 (
            .O(N__60954),
            .I(N__60917));
    InMux I__13978 (
            .O(N__60953),
            .I(N__60914));
    Span4Mux_v I__13977 (
            .O(N__60950),
            .I(N__60911));
    Span4Mux_v I__13976 (
            .O(N__60947),
            .I(N__60906));
    Span4Mux_v I__13975 (
            .O(N__60944),
            .I(N__60906));
    Span4Mux_v I__13974 (
            .O(N__60941),
            .I(N__60903));
    InMux I__13973 (
            .O(N__60940),
            .I(N__60896));
    InMux I__13972 (
            .O(N__60939),
            .I(N__60896));
    InMux I__13971 (
            .O(N__60938),
            .I(N__60896));
    Span4Mux_v I__13970 (
            .O(N__60933),
            .I(N__60893));
    LocalMux I__13969 (
            .O(N__60928),
            .I(N__60890));
    Span4Mux_v I__13968 (
            .O(N__60925),
            .I(N__60887));
    Span4Mux_v I__13967 (
            .O(N__60920),
            .I(N__60884));
    LocalMux I__13966 (
            .O(N__60917),
            .I(N__60879));
    LocalMux I__13965 (
            .O(N__60914),
            .I(N__60879));
    Sp12to4 I__13964 (
            .O(N__60911),
            .I(N__60870));
    Sp12to4 I__13963 (
            .O(N__60906),
            .I(N__60870));
    Sp12to4 I__13962 (
            .O(N__60903),
            .I(N__60870));
    LocalMux I__13961 (
            .O(N__60896),
            .I(N__60870));
    Span4Mux_v I__13960 (
            .O(N__60893),
            .I(N__60867));
    Span4Mux_v I__13959 (
            .O(N__60890),
            .I(N__60864));
    Span4Mux_v I__13958 (
            .O(N__60887),
            .I(N__60861));
    Span4Mux_v I__13957 (
            .O(N__60884),
            .I(N__60858));
    Sp12to4 I__13956 (
            .O(N__60879),
            .I(N__60853));
    Span12Mux_h I__13955 (
            .O(N__60870),
            .I(N__60853));
    Span4Mux_h I__13954 (
            .O(N__60867),
            .I(N__60848));
    Span4Mux_v I__13953 (
            .O(N__60864),
            .I(N__60848));
    Odrv4 I__13952 (
            .O(N__60861),
            .I(aluOut_13));
    Odrv4 I__13951 (
            .O(N__60858),
            .I(aluOut_13));
    Odrv12 I__13950 (
            .O(N__60853),
            .I(aluOut_13));
    Odrv4 I__13949 (
            .O(N__60848),
            .I(aluOut_13));
    InMux I__13948 (
            .O(N__60839),
            .I(N__60836));
    LocalMux I__13947 (
            .O(N__60836),
            .I(N__60832));
    InMux I__13946 (
            .O(N__60835),
            .I(N__60829));
    Span4Mux_h I__13945 (
            .O(N__60832),
            .I(N__60826));
    LocalMux I__13944 (
            .O(N__60829),
            .I(N__60823));
    Odrv4 I__13943 (
            .O(N__60826),
            .I(\ALU.addsub_13 ));
    Odrv12 I__13942 (
            .O(N__60823),
            .I(\ALU.addsub_13 ));
    CascadeMux I__13941 (
            .O(N__60818),
            .I(N__60815));
    InMux I__13940 (
            .O(N__60815),
            .I(N__60809));
    CascadeMux I__13939 (
            .O(N__60814),
            .I(N__60806));
    InMux I__13938 (
            .O(N__60813),
            .I(N__60802));
    CascadeMux I__13937 (
            .O(N__60812),
            .I(N__60799));
    LocalMux I__13936 (
            .O(N__60809),
            .I(N__60796));
    InMux I__13935 (
            .O(N__60806),
            .I(N__60793));
    CascadeMux I__13934 (
            .O(N__60805),
            .I(N__60790));
    LocalMux I__13933 (
            .O(N__60802),
            .I(N__60787));
    InMux I__13932 (
            .O(N__60799),
            .I(N__60784));
    Sp12to4 I__13931 (
            .O(N__60796),
            .I(N__60781));
    LocalMux I__13930 (
            .O(N__60793),
            .I(N__60777));
    InMux I__13929 (
            .O(N__60790),
            .I(N__60774));
    Span4Mux_v I__13928 (
            .O(N__60787),
            .I(N__60769));
    LocalMux I__13927 (
            .O(N__60784),
            .I(N__60769));
    Span12Mux_v I__13926 (
            .O(N__60781),
            .I(N__60766));
    InMux I__13925 (
            .O(N__60780),
            .I(N__60763));
    Span4Mux_v I__13924 (
            .O(N__60777),
            .I(N__60760));
    LocalMux I__13923 (
            .O(N__60774),
            .I(N__60755));
    Span4Mux_h I__13922 (
            .O(N__60769),
            .I(N__60755));
    Span12Mux_h I__13921 (
            .O(N__60766),
            .I(N__60752));
    LocalMux I__13920 (
            .O(N__60763),
            .I(\CONTROL.addrstackptrZ0Z_4 ));
    Odrv4 I__13919 (
            .O(N__60760),
            .I(\CONTROL.addrstackptrZ0Z_4 ));
    Odrv4 I__13918 (
            .O(N__60755),
            .I(\CONTROL.addrstackptrZ0Z_4 ));
    Odrv12 I__13917 (
            .O(N__60752),
            .I(\CONTROL.addrstackptrZ0Z_4 ));
    CascadeMux I__13916 (
            .O(N__60743),
            .I(N__60740));
    InMux I__13915 (
            .O(N__60740),
            .I(N__60737));
    LocalMux I__13914 (
            .O(N__60737),
            .I(N__60731));
    InMux I__13913 (
            .O(N__60736),
            .I(N__60727));
    CascadeMux I__13912 (
            .O(N__60735),
            .I(N__60724));
    CascadeMux I__13911 (
            .O(N__60734),
            .I(N__60720));
    Span4Mux_v I__13910 (
            .O(N__60731),
            .I(N__60717));
    InMux I__13909 (
            .O(N__60730),
            .I(N__60714));
    LocalMux I__13908 (
            .O(N__60727),
            .I(N__60711));
    InMux I__13907 (
            .O(N__60724),
            .I(N__60708));
    InMux I__13906 (
            .O(N__60723),
            .I(N__60705));
    InMux I__13905 (
            .O(N__60720),
            .I(N__60702));
    Span4Mux_h I__13904 (
            .O(N__60717),
            .I(N__60696));
    LocalMux I__13903 (
            .O(N__60714),
            .I(N__60696));
    Span4Mux_h I__13902 (
            .O(N__60711),
            .I(N__60693));
    LocalMux I__13901 (
            .O(N__60708),
            .I(N__60686));
    LocalMux I__13900 (
            .O(N__60705),
            .I(N__60686));
    LocalMux I__13899 (
            .O(N__60702),
            .I(N__60686));
    CascadeMux I__13898 (
            .O(N__60701),
            .I(N__60683));
    Sp12to4 I__13897 (
            .O(N__60696),
            .I(N__60679));
    Sp12to4 I__13896 (
            .O(N__60693),
            .I(N__60676));
    Span4Mux_v I__13895 (
            .O(N__60686),
            .I(N__60673));
    InMux I__13894 (
            .O(N__60683),
            .I(N__60668));
    InMux I__13893 (
            .O(N__60682),
            .I(N__60668));
    Span12Mux_h I__13892 (
            .O(N__60679),
            .I(N__60663));
    Span12Mux_v I__13891 (
            .O(N__60676),
            .I(N__60663));
    Sp12to4 I__13890 (
            .O(N__60673),
            .I(N__60660));
    LocalMux I__13889 (
            .O(N__60668),
            .I(\CONTROL.addrstackptrZ0Z_2 ));
    Odrv12 I__13888 (
            .O(N__60663),
            .I(\CONTROL.addrstackptrZ0Z_2 ));
    Odrv12 I__13887 (
            .O(N__60660),
            .I(\CONTROL.addrstackptrZ0Z_2 ));
    InMux I__13886 (
            .O(N__60653),
            .I(N__60650));
    LocalMux I__13885 (
            .O(N__60650),
            .I(N__60647));
    Span4Mux_v I__13884 (
            .O(N__60647),
            .I(N__60644));
    Span4Mux_h I__13883 (
            .O(N__60644),
            .I(N__60641));
    Span4Mux_h I__13882 (
            .O(N__60641),
            .I(N__60638));
    Span4Mux_v I__13881 (
            .O(N__60638),
            .I(N__60635));
    Span4Mux_v I__13880 (
            .O(N__60635),
            .I(N__60632));
    Odrv4 I__13879 (
            .O(N__60632),
            .I(\CONTROL.g1_1_3 ));
    CascadeMux I__13878 (
            .O(N__60629),
            .I(N__60621));
    CascadeMux I__13877 (
            .O(N__60628),
            .I(N__60618));
    CascadeMux I__13876 (
            .O(N__60627),
            .I(N__60613));
    CascadeMux I__13875 (
            .O(N__60626),
            .I(N__60610));
    InMux I__13874 (
            .O(N__60625),
            .I(N__60606));
    InMux I__13873 (
            .O(N__60624),
            .I(N__60603));
    InMux I__13872 (
            .O(N__60621),
            .I(N__60599));
    InMux I__13871 (
            .O(N__60618),
            .I(N__60595));
    InMux I__13870 (
            .O(N__60617),
            .I(N__60590));
    InMux I__13869 (
            .O(N__60616),
            .I(N__60586));
    InMux I__13868 (
            .O(N__60613),
            .I(N__60580));
    InMux I__13867 (
            .O(N__60610),
            .I(N__60580));
    CascadeMux I__13866 (
            .O(N__60609),
            .I(N__60576));
    LocalMux I__13865 (
            .O(N__60606),
            .I(N__60569));
    LocalMux I__13864 (
            .O(N__60603),
            .I(N__60563));
    InMux I__13863 (
            .O(N__60602),
            .I(N__60560));
    LocalMux I__13862 (
            .O(N__60599),
            .I(N__60557));
    InMux I__13861 (
            .O(N__60598),
            .I(N__60554));
    LocalMux I__13860 (
            .O(N__60595),
            .I(N__60551));
    InMux I__13859 (
            .O(N__60594),
            .I(N__60546));
    InMux I__13858 (
            .O(N__60593),
            .I(N__60546));
    LocalMux I__13857 (
            .O(N__60590),
            .I(N__60536));
    InMux I__13856 (
            .O(N__60589),
            .I(N__60533));
    LocalMux I__13855 (
            .O(N__60586),
            .I(N__60530));
    InMux I__13854 (
            .O(N__60585),
            .I(N__60527));
    LocalMux I__13853 (
            .O(N__60580),
            .I(N__60524));
    InMux I__13852 (
            .O(N__60579),
            .I(N__60521));
    InMux I__13851 (
            .O(N__60576),
            .I(N__60518));
    InMux I__13850 (
            .O(N__60575),
            .I(N__60513));
    InMux I__13849 (
            .O(N__60574),
            .I(N__60513));
    InMux I__13848 (
            .O(N__60573),
            .I(N__60508));
    InMux I__13847 (
            .O(N__60572),
            .I(N__60508));
    Span4Mux_v I__13846 (
            .O(N__60569),
            .I(N__60505));
    InMux I__13845 (
            .O(N__60568),
            .I(N__60500));
    InMux I__13844 (
            .O(N__60567),
            .I(N__60500));
    InMux I__13843 (
            .O(N__60566),
            .I(N__60497));
    Span4Mux_v I__13842 (
            .O(N__60563),
            .I(N__60492));
    LocalMux I__13841 (
            .O(N__60560),
            .I(N__60492));
    Span4Mux_v I__13840 (
            .O(N__60557),
            .I(N__60485));
    LocalMux I__13839 (
            .O(N__60554),
            .I(N__60485));
    Span4Mux_h I__13838 (
            .O(N__60551),
            .I(N__60485));
    LocalMux I__13837 (
            .O(N__60546),
            .I(N__60482));
    InMux I__13836 (
            .O(N__60545),
            .I(N__60471));
    InMux I__13835 (
            .O(N__60544),
            .I(N__60471));
    InMux I__13834 (
            .O(N__60543),
            .I(N__60471));
    InMux I__13833 (
            .O(N__60542),
            .I(N__60471));
    InMux I__13832 (
            .O(N__60541),
            .I(N__60471));
    InMux I__13831 (
            .O(N__60540),
            .I(N__60466));
    InMux I__13830 (
            .O(N__60539),
            .I(N__60466));
    Span4Mux_h I__13829 (
            .O(N__60536),
            .I(N__60461));
    LocalMux I__13828 (
            .O(N__60533),
            .I(N__60461));
    Span4Mux_v I__13827 (
            .O(N__60530),
            .I(N__60454));
    LocalMux I__13826 (
            .O(N__60527),
            .I(N__60454));
    Span4Mux_v I__13825 (
            .O(N__60524),
            .I(N__60454));
    LocalMux I__13824 (
            .O(N__60521),
            .I(N__60451));
    LocalMux I__13823 (
            .O(N__60518),
            .I(N__60448));
    LocalMux I__13822 (
            .O(N__60513),
            .I(N__60445));
    LocalMux I__13821 (
            .O(N__60508),
            .I(N__60438));
    Span4Mux_h I__13820 (
            .O(N__60505),
            .I(N__60438));
    LocalMux I__13819 (
            .O(N__60500),
            .I(N__60438));
    LocalMux I__13818 (
            .O(N__60497),
            .I(N__60433));
    Span4Mux_v I__13817 (
            .O(N__60492),
            .I(N__60433));
    Span4Mux_v I__13816 (
            .O(N__60485),
            .I(N__60430));
    Span4Mux_v I__13815 (
            .O(N__60482),
            .I(N__60427));
    LocalMux I__13814 (
            .O(N__60471),
            .I(N__60418));
    LocalMux I__13813 (
            .O(N__60466),
            .I(N__60418));
    Span4Mux_h I__13812 (
            .O(N__60461),
            .I(N__60418));
    Span4Mux_h I__13811 (
            .O(N__60454),
            .I(N__60418));
    Span12Mux_v I__13810 (
            .O(N__60451),
            .I(N__60415));
    Span4Mux_v I__13809 (
            .O(N__60448),
            .I(N__60412));
    Span4Mux_v I__13808 (
            .O(N__60445),
            .I(N__60407));
    Span4Mux_h I__13807 (
            .O(N__60438),
            .I(N__60407));
    Span4Mux_v I__13806 (
            .O(N__60433),
            .I(N__60402));
    Span4Mux_v I__13805 (
            .O(N__60430),
            .I(N__60402));
    Span4Mux_h I__13804 (
            .O(N__60427),
            .I(N__60397));
    Span4Mux_v I__13803 (
            .O(N__60418),
            .I(N__60397));
    Odrv12 I__13802 (
            .O(N__60415),
            .I(aluOut_0));
    Odrv4 I__13801 (
            .O(N__60412),
            .I(aluOut_0));
    Odrv4 I__13800 (
            .O(N__60407),
            .I(aluOut_0));
    Odrv4 I__13799 (
            .O(N__60402),
            .I(aluOut_0));
    Odrv4 I__13798 (
            .O(N__60397),
            .I(aluOut_0));
    CascadeMux I__13797 (
            .O(N__60386),
            .I(N__60383));
    InMux I__13796 (
            .O(N__60383),
            .I(N__60380));
    LocalMux I__13795 (
            .O(N__60380),
            .I(N__60377));
    Span4Mux_h I__13794 (
            .O(N__60377),
            .I(N__60374));
    Span4Mux_h I__13793 (
            .O(N__60374),
            .I(N__60371));
    Span4Mux_v I__13792 (
            .O(N__60371),
            .I(N__60368));
    Odrv4 I__13791 (
            .O(N__60368),
            .I(\ALU.d_RNI27KBDZ0Z_0 ));
    InMux I__13790 (
            .O(N__60365),
            .I(N__60362));
    LocalMux I__13789 (
            .O(N__60362),
            .I(N__60359));
    Span12Mux_h I__13788 (
            .O(N__60359),
            .I(N__60355));
    InMux I__13787 (
            .O(N__60358),
            .I(N__60352));
    Odrv12 I__13786 (
            .O(N__60355),
            .I(\ALU.addsub_0 ));
    LocalMux I__13785 (
            .O(N__60352),
            .I(\ALU.addsub_0 ));
    InMux I__13784 (
            .O(N__60347),
            .I(\ALU.addsub_cry_0_c_THRU_CO ));
    CascadeMux I__13783 (
            .O(N__60344),
            .I(N__60341));
    InMux I__13782 (
            .O(N__60341),
            .I(N__60338));
    LocalMux I__13781 (
            .O(N__60338),
            .I(N__60335));
    Span4Mux_v I__13780 (
            .O(N__60335),
            .I(N__60332));
    Span4Mux_h I__13779 (
            .O(N__60332),
            .I(N__60329));
    Odrv4 I__13778 (
            .O(N__60329),
            .I(\ALU.d_RNIIEOKOZ0Z_1 ));
    InMux I__13777 (
            .O(N__60326),
            .I(N__60323));
    LocalMux I__13776 (
            .O(N__60323),
            .I(N__60320));
    Span12Mux_v I__13775 (
            .O(N__60320),
            .I(N__60316));
    InMux I__13774 (
            .O(N__60319),
            .I(N__60313));
    Odrv12 I__13773 (
            .O(N__60316),
            .I(\ALU.addsub_1 ));
    LocalMux I__13772 (
            .O(N__60313),
            .I(\ALU.addsub_1 ));
    InMux I__13771 (
            .O(N__60308),
            .I(\ALU.addsub_cry_0 ));
    CascadeMux I__13770 (
            .O(N__60305),
            .I(N__60302));
    InMux I__13769 (
            .O(N__60302),
            .I(N__60299));
    LocalMux I__13768 (
            .O(N__60299),
            .I(N__60296));
    Span12Mux_h I__13767 (
            .O(N__60296),
            .I(N__60293));
    Odrv12 I__13766 (
            .O(N__60293),
            .I(\ALU.d_RNIN178LZ0Z_2 ));
    InMux I__13765 (
            .O(N__60290),
            .I(N__60287));
    LocalMux I__13764 (
            .O(N__60287),
            .I(N__60284));
    Span4Mux_h I__13763 (
            .O(N__60284),
            .I(N__60281));
    Span4Mux_h I__13762 (
            .O(N__60281),
            .I(N__60277));
    InMux I__13761 (
            .O(N__60280),
            .I(N__60274));
    Odrv4 I__13760 (
            .O(N__60277),
            .I(\ALU.addsub_2 ));
    LocalMux I__13759 (
            .O(N__60274),
            .I(\ALU.addsub_2 ));
    InMux I__13758 (
            .O(N__60269),
            .I(\ALU.addsub_cry_1 ));
    InMux I__13757 (
            .O(N__60266),
            .I(N__60257));
    InMux I__13756 (
            .O(N__60265),
            .I(N__60254));
    CascadeMux I__13755 (
            .O(N__60264),
            .I(N__60251));
    CascadeMux I__13754 (
            .O(N__60263),
            .I(N__60248));
    CascadeMux I__13753 (
            .O(N__60262),
            .I(N__60242));
    InMux I__13752 (
            .O(N__60261),
            .I(N__60238));
    InMux I__13751 (
            .O(N__60260),
            .I(N__60233));
    LocalMux I__13750 (
            .O(N__60257),
            .I(N__60228));
    LocalMux I__13749 (
            .O(N__60254),
            .I(N__60228));
    InMux I__13748 (
            .O(N__60251),
            .I(N__60224));
    InMux I__13747 (
            .O(N__60248),
            .I(N__60221));
    CascadeMux I__13746 (
            .O(N__60247),
            .I(N__60215));
    InMux I__13745 (
            .O(N__60246),
            .I(N__60210));
    InMux I__13744 (
            .O(N__60245),
            .I(N__60202));
    InMux I__13743 (
            .O(N__60242),
            .I(N__60199));
    CascadeMux I__13742 (
            .O(N__60241),
            .I(N__60193));
    LocalMux I__13741 (
            .O(N__60238),
            .I(N__60184));
    InMux I__13740 (
            .O(N__60237),
            .I(N__60181));
    InMux I__13739 (
            .O(N__60236),
            .I(N__60178));
    LocalMux I__13738 (
            .O(N__60233),
            .I(N__60173));
    Span4Mux_v I__13737 (
            .O(N__60228),
            .I(N__60173));
    InMux I__13736 (
            .O(N__60227),
            .I(N__60170));
    LocalMux I__13735 (
            .O(N__60224),
            .I(N__60165));
    LocalMux I__13734 (
            .O(N__60221),
            .I(N__60165));
    InMux I__13733 (
            .O(N__60220),
            .I(N__60162));
    InMux I__13732 (
            .O(N__60219),
            .I(N__60159));
    InMux I__13731 (
            .O(N__60218),
            .I(N__60152));
    InMux I__13730 (
            .O(N__60215),
            .I(N__60152));
    InMux I__13729 (
            .O(N__60214),
            .I(N__60147));
    InMux I__13728 (
            .O(N__60213),
            .I(N__60147));
    LocalMux I__13727 (
            .O(N__60210),
            .I(N__60144));
    InMux I__13726 (
            .O(N__60209),
            .I(N__60139));
    InMux I__13725 (
            .O(N__60208),
            .I(N__60139));
    InMux I__13724 (
            .O(N__60207),
            .I(N__60134));
    InMux I__13723 (
            .O(N__60206),
            .I(N__60134));
    CascadeMux I__13722 (
            .O(N__60205),
            .I(N__60130));
    LocalMux I__13721 (
            .O(N__60202),
            .I(N__60127));
    LocalMux I__13720 (
            .O(N__60199),
            .I(N__60124));
    InMux I__13719 (
            .O(N__60198),
            .I(N__60119));
    InMux I__13718 (
            .O(N__60197),
            .I(N__60119));
    InMux I__13717 (
            .O(N__60196),
            .I(N__60109));
    InMux I__13716 (
            .O(N__60193),
            .I(N__60109));
    InMux I__13715 (
            .O(N__60192),
            .I(N__60109));
    InMux I__13714 (
            .O(N__60191),
            .I(N__60109));
    InMux I__13713 (
            .O(N__60190),
            .I(N__60102));
    InMux I__13712 (
            .O(N__60189),
            .I(N__60102));
    InMux I__13711 (
            .O(N__60188),
            .I(N__60102));
    InMux I__13710 (
            .O(N__60187),
            .I(N__60096));
    Span4Mux_v I__13709 (
            .O(N__60184),
            .I(N__60093));
    LocalMux I__13708 (
            .O(N__60181),
            .I(N__60090));
    LocalMux I__13707 (
            .O(N__60178),
            .I(N__60087));
    Span4Mux_h I__13706 (
            .O(N__60173),
            .I(N__60084));
    LocalMux I__13705 (
            .O(N__60170),
            .I(N__60079));
    Span4Mux_v I__13704 (
            .O(N__60165),
            .I(N__60079));
    LocalMux I__13703 (
            .O(N__60162),
            .I(N__60074));
    LocalMux I__13702 (
            .O(N__60159),
            .I(N__60074));
    InMux I__13701 (
            .O(N__60158),
            .I(N__60069));
    InMux I__13700 (
            .O(N__60157),
            .I(N__60069));
    LocalMux I__13699 (
            .O(N__60152),
            .I(N__60066));
    LocalMux I__13698 (
            .O(N__60147),
            .I(N__60057));
    Span4Mux_h I__13697 (
            .O(N__60144),
            .I(N__60057));
    LocalMux I__13696 (
            .O(N__60139),
            .I(N__60057));
    LocalMux I__13695 (
            .O(N__60134),
            .I(N__60057));
    InMux I__13694 (
            .O(N__60133),
            .I(N__60052));
    InMux I__13693 (
            .O(N__60130),
            .I(N__60052));
    Span4Mux_v I__13692 (
            .O(N__60127),
            .I(N__60045));
    Span4Mux_v I__13691 (
            .O(N__60124),
            .I(N__60045));
    LocalMux I__13690 (
            .O(N__60119),
            .I(N__60045));
    InMux I__13689 (
            .O(N__60118),
            .I(N__60042));
    LocalMux I__13688 (
            .O(N__60109),
            .I(N__60037));
    LocalMux I__13687 (
            .O(N__60102),
            .I(N__60037));
    InMux I__13686 (
            .O(N__60101),
            .I(N__60030));
    InMux I__13685 (
            .O(N__60100),
            .I(N__60030));
    InMux I__13684 (
            .O(N__60099),
            .I(N__60030));
    LocalMux I__13683 (
            .O(N__60096),
            .I(N__60027));
    Span4Mux_v I__13682 (
            .O(N__60093),
            .I(N__60024));
    Span4Mux_v I__13681 (
            .O(N__60090),
            .I(N__60017));
    Span4Mux_h I__13680 (
            .O(N__60087),
            .I(N__60017));
    Span4Mux_v I__13679 (
            .O(N__60084),
            .I(N__60017));
    Span4Mux_v I__13678 (
            .O(N__60079),
            .I(N__60010));
    Span4Mux_h I__13677 (
            .O(N__60074),
            .I(N__60010));
    LocalMux I__13676 (
            .O(N__60069),
            .I(N__60010));
    Span4Mux_h I__13675 (
            .O(N__60066),
            .I(N__60007));
    Span4Mux_h I__13674 (
            .O(N__60057),
            .I(N__60004));
    LocalMux I__13673 (
            .O(N__60052),
            .I(N__59999));
    Span4Mux_h I__13672 (
            .O(N__60045),
            .I(N__59999));
    LocalMux I__13671 (
            .O(N__60042),
            .I(N__59992));
    Span4Mux_v I__13670 (
            .O(N__60037),
            .I(N__59992));
    LocalMux I__13669 (
            .O(N__60030),
            .I(N__59992));
    Span12Mux_v I__13668 (
            .O(N__60027),
            .I(N__59989));
    Span4Mux_h I__13667 (
            .O(N__60024),
            .I(N__59986));
    Span4Mux_h I__13666 (
            .O(N__60017),
            .I(N__59983));
    Span4Mux_v I__13665 (
            .O(N__60010),
            .I(N__59980));
    Span4Mux_h I__13664 (
            .O(N__60007),
            .I(N__59975));
    Span4Mux_v I__13663 (
            .O(N__60004),
            .I(N__59975));
    Span4Mux_v I__13662 (
            .O(N__59999),
            .I(N__59970));
    Span4Mux_h I__13661 (
            .O(N__59992),
            .I(N__59970));
    Odrv12 I__13660 (
            .O(N__59989),
            .I(aluOut_3));
    Odrv4 I__13659 (
            .O(N__59986),
            .I(aluOut_3));
    Odrv4 I__13658 (
            .O(N__59983),
            .I(aluOut_3));
    Odrv4 I__13657 (
            .O(N__59980),
            .I(aluOut_3));
    Odrv4 I__13656 (
            .O(N__59975),
            .I(aluOut_3));
    Odrv4 I__13655 (
            .O(N__59970),
            .I(aluOut_3));
    CascadeMux I__13654 (
            .O(N__59957),
            .I(N__59954));
    InMux I__13653 (
            .O(N__59954),
            .I(N__59951));
    LocalMux I__13652 (
            .O(N__59951),
            .I(N__59948));
    Span4Mux_h I__13651 (
            .O(N__59948),
            .I(N__59945));
    Span4Mux_v I__13650 (
            .O(N__59945),
            .I(N__59942));
    Sp12to4 I__13649 (
            .O(N__59942),
            .I(N__59939));
    Odrv12 I__13648 (
            .O(N__59939),
            .I(\ALU.d_RNI04H8GZ0Z_3 ));
    InMux I__13647 (
            .O(N__59936),
            .I(N__59933));
    LocalMux I__13646 (
            .O(N__59933),
            .I(N__59930));
    Span4Mux_v I__13645 (
            .O(N__59930),
            .I(N__59926));
    InMux I__13644 (
            .O(N__59929),
            .I(N__59923));
    Span4Mux_h I__13643 (
            .O(N__59926),
            .I(N__59920));
    LocalMux I__13642 (
            .O(N__59923),
            .I(\ALU.addsub_3 ));
    Odrv4 I__13641 (
            .O(N__59920),
            .I(\ALU.addsub_3 ));
    InMux I__13640 (
            .O(N__59915),
            .I(\ALU.addsub_cry_2 ));
    CascadeMux I__13639 (
            .O(N__59912),
            .I(N__59907));
    CascadeMux I__13638 (
            .O(N__59911),
            .I(N__59904));
    InMux I__13637 (
            .O(N__59910),
            .I(N__59899));
    InMux I__13636 (
            .O(N__59907),
            .I(N__59895));
    InMux I__13635 (
            .O(N__59904),
            .I(N__59891));
    InMux I__13634 (
            .O(N__59903),
            .I(N__59888));
    CascadeMux I__13633 (
            .O(N__59902),
            .I(N__59885));
    LocalMux I__13632 (
            .O(N__59899),
            .I(N__59878));
    InMux I__13631 (
            .O(N__59898),
            .I(N__59875));
    LocalMux I__13630 (
            .O(N__59895),
            .I(N__59870));
    InMux I__13629 (
            .O(N__59894),
            .I(N__59867));
    LocalMux I__13628 (
            .O(N__59891),
            .I(N__59861));
    LocalMux I__13627 (
            .O(N__59888),
            .I(N__59858));
    InMux I__13626 (
            .O(N__59885),
            .I(N__59853));
    InMux I__13625 (
            .O(N__59884),
            .I(N__59853));
    InMux I__13624 (
            .O(N__59883),
            .I(N__59850));
    InMux I__13623 (
            .O(N__59882),
            .I(N__59846));
    InMux I__13622 (
            .O(N__59881),
            .I(N__59843));
    Span4Mux_v I__13621 (
            .O(N__59878),
            .I(N__59837));
    LocalMux I__13620 (
            .O(N__59875),
            .I(N__59834));
    InMux I__13619 (
            .O(N__59874),
            .I(N__59830));
    InMux I__13618 (
            .O(N__59873),
            .I(N__59827));
    Span4Mux_v I__13617 (
            .O(N__59870),
            .I(N__59824));
    LocalMux I__13616 (
            .O(N__59867),
            .I(N__59821));
    CascadeMux I__13615 (
            .O(N__59866),
            .I(N__59818));
    InMux I__13614 (
            .O(N__59865),
            .I(N__59814));
    InMux I__13613 (
            .O(N__59864),
            .I(N__59811));
    Span4Mux_v I__13612 (
            .O(N__59861),
            .I(N__59806));
    Span4Mux_v I__13611 (
            .O(N__59858),
            .I(N__59806));
    LocalMux I__13610 (
            .O(N__59853),
            .I(N__59803));
    LocalMux I__13609 (
            .O(N__59850),
            .I(N__59797));
    InMux I__13608 (
            .O(N__59849),
            .I(N__59794));
    LocalMux I__13607 (
            .O(N__59846),
            .I(N__59791));
    LocalMux I__13606 (
            .O(N__59843),
            .I(N__59788));
    InMux I__13605 (
            .O(N__59842),
            .I(N__59785));
    InMux I__13604 (
            .O(N__59841),
            .I(N__59780));
    InMux I__13603 (
            .O(N__59840),
            .I(N__59780));
    Span4Mux_h I__13602 (
            .O(N__59837),
            .I(N__59775));
    Span4Mux_v I__13601 (
            .O(N__59834),
            .I(N__59775));
    InMux I__13600 (
            .O(N__59833),
            .I(N__59772));
    LocalMux I__13599 (
            .O(N__59830),
            .I(N__59769));
    LocalMux I__13598 (
            .O(N__59827),
            .I(N__59766));
    Span4Mux_h I__13597 (
            .O(N__59824),
            .I(N__59761));
    Span4Mux_v I__13596 (
            .O(N__59821),
            .I(N__59761));
    InMux I__13595 (
            .O(N__59818),
            .I(N__59756));
    InMux I__13594 (
            .O(N__59817),
            .I(N__59756));
    LocalMux I__13593 (
            .O(N__59814),
            .I(N__59747));
    LocalMux I__13592 (
            .O(N__59811),
            .I(N__59747));
    Span4Mux_h I__13591 (
            .O(N__59806),
            .I(N__59747));
    Span4Mux_v I__13590 (
            .O(N__59803),
            .I(N__59747));
    InMux I__13589 (
            .O(N__59802),
            .I(N__59742));
    InMux I__13588 (
            .O(N__59801),
            .I(N__59742));
    InMux I__13587 (
            .O(N__59800),
            .I(N__59739));
    Span12Mux_v I__13586 (
            .O(N__59797),
            .I(N__59732));
    LocalMux I__13585 (
            .O(N__59794),
            .I(N__59732));
    Span12Mux_s9_h I__13584 (
            .O(N__59791),
            .I(N__59732));
    Sp12to4 I__13583 (
            .O(N__59788),
            .I(N__59725));
    LocalMux I__13582 (
            .O(N__59785),
            .I(N__59725));
    LocalMux I__13581 (
            .O(N__59780),
            .I(N__59725));
    Span4Mux_h I__13580 (
            .O(N__59775),
            .I(N__59718));
    LocalMux I__13579 (
            .O(N__59772),
            .I(N__59718));
    Span4Mux_v I__13578 (
            .O(N__59769),
            .I(N__59718));
    Span4Mux_v I__13577 (
            .O(N__59766),
            .I(N__59713));
    Span4Mux_v I__13576 (
            .O(N__59761),
            .I(N__59713));
    LocalMux I__13575 (
            .O(N__59756),
            .I(N__59708));
    Span4Mux_h I__13574 (
            .O(N__59747),
            .I(N__59708));
    LocalMux I__13573 (
            .O(N__59742),
            .I(aluOut_4));
    LocalMux I__13572 (
            .O(N__59739),
            .I(aluOut_4));
    Odrv12 I__13571 (
            .O(N__59732),
            .I(aluOut_4));
    Odrv12 I__13570 (
            .O(N__59725),
            .I(aluOut_4));
    Odrv4 I__13569 (
            .O(N__59718),
            .I(aluOut_4));
    Odrv4 I__13568 (
            .O(N__59713),
            .I(aluOut_4));
    Odrv4 I__13567 (
            .O(N__59708),
            .I(aluOut_4));
    CascadeMux I__13566 (
            .O(N__59693),
            .I(N__59690));
    InMux I__13565 (
            .O(N__59690),
            .I(N__59687));
    LocalMux I__13564 (
            .O(N__59687),
            .I(N__59684));
    Span4Mux_v I__13563 (
            .O(N__59684),
            .I(N__59681));
    Sp12to4 I__13562 (
            .O(N__59681),
            .I(N__59678));
    Span12Mux_h I__13561 (
            .O(N__59678),
            .I(N__59675));
    Odrv12 I__13560 (
            .O(N__59675),
            .I(\ALU.d_RNI7BF7IZ0Z_4 ));
    InMux I__13559 (
            .O(N__59672),
            .I(N__59669));
    LocalMux I__13558 (
            .O(N__59669),
            .I(N__59666));
    Span12Mux_v I__13557 (
            .O(N__59666),
            .I(N__59662));
    InMux I__13556 (
            .O(N__59665),
            .I(N__59659));
    Span12Mux_h I__13555 (
            .O(N__59662),
            .I(N__59656));
    LocalMux I__13554 (
            .O(N__59659),
            .I(N__59653));
    Odrv12 I__13553 (
            .O(N__59656),
            .I(\ALU.addsub_4 ));
    Odrv4 I__13552 (
            .O(N__59653),
            .I(\ALU.addsub_4 ));
    InMux I__13551 (
            .O(N__59648),
            .I(\ALU.addsub_cry_3 ));
    CascadeMux I__13550 (
            .O(N__59645),
            .I(N__59641));
    InMux I__13549 (
            .O(N__59644),
            .I(N__59634));
    InMux I__13548 (
            .O(N__59641),
            .I(N__59629));
    InMux I__13547 (
            .O(N__59640),
            .I(N__59629));
    InMux I__13546 (
            .O(N__59639),
            .I(N__59626));
    InMux I__13545 (
            .O(N__59638),
            .I(N__59621));
    InMux I__13544 (
            .O(N__59637),
            .I(N__59615));
    LocalMux I__13543 (
            .O(N__59634),
            .I(N__59612));
    LocalMux I__13542 (
            .O(N__59629),
            .I(N__59609));
    LocalMux I__13541 (
            .O(N__59626),
            .I(N__59606));
    InMux I__13540 (
            .O(N__59625),
            .I(N__59603));
    CascadeMux I__13539 (
            .O(N__59624),
            .I(N__59596));
    LocalMux I__13538 (
            .O(N__59621),
            .I(N__59592));
    InMux I__13537 (
            .O(N__59620),
            .I(N__59589));
    InMux I__13536 (
            .O(N__59619),
            .I(N__59577));
    InMux I__13535 (
            .O(N__59618),
            .I(N__59577));
    LocalMux I__13534 (
            .O(N__59615),
            .I(N__59574));
    Span4Mux_v I__13533 (
            .O(N__59612),
            .I(N__59567));
    Span4Mux_v I__13532 (
            .O(N__59609),
            .I(N__59567));
    Span4Mux_v I__13531 (
            .O(N__59606),
            .I(N__59567));
    LocalMux I__13530 (
            .O(N__59603),
            .I(N__59564));
    InMux I__13529 (
            .O(N__59602),
            .I(N__59557));
    InMux I__13528 (
            .O(N__59601),
            .I(N__59557));
    InMux I__13527 (
            .O(N__59600),
            .I(N__59557));
    CascadeMux I__13526 (
            .O(N__59599),
            .I(N__59554));
    InMux I__13525 (
            .O(N__59596),
            .I(N__59551));
    InMux I__13524 (
            .O(N__59595),
            .I(N__59546));
    Span4Mux_h I__13523 (
            .O(N__59592),
            .I(N__59541));
    LocalMux I__13522 (
            .O(N__59589),
            .I(N__59541));
    InMux I__13521 (
            .O(N__59588),
            .I(N__59537));
    InMux I__13520 (
            .O(N__59587),
            .I(N__59534));
    InMux I__13519 (
            .O(N__59586),
            .I(N__59531));
    InMux I__13518 (
            .O(N__59585),
            .I(N__59528));
    InMux I__13517 (
            .O(N__59584),
            .I(N__59521));
    InMux I__13516 (
            .O(N__59583),
            .I(N__59521));
    InMux I__13515 (
            .O(N__59582),
            .I(N__59521));
    LocalMux I__13514 (
            .O(N__59577),
            .I(N__59518));
    Span4Mux_v I__13513 (
            .O(N__59574),
            .I(N__59515));
    Span4Mux_h I__13512 (
            .O(N__59567),
            .I(N__59512));
    Span4Mux_h I__13511 (
            .O(N__59564),
            .I(N__59507));
    LocalMux I__13510 (
            .O(N__59557),
            .I(N__59507));
    InMux I__13509 (
            .O(N__59554),
            .I(N__59504));
    LocalMux I__13508 (
            .O(N__59551),
            .I(N__59500));
    InMux I__13507 (
            .O(N__59550),
            .I(N__59497));
    InMux I__13506 (
            .O(N__59549),
            .I(N__59494));
    LocalMux I__13505 (
            .O(N__59546),
            .I(N__59491));
    Span4Mux_h I__13504 (
            .O(N__59541),
            .I(N__59488));
    CascadeMux I__13503 (
            .O(N__59540),
            .I(N__59480));
    LocalMux I__13502 (
            .O(N__59537),
            .I(N__59473));
    LocalMux I__13501 (
            .O(N__59534),
            .I(N__59470));
    LocalMux I__13500 (
            .O(N__59531),
            .I(N__59463));
    LocalMux I__13499 (
            .O(N__59528),
            .I(N__59463));
    LocalMux I__13498 (
            .O(N__59521),
            .I(N__59463));
    Span4Mux_v I__13497 (
            .O(N__59518),
            .I(N__59454));
    Span4Mux_h I__13496 (
            .O(N__59515),
            .I(N__59454));
    Span4Mux_h I__13495 (
            .O(N__59512),
            .I(N__59454));
    Span4Mux_v I__13494 (
            .O(N__59507),
            .I(N__59454));
    LocalMux I__13493 (
            .O(N__59504),
            .I(N__59451));
    InMux I__13492 (
            .O(N__59503),
            .I(N__59448));
    Span4Mux_h I__13491 (
            .O(N__59500),
            .I(N__59439));
    LocalMux I__13490 (
            .O(N__59497),
            .I(N__59439));
    LocalMux I__13489 (
            .O(N__59494),
            .I(N__59439));
    Span4Mux_v I__13488 (
            .O(N__59491),
            .I(N__59439));
    Span4Mux_h I__13487 (
            .O(N__59488),
            .I(N__59436));
    InMux I__13486 (
            .O(N__59487),
            .I(N__59431));
    InMux I__13485 (
            .O(N__59486),
            .I(N__59431));
    InMux I__13484 (
            .O(N__59485),
            .I(N__59424));
    InMux I__13483 (
            .O(N__59484),
            .I(N__59424));
    InMux I__13482 (
            .O(N__59483),
            .I(N__59424));
    InMux I__13481 (
            .O(N__59480),
            .I(N__59413));
    InMux I__13480 (
            .O(N__59479),
            .I(N__59413));
    InMux I__13479 (
            .O(N__59478),
            .I(N__59413));
    InMux I__13478 (
            .O(N__59477),
            .I(N__59413));
    InMux I__13477 (
            .O(N__59476),
            .I(N__59413));
    Span4Mux_h I__13476 (
            .O(N__59473),
            .I(N__59406));
    Span4Mux_v I__13475 (
            .O(N__59470),
            .I(N__59406));
    Span4Mux_h I__13474 (
            .O(N__59463),
            .I(N__59406));
    Span4Mux_h I__13473 (
            .O(N__59454),
            .I(N__59403));
    Odrv12 I__13472 (
            .O(N__59451),
            .I(aluOut_5));
    LocalMux I__13471 (
            .O(N__59448),
            .I(aluOut_5));
    Odrv4 I__13470 (
            .O(N__59439),
            .I(aluOut_5));
    Odrv4 I__13469 (
            .O(N__59436),
            .I(aluOut_5));
    LocalMux I__13468 (
            .O(N__59431),
            .I(aluOut_5));
    LocalMux I__13467 (
            .O(N__59424),
            .I(aluOut_5));
    LocalMux I__13466 (
            .O(N__59413),
            .I(aluOut_5));
    Odrv4 I__13465 (
            .O(N__59406),
            .I(aluOut_5));
    Odrv4 I__13464 (
            .O(N__59403),
            .I(aluOut_5));
    CascadeMux I__13463 (
            .O(N__59384),
            .I(N__59381));
    InMux I__13462 (
            .O(N__59381),
            .I(N__59378));
    LocalMux I__13461 (
            .O(N__59378),
            .I(N__59375));
    Span12Mux_s10_h I__13460 (
            .O(N__59375),
            .I(N__59372));
    Odrv12 I__13459 (
            .O(N__59372),
            .I(\ALU.d_RNI58QFIZ0Z_5 ));
    InMux I__13458 (
            .O(N__59369),
            .I(N__59366));
    LocalMux I__13457 (
            .O(N__59366),
            .I(N__59363));
    Span4Mux_h I__13456 (
            .O(N__59363),
            .I(N__59360));
    Span4Mux_h I__13455 (
            .O(N__59360),
            .I(N__59357));
    Span4Mux_h I__13454 (
            .O(N__59357),
            .I(N__59354));
    Span4Mux_v I__13453 (
            .O(N__59354),
            .I(N__59350));
    InMux I__13452 (
            .O(N__59353),
            .I(N__59347));
    Odrv4 I__13451 (
            .O(N__59350),
            .I(\ALU.addsub_5 ));
    LocalMux I__13450 (
            .O(N__59347),
            .I(\ALU.addsub_5 ));
    InMux I__13449 (
            .O(N__59342),
            .I(\ALU.addsub_cry_4 ));
    InMux I__13448 (
            .O(N__59339),
            .I(N__59335));
    InMux I__13447 (
            .O(N__59338),
            .I(N__59332));
    LocalMux I__13446 (
            .O(N__59335),
            .I(N__59329));
    LocalMux I__13445 (
            .O(N__59332),
            .I(N__59325));
    Span4Mux_v I__13444 (
            .O(N__59329),
            .I(N__59322));
    InMux I__13443 (
            .O(N__59328),
            .I(N__59319));
    Span4Mux_h I__13442 (
            .O(N__59325),
            .I(N__59316));
    Span4Mux_h I__13441 (
            .O(N__59322),
            .I(N__59313));
    LocalMux I__13440 (
            .O(N__59319),
            .I(\ALU.a_15_m2_sZ0Z_15 ));
    Odrv4 I__13439 (
            .O(N__59316),
            .I(\ALU.a_15_m2_sZ0Z_15 ));
    Odrv4 I__13438 (
            .O(N__59313),
            .I(\ALU.a_15_m2_sZ0Z_15 ));
    InMux I__13437 (
            .O(N__59306),
            .I(N__59302));
    InMux I__13436 (
            .O(N__59305),
            .I(N__59299));
    LocalMux I__13435 (
            .O(N__59302),
            .I(N__59292));
    LocalMux I__13434 (
            .O(N__59299),
            .I(N__59283));
    InMux I__13433 (
            .O(N__59298),
            .I(N__59276));
    InMux I__13432 (
            .O(N__59297),
            .I(N__59276));
    InMux I__13431 (
            .O(N__59296),
            .I(N__59271));
    InMux I__13430 (
            .O(N__59295),
            .I(N__59271));
    Span4Mux_v I__13429 (
            .O(N__59292),
            .I(N__59268));
    InMux I__13428 (
            .O(N__59291),
            .I(N__59263));
    InMux I__13427 (
            .O(N__59290),
            .I(N__59259));
    InMux I__13426 (
            .O(N__59289),
            .I(N__59250));
    InMux I__13425 (
            .O(N__59288),
            .I(N__59250));
    InMux I__13424 (
            .O(N__59287),
            .I(N__59250));
    InMux I__13423 (
            .O(N__59286),
            .I(N__59250));
    Span4Mux_v I__13422 (
            .O(N__59283),
            .I(N__59245));
    InMux I__13421 (
            .O(N__59282),
            .I(N__59240));
    InMux I__13420 (
            .O(N__59281),
            .I(N__59240));
    LocalMux I__13419 (
            .O(N__59276),
            .I(N__59235));
    LocalMux I__13418 (
            .O(N__59271),
            .I(N__59235));
    Span4Mux_h I__13417 (
            .O(N__59268),
            .I(N__59232));
    InMux I__13416 (
            .O(N__59267),
            .I(N__59229));
    InMux I__13415 (
            .O(N__59266),
            .I(N__59226));
    LocalMux I__13414 (
            .O(N__59263),
            .I(N__59223));
    InMux I__13413 (
            .O(N__59262),
            .I(N__59220));
    LocalMux I__13412 (
            .O(N__59259),
            .I(N__59215));
    LocalMux I__13411 (
            .O(N__59250),
            .I(N__59215));
    InMux I__13410 (
            .O(N__59249),
            .I(N__59212));
    InMux I__13409 (
            .O(N__59248),
            .I(N__59209));
    Sp12to4 I__13408 (
            .O(N__59245),
            .I(N__59202));
    LocalMux I__13407 (
            .O(N__59240),
            .I(N__59202));
    Span12Mux_v I__13406 (
            .O(N__59235),
            .I(N__59202));
    Span4Mux_v I__13405 (
            .O(N__59232),
            .I(N__59195));
    LocalMux I__13404 (
            .O(N__59229),
            .I(N__59195));
    LocalMux I__13403 (
            .O(N__59226),
            .I(N__59195));
    Span4Mux_h I__13402 (
            .O(N__59223),
            .I(N__59188));
    LocalMux I__13401 (
            .O(N__59220),
            .I(N__59188));
    Span4Mux_h I__13400 (
            .O(N__59215),
            .I(N__59188));
    LocalMux I__13399 (
            .O(N__59212),
            .I(\ALU.a_15_sm0 ));
    LocalMux I__13398 (
            .O(N__59209),
            .I(\ALU.a_15_sm0 ));
    Odrv12 I__13397 (
            .O(N__59202),
            .I(\ALU.a_15_sm0 ));
    Odrv4 I__13396 (
            .O(N__59195),
            .I(\ALU.a_15_sm0 ));
    Odrv4 I__13395 (
            .O(N__59188),
            .I(\ALU.a_15_sm0 ));
    CascadeMux I__13394 (
            .O(N__59177),
            .I(N__59173));
    CascadeMux I__13393 (
            .O(N__59176),
            .I(N__59170));
    InMux I__13392 (
            .O(N__59173),
            .I(N__59166));
    InMux I__13391 (
            .O(N__59170),
            .I(N__59163));
    InMux I__13390 (
            .O(N__59169),
            .I(N__59160));
    LocalMux I__13389 (
            .O(N__59166),
            .I(N__59151));
    LocalMux I__13388 (
            .O(N__59163),
            .I(N__59151));
    LocalMux I__13387 (
            .O(N__59160),
            .I(N__59151));
    InMux I__13386 (
            .O(N__59159),
            .I(N__59146));
    InMux I__13385 (
            .O(N__59158),
            .I(N__59146));
    Span4Mux_v I__13384 (
            .O(N__59151),
            .I(N__59133));
    LocalMux I__13383 (
            .O(N__59146),
            .I(N__59130));
    InMux I__13382 (
            .O(N__59145),
            .I(N__59125));
    InMux I__13381 (
            .O(N__59144),
            .I(N__59125));
    CascadeMux I__13380 (
            .O(N__59143),
            .I(N__59121));
    CascadeMux I__13379 (
            .O(N__59142),
            .I(N__59117));
    CascadeMux I__13378 (
            .O(N__59141),
            .I(N__59114));
    CascadeMux I__13377 (
            .O(N__59140),
            .I(N__59111));
    CascadeMux I__13376 (
            .O(N__59139),
            .I(N__59108));
    CascadeMux I__13375 (
            .O(N__59138),
            .I(N__59103));
    InMux I__13374 (
            .O(N__59137),
            .I(N__59095));
    InMux I__13373 (
            .O(N__59136),
            .I(N__59095));
    Span4Mux_v I__13372 (
            .O(N__59133),
            .I(N__59088));
    Span4Mux_h I__13371 (
            .O(N__59130),
            .I(N__59088));
    LocalMux I__13370 (
            .O(N__59125),
            .I(N__59088));
    InMux I__13369 (
            .O(N__59124),
            .I(N__59085));
    InMux I__13368 (
            .O(N__59121),
            .I(N__59082));
    CascadeMux I__13367 (
            .O(N__59120),
            .I(N__59079));
    InMux I__13366 (
            .O(N__59117),
            .I(N__59076));
    InMux I__13365 (
            .O(N__59114),
            .I(N__59073));
    InMux I__13364 (
            .O(N__59111),
            .I(N__59070));
    InMux I__13363 (
            .O(N__59108),
            .I(N__59067));
    InMux I__13362 (
            .O(N__59107),
            .I(N__59059));
    InMux I__13361 (
            .O(N__59106),
            .I(N__59059));
    InMux I__13360 (
            .O(N__59103),
            .I(N__59059));
    InMux I__13359 (
            .O(N__59102),
            .I(N__59056));
    InMux I__13358 (
            .O(N__59101),
            .I(N__59051));
    InMux I__13357 (
            .O(N__59100),
            .I(N__59051));
    LocalMux I__13356 (
            .O(N__59095),
            .I(N__59045));
    Span4Mux_h I__13355 (
            .O(N__59088),
            .I(N__59037));
    LocalMux I__13354 (
            .O(N__59085),
            .I(N__59037));
    LocalMux I__13353 (
            .O(N__59082),
            .I(N__59034));
    InMux I__13352 (
            .O(N__59079),
            .I(N__59031));
    LocalMux I__13351 (
            .O(N__59076),
            .I(N__59024));
    LocalMux I__13350 (
            .O(N__59073),
            .I(N__59024));
    LocalMux I__13349 (
            .O(N__59070),
            .I(N__59024));
    LocalMux I__13348 (
            .O(N__59067),
            .I(N__59021));
    InMux I__13347 (
            .O(N__59066),
            .I(N__59018));
    LocalMux I__13346 (
            .O(N__59059),
            .I(N__59013));
    LocalMux I__13345 (
            .O(N__59056),
            .I(N__59013));
    LocalMux I__13344 (
            .O(N__59051),
            .I(N__59010));
    CascadeMux I__13343 (
            .O(N__59050),
            .I(N__59006));
    CascadeMux I__13342 (
            .O(N__59049),
            .I(N__59002));
    CascadeMux I__13341 (
            .O(N__59048),
            .I(N__58998));
    Span4Mux_v I__13340 (
            .O(N__59045),
            .I(N__58995));
    InMux I__13339 (
            .O(N__59044),
            .I(N__58988));
    InMux I__13338 (
            .O(N__59043),
            .I(N__58988));
    InMux I__13337 (
            .O(N__59042),
            .I(N__58988));
    Span4Mux_v I__13336 (
            .O(N__59037),
            .I(N__58984));
    Span4Mux_v I__13335 (
            .O(N__59034),
            .I(N__58981));
    LocalMux I__13334 (
            .O(N__59031),
            .I(N__58976));
    Span4Mux_v I__13333 (
            .O(N__59024),
            .I(N__58976));
    Span4Mux_v I__13332 (
            .O(N__59021),
            .I(N__58971));
    LocalMux I__13331 (
            .O(N__59018),
            .I(N__58971));
    Span4Mux_v I__13330 (
            .O(N__59013),
            .I(N__58968));
    Span4Mux_h I__13329 (
            .O(N__59010),
            .I(N__58965));
    InMux I__13328 (
            .O(N__59009),
            .I(N__58958));
    InMux I__13327 (
            .O(N__59006),
            .I(N__58958));
    InMux I__13326 (
            .O(N__59005),
            .I(N__58958));
    InMux I__13325 (
            .O(N__59002),
            .I(N__58951));
    InMux I__13324 (
            .O(N__59001),
            .I(N__58951));
    InMux I__13323 (
            .O(N__58998),
            .I(N__58951));
    Span4Mux_h I__13322 (
            .O(N__58995),
            .I(N__58946));
    LocalMux I__13321 (
            .O(N__58988),
            .I(N__58946));
    InMux I__13320 (
            .O(N__58987),
            .I(N__58943));
    Sp12to4 I__13319 (
            .O(N__58984),
            .I(N__58940));
    Span4Mux_h I__13318 (
            .O(N__58981),
            .I(N__58933));
    Span4Mux_v I__13317 (
            .O(N__58976),
            .I(N__58933));
    Span4Mux_v I__13316 (
            .O(N__58971),
            .I(N__58933));
    Span4Mux_v I__13315 (
            .O(N__58968),
            .I(N__58930));
    Span4Mux_v I__13314 (
            .O(N__58965),
            .I(N__58927));
    LocalMux I__13313 (
            .O(N__58958),
            .I(N__58920));
    LocalMux I__13312 (
            .O(N__58951),
            .I(N__58920));
    Span4Mux_h I__13311 (
            .O(N__58946),
            .I(N__58920));
    LocalMux I__13310 (
            .O(N__58943),
            .I(N__58915));
    Span12Mux_h I__13309 (
            .O(N__58940),
            .I(N__58915));
    Sp12to4 I__13308 (
            .O(N__58933),
            .I(N__58910));
    Sp12to4 I__13307 (
            .O(N__58930),
            .I(N__58910));
    Span4Mux_v I__13306 (
            .O(N__58927),
            .I(N__58907));
    Span4Mux_v I__13305 (
            .O(N__58920),
            .I(N__58904));
    Span12Mux_v I__13304 (
            .O(N__58915),
            .I(N__58899));
    Span12Mux_h I__13303 (
            .O(N__58910),
            .I(N__58899));
    Span4Mux_h I__13302 (
            .O(N__58907),
            .I(N__58894));
    Span4Mux_v I__13301 (
            .O(N__58904),
            .I(N__58894));
    Odrv12 I__13300 (
            .O(N__58899),
            .I(aluOperation_1));
    Odrv4 I__13299 (
            .O(N__58894),
            .I(aluOperation_1));
    InMux I__13298 (
            .O(N__58889),
            .I(N__58881));
    InMux I__13297 (
            .O(N__58888),
            .I(N__58878));
    InMux I__13296 (
            .O(N__58887),
            .I(N__58874));
    InMux I__13295 (
            .O(N__58886),
            .I(N__58871));
    InMux I__13294 (
            .O(N__58885),
            .I(N__58868));
    InMux I__13293 (
            .O(N__58884),
            .I(N__58865));
    LocalMux I__13292 (
            .O(N__58881),
            .I(N__58861));
    LocalMux I__13291 (
            .O(N__58878),
            .I(N__58858));
    InMux I__13290 (
            .O(N__58877),
            .I(N__58855));
    LocalMux I__13289 (
            .O(N__58874),
            .I(N__58850));
    LocalMux I__13288 (
            .O(N__58871),
            .I(N__58850));
    LocalMux I__13287 (
            .O(N__58868),
            .I(N__58845));
    LocalMux I__13286 (
            .O(N__58865),
            .I(N__58845));
    InMux I__13285 (
            .O(N__58864),
            .I(N__58842));
    Span4Mux_h I__13284 (
            .O(N__58861),
            .I(N__58839));
    Span4Mux_h I__13283 (
            .O(N__58858),
            .I(N__58836));
    LocalMux I__13282 (
            .O(N__58855),
            .I(N__58831));
    Span4Mux_v I__13281 (
            .O(N__58850),
            .I(N__58831));
    Span4Mux_v I__13280 (
            .O(N__58845),
            .I(N__58828));
    LocalMux I__13279 (
            .O(N__58842),
            .I(\ALU.a_15_ns_1_7 ));
    Odrv4 I__13278 (
            .O(N__58839),
            .I(\ALU.a_15_ns_1_7 ));
    Odrv4 I__13277 (
            .O(N__58836),
            .I(\ALU.a_15_ns_1_7 ));
    Odrv4 I__13276 (
            .O(N__58831),
            .I(\ALU.a_15_ns_1_7 ));
    Odrv4 I__13275 (
            .O(N__58828),
            .I(\ALU.a_15_ns_1_7 ));
    InMux I__13274 (
            .O(N__58817),
            .I(N__58813));
    InMux I__13273 (
            .O(N__58816),
            .I(N__58809));
    LocalMux I__13272 (
            .O(N__58813),
            .I(N__58805));
    InMux I__13271 (
            .O(N__58812),
            .I(N__58802));
    LocalMux I__13270 (
            .O(N__58809),
            .I(N__58796));
    InMux I__13269 (
            .O(N__58808),
            .I(N__58793));
    Span4Mux_h I__13268 (
            .O(N__58805),
            .I(N__58790));
    LocalMux I__13267 (
            .O(N__58802),
            .I(N__58787));
    InMux I__13266 (
            .O(N__58801),
            .I(N__58784));
    InMux I__13265 (
            .O(N__58800),
            .I(N__58781));
    InMux I__13264 (
            .O(N__58799),
            .I(N__58778));
    Span4Mux_v I__13263 (
            .O(N__58796),
            .I(N__58773));
    LocalMux I__13262 (
            .O(N__58793),
            .I(N__58773));
    Span4Mux_h I__13261 (
            .O(N__58790),
            .I(N__58768));
    Span4Mux_v I__13260 (
            .O(N__58787),
            .I(N__58768));
    LocalMux I__13259 (
            .O(N__58784),
            .I(\ALU.mult_388_c_RNIPGN6QZ0Z7 ));
    LocalMux I__13258 (
            .O(N__58781),
            .I(\ALU.mult_388_c_RNIPGN6QZ0Z7 ));
    LocalMux I__13257 (
            .O(N__58778),
            .I(\ALU.mult_388_c_RNIPGN6QZ0Z7 ));
    Odrv4 I__13256 (
            .O(N__58773),
            .I(\ALU.mult_388_c_RNIPGN6QZ0Z7 ));
    Odrv4 I__13255 (
            .O(N__58768),
            .I(\ALU.mult_388_c_RNIPGN6QZ0Z7 ));
    InMux I__13254 (
            .O(N__58757),
            .I(N__58753));
    CascadeMux I__13253 (
            .O(N__58756),
            .I(N__58749));
    LocalMux I__13252 (
            .O(N__58753),
            .I(N__58746));
    InMux I__13251 (
            .O(N__58752),
            .I(N__58742));
    InMux I__13250 (
            .O(N__58749),
            .I(N__58736));
    Span4Mux_v I__13249 (
            .O(N__58746),
            .I(N__58733));
    InMux I__13248 (
            .O(N__58745),
            .I(N__58730));
    LocalMux I__13247 (
            .O(N__58742),
            .I(N__58727));
    InMux I__13246 (
            .O(N__58741),
            .I(N__58724));
    InMux I__13245 (
            .O(N__58740),
            .I(N__58721));
    InMux I__13244 (
            .O(N__58739),
            .I(N__58718));
    LocalMux I__13243 (
            .O(N__58736),
            .I(N__58714));
    Span4Mux_h I__13242 (
            .O(N__58733),
            .I(N__58709));
    LocalMux I__13241 (
            .O(N__58730),
            .I(N__58709));
    Span4Mux_v I__13240 (
            .O(N__58727),
            .I(N__58706));
    LocalMux I__13239 (
            .O(N__58724),
            .I(N__58699));
    LocalMux I__13238 (
            .O(N__58721),
            .I(N__58699));
    LocalMux I__13237 (
            .O(N__58718),
            .I(N__58699));
    InMux I__13236 (
            .O(N__58717),
            .I(N__58696));
    Span4Mux_v I__13235 (
            .O(N__58714),
            .I(N__58691));
    Span4Mux_v I__13234 (
            .O(N__58709),
            .I(N__58691));
    Span4Mux_h I__13233 (
            .O(N__58706),
            .I(N__58684));
    Span4Mux_v I__13232 (
            .O(N__58699),
            .I(N__58684));
    LocalMux I__13231 (
            .O(N__58696),
            .I(N__58684));
    Odrv4 I__13230 (
            .O(N__58691),
            .I(\ALU.rshift_3 ));
    Odrv4 I__13229 (
            .O(N__58684),
            .I(\ALU.rshift_3 ));
    InMux I__13228 (
            .O(N__58679),
            .I(N__58673));
    InMux I__13227 (
            .O(N__58678),
            .I(N__58670));
    InMux I__13226 (
            .O(N__58677),
            .I(N__58667));
    InMux I__13225 (
            .O(N__58676),
            .I(N__58660));
    LocalMux I__13224 (
            .O(N__58673),
            .I(N__58657));
    LocalMux I__13223 (
            .O(N__58670),
            .I(N__58654));
    LocalMux I__13222 (
            .O(N__58667),
            .I(N__58651));
    InMux I__13221 (
            .O(N__58666),
            .I(N__58648));
    InMux I__13220 (
            .O(N__58665),
            .I(N__58645));
    InMux I__13219 (
            .O(N__58664),
            .I(N__58642));
    InMux I__13218 (
            .O(N__58663),
            .I(N__58639));
    LocalMux I__13217 (
            .O(N__58660),
            .I(N__58636));
    Span4Mux_v I__13216 (
            .O(N__58657),
            .I(N__58633));
    Span4Mux_h I__13215 (
            .O(N__58654),
            .I(N__58630));
    Span12Mux_h I__13214 (
            .O(N__58651),
            .I(N__58627));
    LocalMux I__13213 (
            .O(N__58648),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    LocalMux I__13212 (
            .O(N__58645),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    LocalMux I__13211 (
            .O(N__58642),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    LocalMux I__13210 (
            .O(N__58639),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    Odrv4 I__13209 (
            .O(N__58636),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    Odrv4 I__13208 (
            .O(N__58633),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    Odrv4 I__13207 (
            .O(N__58630),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    Odrv12 I__13206 (
            .O(N__58627),
            .I(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ));
    InMux I__13205 (
            .O(N__58610),
            .I(N__58607));
    LocalMux I__13204 (
            .O(N__58607),
            .I(N__58603));
    InMux I__13203 (
            .O(N__58606),
            .I(N__58599));
    Span4Mux_v I__13202 (
            .O(N__58603),
            .I(N__58596));
    InMux I__13201 (
            .O(N__58602),
            .I(N__58593));
    LocalMux I__13200 (
            .O(N__58599),
            .I(N__58590));
    Span4Mux_h I__13199 (
            .O(N__58596),
            .I(N__58585));
    LocalMux I__13198 (
            .O(N__58593),
            .I(N__58585));
    Span4Mux_h I__13197 (
            .O(N__58590),
            .I(N__58582));
    Span4Mux_h I__13196 (
            .O(N__58585),
            .I(N__58579));
    Span4Mux_h I__13195 (
            .O(N__58582),
            .I(N__58576));
    Span4Mux_v I__13194 (
            .O(N__58579),
            .I(N__58573));
    Span4Mux_v I__13193 (
            .O(N__58576),
            .I(N__58570));
    Odrv4 I__13192 (
            .O(N__58573),
            .I(h_3));
    Odrv4 I__13191 (
            .O(N__58570),
            .I(h_3));
    CascadeMux I__13190 (
            .O(N__58565),
            .I(N__58559));
    CascadeMux I__13189 (
            .O(N__58564),
            .I(N__58556));
    CascadeMux I__13188 (
            .O(N__58563),
            .I(N__58553));
    InMux I__13187 (
            .O(N__58562),
            .I(N__58548));
    InMux I__13186 (
            .O(N__58559),
            .I(N__58544));
    InMux I__13185 (
            .O(N__58556),
            .I(N__58541));
    InMux I__13184 (
            .O(N__58553),
            .I(N__58538));
    InMux I__13183 (
            .O(N__58552),
            .I(N__58535));
    CascadeMux I__13182 (
            .O(N__58551),
            .I(N__58530));
    LocalMux I__13181 (
            .O(N__58548),
            .I(N__58527));
    CascadeMux I__13180 (
            .O(N__58547),
            .I(N__58521));
    LocalMux I__13179 (
            .O(N__58544),
            .I(N__58516));
    LocalMux I__13178 (
            .O(N__58541),
            .I(N__58516));
    LocalMux I__13177 (
            .O(N__58538),
            .I(N__58511));
    LocalMux I__13176 (
            .O(N__58535),
            .I(N__58511));
    InMux I__13175 (
            .O(N__58534),
            .I(N__58505));
    InMux I__13174 (
            .O(N__58533),
            .I(N__58505));
    InMux I__13173 (
            .O(N__58530),
            .I(N__58502));
    Span4Mux_v I__13172 (
            .O(N__58527),
            .I(N__58499));
    InMux I__13171 (
            .O(N__58526),
            .I(N__58491));
    InMux I__13170 (
            .O(N__58525),
            .I(N__58488));
    InMux I__13169 (
            .O(N__58524),
            .I(N__58485));
    InMux I__13168 (
            .O(N__58521),
            .I(N__58482));
    Span4Mux_v I__13167 (
            .O(N__58516),
            .I(N__58479));
    Span4Mux_h I__13166 (
            .O(N__58511),
            .I(N__58476));
    InMux I__13165 (
            .O(N__58510),
            .I(N__58473));
    LocalMux I__13164 (
            .O(N__58505),
            .I(N__58470));
    LocalMux I__13163 (
            .O(N__58502),
            .I(N__58465));
    Sp12to4 I__13162 (
            .O(N__58499),
            .I(N__58465));
    InMux I__13161 (
            .O(N__58498),
            .I(N__58462));
    InMux I__13160 (
            .O(N__58497),
            .I(N__58457));
    InMux I__13159 (
            .O(N__58496),
            .I(N__58457));
    InMux I__13158 (
            .O(N__58495),
            .I(N__58452));
    InMux I__13157 (
            .O(N__58494),
            .I(N__58449));
    LocalMux I__13156 (
            .O(N__58491),
            .I(N__58444));
    LocalMux I__13155 (
            .O(N__58488),
            .I(N__58444));
    LocalMux I__13154 (
            .O(N__58485),
            .I(N__58439));
    LocalMux I__13153 (
            .O(N__58482),
            .I(N__58439));
    Span4Mux_h I__13152 (
            .O(N__58479),
            .I(N__58434));
    Span4Mux_v I__13151 (
            .O(N__58476),
            .I(N__58434));
    LocalMux I__13150 (
            .O(N__58473),
            .I(N__58431));
    Span4Mux_v I__13149 (
            .O(N__58470),
            .I(N__58428));
    Span12Mux_h I__13148 (
            .O(N__58465),
            .I(N__58423));
    LocalMux I__13147 (
            .O(N__58462),
            .I(N__58423));
    LocalMux I__13146 (
            .O(N__58457),
            .I(N__58420));
    InMux I__13145 (
            .O(N__58456),
            .I(N__58417));
    InMux I__13144 (
            .O(N__58455),
            .I(N__58414));
    LocalMux I__13143 (
            .O(N__58452),
            .I(N__58409));
    LocalMux I__13142 (
            .O(N__58449),
            .I(N__58409));
    Span12Mux_v I__13141 (
            .O(N__58444),
            .I(N__58406));
    Span12Mux_v I__13140 (
            .O(N__58439),
            .I(N__58403));
    Span4Mux_v I__13139 (
            .O(N__58434),
            .I(N__58396));
    Span4Mux_v I__13138 (
            .O(N__58431),
            .I(N__58396));
    Span4Mux_h I__13137 (
            .O(N__58428),
            .I(N__58396));
    Span12Mux_v I__13136 (
            .O(N__58423),
            .I(N__58393));
    Span4Mux_h I__13135 (
            .O(N__58420),
            .I(N__58390));
    LocalMux I__13134 (
            .O(N__58417),
            .I(\ALU.a_15_sZ0Z_13 ));
    LocalMux I__13133 (
            .O(N__58414),
            .I(\ALU.a_15_sZ0Z_13 ));
    Odrv4 I__13132 (
            .O(N__58409),
            .I(\ALU.a_15_sZ0Z_13 ));
    Odrv12 I__13131 (
            .O(N__58406),
            .I(\ALU.a_15_sZ0Z_13 ));
    Odrv12 I__13130 (
            .O(N__58403),
            .I(\ALU.a_15_sZ0Z_13 ));
    Odrv4 I__13129 (
            .O(N__58396),
            .I(\ALU.a_15_sZ0Z_13 ));
    Odrv12 I__13128 (
            .O(N__58393),
            .I(\ALU.a_15_sZ0Z_13 ));
    Odrv4 I__13127 (
            .O(N__58390),
            .I(\ALU.a_15_sZ0Z_13 ));
    CascadeMux I__13126 (
            .O(N__58373),
            .I(N__58367));
    InMux I__13125 (
            .O(N__58372),
            .I(N__58362));
    InMux I__13124 (
            .O(N__58371),
            .I(N__58359));
    InMux I__13123 (
            .O(N__58370),
            .I(N__58356));
    InMux I__13122 (
            .O(N__58367),
            .I(N__58353));
    InMux I__13121 (
            .O(N__58366),
            .I(N__58350));
    InMux I__13120 (
            .O(N__58365),
            .I(N__58347));
    LocalMux I__13119 (
            .O(N__58362),
            .I(N__58344));
    LocalMux I__13118 (
            .O(N__58359),
            .I(N__58340));
    LocalMux I__13117 (
            .O(N__58356),
            .I(N__58337));
    LocalMux I__13116 (
            .O(N__58353),
            .I(N__58330));
    LocalMux I__13115 (
            .O(N__58350),
            .I(N__58330));
    LocalMux I__13114 (
            .O(N__58347),
            .I(N__58330));
    Span4Mux_h I__13113 (
            .O(N__58344),
            .I(N__58327));
    InMux I__13112 (
            .O(N__58343),
            .I(N__58324));
    Span4Mux_h I__13111 (
            .O(N__58340),
            .I(N__58321));
    Span4Mux_h I__13110 (
            .O(N__58337),
            .I(N__58318));
    Span4Mux_v I__13109 (
            .O(N__58330),
            .I(N__58315));
    Span4Mux_h I__13108 (
            .O(N__58327),
            .I(N__58312));
    LocalMux I__13107 (
            .O(N__58324),
            .I(\ALU.c_RNIO0KOKEZ0Z_10 ));
    Odrv4 I__13106 (
            .O(N__58321),
            .I(\ALU.c_RNIO0KOKEZ0Z_10 ));
    Odrv4 I__13105 (
            .O(N__58318),
            .I(\ALU.c_RNIO0KOKEZ0Z_10 ));
    Odrv4 I__13104 (
            .O(N__58315),
            .I(\ALU.c_RNIO0KOKEZ0Z_10 ));
    Odrv4 I__13103 (
            .O(N__58312),
            .I(\ALU.c_RNIO0KOKEZ0Z_10 ));
    InMux I__13102 (
            .O(N__58301),
            .I(N__58296));
    InMux I__13101 (
            .O(N__58300),
            .I(N__58291));
    InMux I__13100 (
            .O(N__58299),
            .I(N__58288));
    LocalMux I__13099 (
            .O(N__58296),
            .I(N__58285));
    InMux I__13098 (
            .O(N__58295),
            .I(N__58280));
    InMux I__13097 (
            .O(N__58294),
            .I(N__58277));
    LocalMux I__13096 (
            .O(N__58291),
            .I(N__58274));
    LocalMux I__13095 (
            .O(N__58288),
            .I(N__58271));
    Span4Mux_v I__13094 (
            .O(N__58285),
            .I(N__58268));
    InMux I__13093 (
            .O(N__58284),
            .I(N__58265));
    InMux I__13092 (
            .O(N__58283),
            .I(N__58262));
    LocalMux I__13091 (
            .O(N__58280),
            .I(N__58255));
    LocalMux I__13090 (
            .O(N__58277),
            .I(N__58255));
    Span4Mux_h I__13089 (
            .O(N__58274),
            .I(N__58255));
    Span4Mux_v I__13088 (
            .O(N__58271),
            .I(N__58250));
    Span4Mux_h I__13087 (
            .O(N__58268),
            .I(N__58250));
    LocalMux I__13086 (
            .O(N__58265),
            .I(\ALU.mult_549_c_RNIE7260OZ0 ));
    LocalMux I__13085 (
            .O(N__58262),
            .I(\ALU.mult_549_c_RNIE7260OZ0 ));
    Odrv4 I__13084 (
            .O(N__58255),
            .I(\ALU.mult_549_c_RNIE7260OZ0 ));
    Odrv4 I__13083 (
            .O(N__58250),
            .I(\ALU.mult_549_c_RNIE7260OZ0 ));
    CascadeMux I__13082 (
            .O(N__58241),
            .I(N__58238));
    InMux I__13081 (
            .O(N__58238),
            .I(N__58235));
    LocalMux I__13080 (
            .O(N__58235),
            .I(N__58231));
    InMux I__13079 (
            .O(N__58234),
            .I(N__58228));
    Span4Mux_v I__13078 (
            .O(N__58231),
            .I(N__58222));
    LocalMux I__13077 (
            .O(N__58228),
            .I(N__58222));
    InMux I__13076 (
            .O(N__58227),
            .I(N__58219));
    Span4Mux_v I__13075 (
            .O(N__58222),
            .I(N__58216));
    LocalMux I__13074 (
            .O(N__58219),
            .I(N__58213));
    Span4Mux_h I__13073 (
            .O(N__58216),
            .I(N__58210));
    Span4Mux_v I__13072 (
            .O(N__58213),
            .I(N__58207));
    Sp12to4 I__13071 (
            .O(N__58210),
            .I(N__58202));
    Sp12to4 I__13070 (
            .O(N__58207),
            .I(N__58202));
    Span12Mux_h I__13069 (
            .O(N__58202),
            .I(N__58199));
    Odrv12 I__13068 (
            .O(N__58199),
            .I(h_10));
    InMux I__13067 (
            .O(N__58196),
            .I(N__58191));
    InMux I__13066 (
            .O(N__58195),
            .I(N__58185));
    InMux I__13065 (
            .O(N__58194),
            .I(N__58181));
    LocalMux I__13064 (
            .O(N__58191),
            .I(N__58178));
    InMux I__13063 (
            .O(N__58190),
            .I(N__58175));
    InMux I__13062 (
            .O(N__58189),
            .I(N__58172));
    InMux I__13061 (
            .O(N__58188),
            .I(N__58169));
    LocalMux I__13060 (
            .O(N__58185),
            .I(N__58166));
    InMux I__13059 (
            .O(N__58184),
            .I(N__58162));
    LocalMux I__13058 (
            .O(N__58181),
            .I(N__58159));
    Span4Mux_v I__13057 (
            .O(N__58178),
            .I(N__58150));
    LocalMux I__13056 (
            .O(N__58175),
            .I(N__58150));
    LocalMux I__13055 (
            .O(N__58172),
            .I(N__58150));
    LocalMux I__13054 (
            .O(N__58169),
            .I(N__58150));
    Span4Mux_v I__13053 (
            .O(N__58166),
            .I(N__58147));
    InMux I__13052 (
            .O(N__58165),
            .I(N__58144));
    LocalMux I__13051 (
            .O(N__58162),
            .I(N__58139));
    Span4Mux_h I__13050 (
            .O(N__58159),
            .I(N__58139));
    Span4Mux_v I__13049 (
            .O(N__58150),
            .I(N__58134));
    Span4Mux_h I__13048 (
            .O(N__58147),
            .I(N__58134));
    LocalMux I__13047 (
            .O(N__58144),
            .I(\ALU.c_RNIBN2FN8Z0Z_11 ));
    Odrv4 I__13046 (
            .O(N__58139),
            .I(\ALU.c_RNIBN2FN8Z0Z_11 ));
    Odrv4 I__13045 (
            .O(N__58134),
            .I(\ALU.c_RNIBN2FN8Z0Z_11 ));
    CascadeMux I__13044 (
            .O(N__58127),
            .I(N__58123));
    CascadeMux I__13043 (
            .O(N__58126),
            .I(N__58120));
    InMux I__13042 (
            .O(N__58123),
            .I(N__58115));
    InMux I__13041 (
            .O(N__58120),
            .I(N__58112));
    InMux I__13040 (
            .O(N__58119),
            .I(N__58105));
    InMux I__13039 (
            .O(N__58118),
            .I(N__58102));
    LocalMux I__13038 (
            .O(N__58115),
            .I(N__58099));
    LocalMux I__13037 (
            .O(N__58112),
            .I(N__58096));
    InMux I__13036 (
            .O(N__58111),
            .I(N__58093));
    InMux I__13035 (
            .O(N__58110),
            .I(N__58090));
    InMux I__13034 (
            .O(N__58109),
            .I(N__58087));
    InMux I__13033 (
            .O(N__58108),
            .I(N__58084));
    LocalMux I__13032 (
            .O(N__58105),
            .I(N__58081));
    LocalMux I__13031 (
            .O(N__58102),
            .I(N__58076));
    Span4Mux_h I__13030 (
            .O(N__58099),
            .I(N__58076));
    Span4Mux_h I__13029 (
            .O(N__58096),
            .I(N__58073));
    LocalMux I__13028 (
            .O(N__58093),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ));
    LocalMux I__13027 (
            .O(N__58090),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ));
    LocalMux I__13026 (
            .O(N__58087),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ));
    LocalMux I__13025 (
            .O(N__58084),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ));
    Odrv4 I__13024 (
            .O(N__58081),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ));
    Odrv4 I__13023 (
            .O(N__58076),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ));
    Odrv4 I__13022 (
            .O(N__58073),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ));
    InMux I__13021 (
            .O(N__58058),
            .I(N__58053));
    InMux I__13020 (
            .O(N__58057),
            .I(N__58046));
    InMux I__13019 (
            .O(N__58056),
            .I(N__58043));
    LocalMux I__13018 (
            .O(N__58053),
            .I(N__58040));
    InMux I__13017 (
            .O(N__58052),
            .I(N__58037));
    InMux I__13016 (
            .O(N__58051),
            .I(N__58034));
    InMux I__13015 (
            .O(N__58050),
            .I(N__58031));
    InMux I__13014 (
            .O(N__58049),
            .I(N__58028));
    LocalMux I__13013 (
            .O(N__58046),
            .I(N__58025));
    LocalMux I__13012 (
            .O(N__58043),
            .I(N__58022));
    Span4Mux_v I__13011 (
            .O(N__58040),
            .I(N__58019));
    LocalMux I__13010 (
            .O(N__58037),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0 ));
    LocalMux I__13009 (
            .O(N__58034),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0 ));
    LocalMux I__13008 (
            .O(N__58031),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0 ));
    LocalMux I__13007 (
            .O(N__58028),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0 ));
    Odrv4 I__13006 (
            .O(N__58025),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0 ));
    Odrv12 I__13005 (
            .O(N__58022),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0 ));
    Odrv4 I__13004 (
            .O(N__58019),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0 ));
    CascadeMux I__13003 (
            .O(N__58004),
            .I(N__58001));
    InMux I__13002 (
            .O(N__58001),
            .I(N__57998));
    LocalMux I__13001 (
            .O(N__57998),
            .I(N__57994));
    InMux I__13000 (
            .O(N__57997),
            .I(N__57991));
    Span4Mux_v I__12999 (
            .O(N__57994),
            .I(N__57988));
    LocalMux I__12998 (
            .O(N__57991),
            .I(N__57985));
    Span4Mux_h I__12997 (
            .O(N__57988),
            .I(N__57982));
    Span4Mux_v I__12996 (
            .O(N__57985),
            .I(N__57978));
    Span4Mux_v I__12995 (
            .O(N__57982),
            .I(N__57975));
    InMux I__12994 (
            .O(N__57981),
            .I(N__57972));
    Span4Mux_h I__12993 (
            .O(N__57978),
            .I(N__57969));
    Sp12to4 I__12992 (
            .O(N__57975),
            .I(N__57964));
    LocalMux I__12991 (
            .O(N__57972),
            .I(N__57964));
    Span4Mux_h I__12990 (
            .O(N__57969),
            .I(N__57961));
    Span12Mux_h I__12989 (
            .O(N__57964),
            .I(N__57958));
    Span4Mux_v I__12988 (
            .O(N__57961),
            .I(N__57955));
    Odrv12 I__12987 (
            .O(N__57958),
            .I(h_11));
    Odrv4 I__12986 (
            .O(N__57955),
            .I(h_11));
    InMux I__12985 (
            .O(N__57950),
            .I(N__57947));
    LocalMux I__12984 (
            .O(N__57947),
            .I(N__57943));
    InMux I__12983 (
            .O(N__57946),
            .I(N__57940));
    Span4Mux_v I__12982 (
            .O(N__57943),
            .I(N__57935));
    LocalMux I__12981 (
            .O(N__57940),
            .I(N__57935));
    Span4Mux_v I__12980 (
            .O(N__57935),
            .I(N__57931));
    InMux I__12979 (
            .O(N__57934),
            .I(N__57928));
    Span4Mux_h I__12978 (
            .O(N__57931),
            .I(N__57925));
    LocalMux I__12977 (
            .O(N__57928),
            .I(N__57922));
    Span4Mux_h I__12976 (
            .O(N__57925),
            .I(N__57917));
    Span4Mux_v I__12975 (
            .O(N__57922),
            .I(N__57917));
    Sp12to4 I__12974 (
            .O(N__57917),
            .I(N__57914));
    Span12Mux_h I__12973 (
            .O(N__57914),
            .I(N__57911));
    Odrv12 I__12972 (
            .O(N__57911),
            .I(h_12));
    InMux I__12971 (
            .O(N__57908),
            .I(N__57905));
    LocalMux I__12970 (
            .O(N__57905),
            .I(N__57902));
    Span4Mux_v I__12969 (
            .O(N__57902),
            .I(N__57899));
    Span4Mux_h I__12968 (
            .O(N__57899),
            .I(N__57896));
    Span4Mux_v I__12967 (
            .O(N__57896),
            .I(N__57893));
    Sp12to4 I__12966 (
            .O(N__57893),
            .I(N__57888));
    InMux I__12965 (
            .O(N__57892),
            .I(N__57885));
    InMux I__12964 (
            .O(N__57891),
            .I(N__57882));
    Span12Mux_h I__12963 (
            .O(N__57888),
            .I(N__57877));
    LocalMux I__12962 (
            .O(N__57885),
            .I(N__57877));
    LocalMux I__12961 (
            .O(N__57882),
            .I(N__57872));
    Span12Mux_v I__12960 (
            .O(N__57877),
            .I(N__57872));
    Odrv12 I__12959 (
            .O(N__57872),
            .I(h_13));
    CascadeMux I__12958 (
            .O(N__57869),
            .I(N__57866));
    InMux I__12957 (
            .O(N__57866),
            .I(N__57863));
    LocalMux I__12956 (
            .O(N__57863),
            .I(N__57860));
    Span4Mux_v I__12955 (
            .O(N__57860),
            .I(N__57856));
    InMux I__12954 (
            .O(N__57859),
            .I(N__57853));
    Span4Mux_h I__12953 (
            .O(N__57856),
            .I(N__57849));
    LocalMux I__12952 (
            .O(N__57853),
            .I(N__57846));
    InMux I__12951 (
            .O(N__57852),
            .I(N__57843));
    Span4Mux_h I__12950 (
            .O(N__57849),
            .I(N__57840));
    Span4Mux_v I__12949 (
            .O(N__57846),
            .I(N__57835));
    LocalMux I__12948 (
            .O(N__57843),
            .I(N__57835));
    Span4Mux_h I__12947 (
            .O(N__57840),
            .I(N__57830));
    Span4Mux_h I__12946 (
            .O(N__57835),
            .I(N__57830));
    Span4Mux_h I__12945 (
            .O(N__57830),
            .I(N__57827));
    Span4Mux_h I__12944 (
            .O(N__57827),
            .I(N__57824));
    Odrv4 I__12943 (
            .O(N__57824),
            .I(h_14));
    InMux I__12942 (
            .O(N__57821),
            .I(N__57816));
    InMux I__12941 (
            .O(N__57820),
            .I(N__57813));
    InMux I__12940 (
            .O(N__57819),
            .I(N__57810));
    LocalMux I__12939 (
            .O(N__57816),
            .I(N__57805));
    LocalMux I__12938 (
            .O(N__57813),
            .I(N__57802));
    LocalMux I__12937 (
            .O(N__57810),
            .I(N__57798));
    InMux I__12936 (
            .O(N__57809),
            .I(N__57793));
    InMux I__12935 (
            .O(N__57808),
            .I(N__57793));
    Span4Mux_v I__12934 (
            .O(N__57805),
            .I(N__57788));
    Span4Mux_v I__12933 (
            .O(N__57802),
            .I(N__57785));
    InMux I__12932 (
            .O(N__57801),
            .I(N__57782));
    Span4Mux_h I__12931 (
            .O(N__57798),
            .I(N__57777));
    LocalMux I__12930 (
            .O(N__57793),
            .I(N__57777));
    InMux I__12929 (
            .O(N__57792),
            .I(N__57774));
    InMux I__12928 (
            .O(N__57791),
            .I(N__57771));
    Span4Mux_v I__12927 (
            .O(N__57788),
            .I(N__57768));
    Sp12to4 I__12926 (
            .O(N__57785),
            .I(N__57765));
    LocalMux I__12925 (
            .O(N__57782),
            .I(N__57762));
    Span4Mux_v I__12924 (
            .O(N__57777),
            .I(N__57758));
    LocalMux I__12923 (
            .O(N__57774),
            .I(N__57755));
    LocalMux I__12922 (
            .O(N__57771),
            .I(N__57752));
    Span4Mux_v I__12921 (
            .O(N__57768),
            .I(N__57748));
    Span12Mux_h I__12920 (
            .O(N__57765),
            .I(N__57743));
    Sp12to4 I__12919 (
            .O(N__57762),
            .I(N__57743));
    InMux I__12918 (
            .O(N__57761),
            .I(N__57740));
    Sp12to4 I__12917 (
            .O(N__57758),
            .I(N__57737));
    Span4Mux_h I__12916 (
            .O(N__57755),
            .I(N__57732));
    Span4Mux_h I__12915 (
            .O(N__57752),
            .I(N__57732));
    InMux I__12914 (
            .O(N__57751),
            .I(N__57729));
    Span4Mux_h I__12913 (
            .O(N__57748),
            .I(N__57725));
    Span12Mux_v I__12912 (
            .O(N__57743),
            .I(N__57722));
    LocalMux I__12911 (
            .O(N__57740),
            .I(N__57715));
    Span12Mux_h I__12910 (
            .O(N__57737),
            .I(N__57715));
    Sp12to4 I__12909 (
            .O(N__57732),
            .I(N__57715));
    LocalMux I__12908 (
            .O(N__57729),
            .I(N__57712));
    InMux I__12907 (
            .O(N__57728),
            .I(N__57709));
    Span4Mux_v I__12906 (
            .O(N__57725),
            .I(N__57706));
    Span12Mux_h I__12905 (
            .O(N__57722),
            .I(N__57703));
    Span12Mux_v I__12904 (
            .O(N__57715),
            .I(N__57700));
    Span4Mux_h I__12903 (
            .O(N__57712),
            .I(N__57697));
    LocalMux I__12902 (
            .O(N__57709),
            .I(\CONTROL.addrstack_1 ));
    Odrv4 I__12901 (
            .O(N__57706),
            .I(\CONTROL.addrstack_1 ));
    Odrv12 I__12900 (
            .O(N__57703),
            .I(\CONTROL.addrstack_1 ));
    Odrv12 I__12899 (
            .O(N__57700),
            .I(\CONTROL.addrstack_1 ));
    Odrv4 I__12898 (
            .O(N__57697),
            .I(\CONTROL.addrstack_1 ));
    CascadeMux I__12897 (
            .O(N__57686),
            .I(N__57682));
    InMux I__12896 (
            .O(N__57685),
            .I(N__57679));
    InMux I__12895 (
            .O(N__57682),
            .I(N__57676));
    LocalMux I__12894 (
            .O(N__57679),
            .I(N__57672));
    LocalMux I__12893 (
            .O(N__57676),
            .I(N__57669));
    InMux I__12892 (
            .O(N__57675),
            .I(N__57666));
    Span4Mux_h I__12891 (
            .O(N__57672),
            .I(N__57661));
    Span4Mux_v I__12890 (
            .O(N__57669),
            .I(N__57661));
    LocalMux I__12889 (
            .O(N__57666),
            .I(N__57658));
    Span4Mux_v I__12888 (
            .O(N__57661),
            .I(N__57655));
    Span12Mux_v I__12887 (
            .O(N__57658),
            .I(N__57652));
    Span4Mux_h I__12886 (
            .O(N__57655),
            .I(N__57649));
    Span12Mux_h I__12885 (
            .O(N__57652),
            .I(N__57646));
    Span4Mux_h I__12884 (
            .O(N__57649),
            .I(N__57643));
    Odrv12 I__12883 (
            .O(N__57646),
            .I(f_12));
    Odrv4 I__12882 (
            .O(N__57643),
            .I(f_12));
    CascadeMux I__12881 (
            .O(N__57638),
            .I(N__57635));
    InMux I__12880 (
            .O(N__57635),
            .I(N__57632));
    LocalMux I__12879 (
            .O(N__57632),
            .I(N__57628));
    InMux I__12878 (
            .O(N__57631),
            .I(N__57625));
    Span4Mux_v I__12877 (
            .O(N__57628),
            .I(N__57622));
    LocalMux I__12876 (
            .O(N__57625),
            .I(N__57616));
    Span4Mux_v I__12875 (
            .O(N__57622),
            .I(N__57616));
    InMux I__12874 (
            .O(N__57621),
            .I(N__57613));
    Span4Mux_h I__12873 (
            .O(N__57616),
            .I(N__57610));
    LocalMux I__12872 (
            .O(N__57613),
            .I(N__57607));
    Span4Mux_h I__12871 (
            .O(N__57610),
            .I(N__57604));
    Span12Mux_h I__12870 (
            .O(N__57607),
            .I(N__57601));
    Span4Mux_h I__12869 (
            .O(N__57604),
            .I(N__57598));
    Odrv12 I__12868 (
            .O(N__57601),
            .I(f_13));
    Odrv4 I__12867 (
            .O(N__57598),
            .I(f_13));
    CascadeMux I__12866 (
            .O(N__57593),
            .I(N__57590));
    InMux I__12865 (
            .O(N__57590),
            .I(N__57587));
    LocalMux I__12864 (
            .O(N__57587),
            .I(N__57583));
    CascadeMux I__12863 (
            .O(N__57586),
            .I(N__57579));
    Span4Mux_v I__12862 (
            .O(N__57583),
            .I(N__57576));
    InMux I__12861 (
            .O(N__57582),
            .I(N__57573));
    InMux I__12860 (
            .O(N__57579),
            .I(N__57570));
    Span4Mux_h I__12859 (
            .O(N__57576),
            .I(N__57567));
    LocalMux I__12858 (
            .O(N__57573),
            .I(N__57564));
    LocalMux I__12857 (
            .O(N__57570),
            .I(N__57561));
    Sp12to4 I__12856 (
            .O(N__57567),
            .I(N__57558));
    Span4Mux_h I__12855 (
            .O(N__57564),
            .I(N__57555));
    Span4Mux_v I__12854 (
            .O(N__57561),
            .I(N__57552));
    Span12Mux_s9_v I__12853 (
            .O(N__57558),
            .I(N__57549));
    Span4Mux_h I__12852 (
            .O(N__57555),
            .I(N__57546));
    Span4Mux_h I__12851 (
            .O(N__57552),
            .I(N__57543));
    Span12Mux_v I__12850 (
            .O(N__57549),
            .I(N__57540));
    Span4Mux_v I__12849 (
            .O(N__57546),
            .I(N__57537));
    Span4Mux_v I__12848 (
            .O(N__57543),
            .I(N__57534));
    Odrv12 I__12847 (
            .O(N__57540),
            .I(f_14));
    Odrv4 I__12846 (
            .O(N__57537),
            .I(f_14));
    Odrv4 I__12845 (
            .O(N__57534),
            .I(f_14));
    CascadeMux I__12844 (
            .O(N__57527),
            .I(N__57524));
    InMux I__12843 (
            .O(N__57524),
            .I(N__57518));
    InMux I__12842 (
            .O(N__57523),
            .I(N__57518));
    LocalMux I__12841 (
            .O(N__57518),
            .I(N__57515));
    Span4Mux_v I__12840 (
            .O(N__57515),
            .I(N__57511));
    InMux I__12839 (
            .O(N__57514),
            .I(N__57508));
    Odrv4 I__12838 (
            .O(N__57511),
            .I(\ALU.log_1_14 ));
    LocalMux I__12837 (
            .O(N__57508),
            .I(\ALU.log_1_14 ));
    InMux I__12836 (
            .O(N__57503),
            .I(N__57500));
    LocalMux I__12835 (
            .O(N__57500),
            .I(N__57497));
    Span4Mux_h I__12834 (
            .O(N__57497),
            .I(N__57494));
    Span4Mux_h I__12833 (
            .O(N__57494),
            .I(N__57491));
    Odrv4 I__12832 (
            .O(N__57491),
            .I(\ALU.a_15_m0_14 ));
    CascadeMux I__12831 (
            .O(N__57488),
            .I(\ALU.addsub_cry_13_c_RNIBVHEA1Z0Z_0_cascade_ ));
    InMux I__12830 (
            .O(N__57485),
            .I(N__57482));
    LocalMux I__12829 (
            .O(N__57482),
            .I(\ALU.addsub_cry_13_c_RNIBVHEAZ0Z1 ));
    CascadeMux I__12828 (
            .O(N__57479),
            .I(\ALU.addsub_cry_13_c_RNIJMTGAZ0Z5_cascade_ ));
    InMux I__12827 (
            .O(N__57476),
            .I(N__57473));
    LocalMux I__12826 (
            .O(N__57473),
            .I(N__57470));
    Span4Mux_h I__12825 (
            .O(N__57470),
            .I(N__57467));
    Span4Mux_h I__12824 (
            .O(N__57467),
            .I(N__57464));
    Odrv4 I__12823 (
            .O(N__57464),
            .I(\ALU.mult_14 ));
    CascadeMux I__12822 (
            .O(N__57461),
            .I(\ALU.a_15_ns_rn_0_14_cascade_ ));
    InMux I__12821 (
            .O(N__57458),
            .I(N__57455));
    LocalMux I__12820 (
            .O(N__57455),
            .I(N__57451));
    InMux I__12819 (
            .O(N__57454),
            .I(N__57448));
    Span4Mux_v I__12818 (
            .O(N__57451),
            .I(N__57445));
    LocalMux I__12817 (
            .O(N__57448),
            .I(N__57442));
    Span4Mux_h I__12816 (
            .O(N__57445),
            .I(N__57439));
    Span4Mux_h I__12815 (
            .O(N__57442),
            .I(N__57436));
    Span4Mux_h I__12814 (
            .O(N__57439),
            .I(N__57433));
    Span4Mux_v I__12813 (
            .O(N__57436),
            .I(N__57430));
    Span4Mux_v I__12812 (
            .O(N__57433),
            .I(N__57427));
    Odrv4 I__12811 (
            .O(N__57430),
            .I(\ALU.aZ0Z_14 ));
    Odrv4 I__12810 (
            .O(N__57427),
            .I(\ALU.aZ0Z_14 ));
    InMux I__12809 (
            .O(N__57422),
            .I(N__57416));
    InMux I__12808 (
            .O(N__57421),
            .I(N__57413));
    InMux I__12807 (
            .O(N__57420),
            .I(N__57407));
    InMux I__12806 (
            .O(N__57419),
            .I(N__57407));
    LocalMux I__12805 (
            .O(N__57416),
            .I(N__57400));
    LocalMux I__12804 (
            .O(N__57413),
            .I(N__57400));
    CascadeMux I__12803 (
            .O(N__57412),
            .I(N__57397));
    LocalMux I__12802 (
            .O(N__57407),
            .I(N__57393));
    InMux I__12801 (
            .O(N__57406),
            .I(N__57390));
    CascadeMux I__12800 (
            .O(N__57405),
            .I(N__57385));
    Span4Mux_h I__12799 (
            .O(N__57400),
            .I(N__57379));
    InMux I__12798 (
            .O(N__57397),
            .I(N__57373));
    InMux I__12797 (
            .O(N__57396),
            .I(N__57373));
    Span4Mux_v I__12796 (
            .O(N__57393),
            .I(N__57368));
    LocalMux I__12795 (
            .O(N__57390),
            .I(N__57365));
    InMux I__12794 (
            .O(N__57389),
            .I(N__57360));
    InMux I__12793 (
            .O(N__57388),
            .I(N__57360));
    InMux I__12792 (
            .O(N__57385),
            .I(N__57355));
    InMux I__12791 (
            .O(N__57384),
            .I(N__57355));
    CascadeMux I__12790 (
            .O(N__57383),
            .I(N__57352));
    InMux I__12789 (
            .O(N__57382),
            .I(N__57346));
    Span4Mux_h I__12788 (
            .O(N__57379),
            .I(N__57343));
    InMux I__12787 (
            .O(N__57378),
            .I(N__57340));
    LocalMux I__12786 (
            .O(N__57373),
            .I(N__57337));
    InMux I__12785 (
            .O(N__57372),
            .I(N__57332));
    InMux I__12784 (
            .O(N__57371),
            .I(N__57332));
    Span4Mux_h I__12783 (
            .O(N__57368),
            .I(N__57329));
    Span4Mux_h I__12782 (
            .O(N__57365),
            .I(N__57322));
    LocalMux I__12781 (
            .O(N__57360),
            .I(N__57322));
    LocalMux I__12780 (
            .O(N__57355),
            .I(N__57322));
    InMux I__12779 (
            .O(N__57352),
            .I(N__57316));
    InMux I__12778 (
            .O(N__57351),
            .I(N__57316));
    InMux I__12777 (
            .O(N__57350),
            .I(N__57311));
    InMux I__12776 (
            .O(N__57349),
            .I(N__57311));
    LocalMux I__12775 (
            .O(N__57346),
            .I(N__57300));
    Span4Mux_v I__12774 (
            .O(N__57343),
            .I(N__57300));
    LocalMux I__12773 (
            .O(N__57340),
            .I(N__57300));
    Span4Mux_v I__12772 (
            .O(N__57337),
            .I(N__57300));
    LocalMux I__12771 (
            .O(N__57332),
            .I(N__57300));
    Span4Mux_v I__12770 (
            .O(N__57329),
            .I(N__57295));
    Span4Mux_h I__12769 (
            .O(N__57322),
            .I(N__57295));
    InMux I__12768 (
            .O(N__57321),
            .I(N__57292));
    LocalMux I__12767 (
            .O(N__57316),
            .I(N__57285));
    LocalMux I__12766 (
            .O(N__57311),
            .I(N__57285));
    Span4Mux_v I__12765 (
            .O(N__57300),
            .I(N__57285));
    Span4Mux_h I__12764 (
            .O(N__57295),
            .I(N__57282));
    LocalMux I__12763 (
            .O(N__57292),
            .I(N__57279));
    Span4Mux_h I__12762 (
            .O(N__57285),
            .I(N__57276));
    Span4Mux_h I__12761 (
            .O(N__57282),
            .I(N__57273));
    Sp12to4 I__12760 (
            .O(N__57279),
            .I(N__57270));
    Span4Mux_h I__12759 (
            .O(N__57276),
            .I(N__57267));
    Sp12to4 I__12758 (
            .O(N__57273),
            .I(N__57264));
    Span12Mux_s11_v I__12757 (
            .O(N__57270),
            .I(N__57261));
    Span4Mux_h I__12756 (
            .O(N__57267),
            .I(N__57258));
    Span12Mux_s11_v I__12755 (
            .O(N__57264),
            .I(N__57255));
    Odrv12 I__12754 (
            .O(N__57261),
            .I(\ALU.a_15_sZ0Z_3 ));
    Odrv4 I__12753 (
            .O(N__57258),
            .I(\ALU.a_15_sZ0Z_3 ));
    Odrv12 I__12752 (
            .O(N__57255),
            .I(\ALU.a_15_sZ0Z_3 ));
    InMux I__12751 (
            .O(N__57248),
            .I(N__57245));
    LocalMux I__12750 (
            .O(N__57245),
            .I(\ALU.log_1_3 ));
    InMux I__12749 (
            .O(N__57242),
            .I(N__57239));
    LocalMux I__12748 (
            .O(N__57239),
            .I(N__57235));
    InMux I__12747 (
            .O(N__57238),
            .I(N__57232));
    Span4Mux_h I__12746 (
            .O(N__57235),
            .I(N__57228));
    LocalMux I__12745 (
            .O(N__57232),
            .I(N__57224));
    InMux I__12744 (
            .O(N__57231),
            .I(N__57221));
    Span4Mux_v I__12743 (
            .O(N__57228),
            .I(N__57218));
    InMux I__12742 (
            .O(N__57227),
            .I(N__57215));
    Span4Mux_v I__12741 (
            .O(N__57224),
            .I(N__57212));
    LocalMux I__12740 (
            .O(N__57221),
            .I(N__57209));
    Span4Mux_h I__12739 (
            .O(N__57218),
            .I(N__57204));
    LocalMux I__12738 (
            .O(N__57215),
            .I(N__57204));
    Span4Mux_v I__12737 (
            .O(N__57212),
            .I(N__57199));
    Span4Mux_h I__12736 (
            .O(N__57209),
            .I(N__57199));
    Span4Mux_h I__12735 (
            .O(N__57204),
            .I(N__57196));
    Span4Mux_v I__12734 (
            .O(N__57199),
            .I(N__57193));
    Span4Mux_h I__12733 (
            .O(N__57196),
            .I(N__57190));
    Odrv4 I__12732 (
            .O(N__57193),
            .I(\ALU.lshift62_2 ));
    Odrv4 I__12731 (
            .O(N__57190),
            .I(\ALU.lshift62_2 ));
    InMux I__12730 (
            .O(N__57185),
            .I(N__57182));
    LocalMux I__12729 (
            .O(N__57182),
            .I(N__57179));
    Odrv12 I__12728 (
            .O(N__57179),
            .I(\ALU.mult_558_c_RNIB3E8DCZ0 ));
    CascadeMux I__12727 (
            .O(N__57176),
            .I(\ALU.a_15_d_ns_1_13_cascade_ ));
    CascadeMux I__12726 (
            .O(N__57173),
            .I(\ALU.mult_558_c_RNIB75F9GZ0_cascade_ ));
    InMux I__12725 (
            .O(N__57170),
            .I(N__57167));
    LocalMux I__12724 (
            .O(N__57167),
            .I(N__57163));
    InMux I__12723 (
            .O(N__57166),
            .I(N__57160));
    Span4Mux_v I__12722 (
            .O(N__57163),
            .I(N__57157));
    LocalMux I__12721 (
            .O(N__57160),
            .I(N__57154));
    Span4Mux_h I__12720 (
            .O(N__57157),
            .I(N__57151));
    Span4Mux_v I__12719 (
            .O(N__57154),
            .I(N__57148));
    Span4Mux_v I__12718 (
            .O(N__57151),
            .I(N__57145));
    Sp12to4 I__12717 (
            .O(N__57148),
            .I(N__57142));
    Sp12to4 I__12716 (
            .O(N__57145),
            .I(N__57137));
    Span12Mux_h I__12715 (
            .O(N__57142),
            .I(N__57137));
    Odrv12 I__12714 (
            .O(N__57137),
            .I(\ALU.aZ0Z_13 ));
    InMux I__12713 (
            .O(N__57134),
            .I(N__57131));
    LocalMux I__12712 (
            .O(N__57131),
            .I(N__57128));
    Span4Mux_v I__12711 (
            .O(N__57128),
            .I(N__57125));
    Odrv4 I__12710 (
            .O(N__57125),
            .I(\ALU.d_RNIJ7J1M5_0Z0Z_2 ));
    CascadeMux I__12709 (
            .O(N__57122),
            .I(N__57118));
    InMux I__12708 (
            .O(N__57121),
            .I(N__57113));
    InMux I__12707 (
            .O(N__57118),
            .I(N__57113));
    LocalMux I__12706 (
            .O(N__57113),
            .I(\ALU.a_15_m3_d_sZ0Z_8 ));
    InMux I__12705 (
            .O(N__57110),
            .I(N__57104));
    InMux I__12704 (
            .O(N__57109),
            .I(N__57104));
    LocalMux I__12703 (
            .O(N__57104),
            .I(N__57101));
    Span4Mux_v I__12702 (
            .O(N__57101),
            .I(N__57098));
    Span4Mux_v I__12701 (
            .O(N__57098),
            .I(N__57095));
    Sp12to4 I__12700 (
            .O(N__57095),
            .I(N__57091));
    InMux I__12699 (
            .O(N__57094),
            .I(N__57088));
    Span12Mux_h I__12698 (
            .O(N__57091),
            .I(N__57085));
    LocalMux I__12697 (
            .O(N__57088),
            .I(N__57082));
    Odrv12 I__12696 (
            .O(N__57085),
            .I(bus_0_8));
    Odrv4 I__12695 (
            .O(N__57082),
            .I(bus_0_8));
    CascadeMux I__12694 (
            .O(N__57077),
            .I(\ALU.a_15_m3_d_sZ0Z_8_cascade_ ));
    InMux I__12693 (
            .O(N__57074),
            .I(N__57068));
    InMux I__12692 (
            .O(N__57073),
            .I(N__57068));
    LocalMux I__12691 (
            .O(N__57068),
            .I(\ALU.d_RNI12L8C5Z0Z_2 ));
    InMux I__12690 (
            .O(N__57065),
            .I(N__57062));
    LocalMux I__12689 (
            .O(N__57062),
            .I(N__57059));
    Span4Mux_v I__12688 (
            .O(N__57059),
            .I(N__57056));
    Odrv4 I__12687 (
            .O(N__57056),
            .I(\ALU.d_RNIJ7J1M5Z0Z_2 ));
    InMux I__12686 (
            .O(N__57053),
            .I(N__57050));
    LocalMux I__12685 (
            .O(N__57050),
            .I(N__57047));
    Span4Mux_h I__12684 (
            .O(N__57047),
            .I(N__57043));
    InMux I__12683 (
            .O(N__57046),
            .I(N__57040));
    Span4Mux_h I__12682 (
            .O(N__57043),
            .I(N__57034));
    LocalMux I__12681 (
            .O(N__57040),
            .I(N__57034));
    InMux I__12680 (
            .O(N__57039),
            .I(N__57025));
    Span4Mux_v I__12679 (
            .O(N__57034),
            .I(N__57021));
    InMux I__12678 (
            .O(N__57033),
            .I(N__57016));
    InMux I__12677 (
            .O(N__57032),
            .I(N__57016));
    InMux I__12676 (
            .O(N__57031),
            .I(N__57012));
    CascadeMux I__12675 (
            .O(N__57030),
            .I(N__57009));
    CascadeMux I__12674 (
            .O(N__57029),
            .I(N__57006));
    CascadeMux I__12673 (
            .O(N__57028),
            .I(N__57003));
    LocalMux I__12672 (
            .O(N__57025),
            .I(N__57000));
    CascadeMux I__12671 (
            .O(N__57024),
            .I(N__56997));
    Span4Mux_v I__12670 (
            .O(N__57021),
            .I(N__56994));
    LocalMux I__12669 (
            .O(N__57016),
            .I(N__56991));
    InMux I__12668 (
            .O(N__57015),
            .I(N__56988));
    LocalMux I__12667 (
            .O(N__57012),
            .I(N__56984));
    InMux I__12666 (
            .O(N__57009),
            .I(N__56977));
    InMux I__12665 (
            .O(N__57006),
            .I(N__56977));
    InMux I__12664 (
            .O(N__57003),
            .I(N__56977));
    Span4Mux_h I__12663 (
            .O(N__57000),
            .I(N__56974));
    InMux I__12662 (
            .O(N__56997),
            .I(N__56971));
    Span4Mux_h I__12661 (
            .O(N__56994),
            .I(N__56966));
    Span4Mux_v I__12660 (
            .O(N__56991),
            .I(N__56966));
    LocalMux I__12659 (
            .O(N__56988),
            .I(N__56963));
    InMux I__12658 (
            .O(N__56987),
            .I(N__56960));
    Span4Mux_h I__12657 (
            .O(N__56984),
            .I(N__56955));
    LocalMux I__12656 (
            .O(N__56977),
            .I(N__56955));
    Odrv4 I__12655 (
            .O(N__56974),
            .I(\ALU.status_19_10 ));
    LocalMux I__12654 (
            .O(N__56971),
            .I(\ALU.status_19_10 ));
    Odrv4 I__12653 (
            .O(N__56966),
            .I(\ALU.status_19_10 ));
    Odrv12 I__12652 (
            .O(N__56963),
            .I(\ALU.status_19_10 ));
    LocalMux I__12651 (
            .O(N__56960),
            .I(\ALU.status_19_10 ));
    Odrv4 I__12650 (
            .O(N__56955),
            .I(\ALU.status_19_10 ));
    CascadeMux I__12649 (
            .O(N__56942),
            .I(N__56939));
    InMux I__12648 (
            .O(N__56939),
            .I(N__56936));
    LocalMux I__12647 (
            .O(N__56936),
            .I(\ALU.aluOut_i_11 ));
    InMux I__12646 (
            .O(N__56933),
            .I(N__56930));
    LocalMux I__12645 (
            .O(N__56930),
            .I(N__56925));
    InMux I__12644 (
            .O(N__56929),
            .I(N__56920));
    InMux I__12643 (
            .O(N__56928),
            .I(N__56920));
    Span4Mux_h I__12642 (
            .O(N__56925),
            .I(N__56917));
    LocalMux I__12641 (
            .O(N__56920),
            .I(N__56914));
    Span4Mux_h I__12640 (
            .O(N__56917),
            .I(N__56911));
    Span4Mux_v I__12639 (
            .O(N__56914),
            .I(N__56906));
    Span4Mux_h I__12638 (
            .O(N__56911),
            .I(N__56901));
    InMux I__12637 (
            .O(N__56910),
            .I(N__56895));
    InMux I__12636 (
            .O(N__56909),
            .I(N__56895));
    Span4Mux_h I__12635 (
            .O(N__56906),
            .I(N__56892));
    InMux I__12634 (
            .O(N__56905),
            .I(N__56889));
    InMux I__12633 (
            .O(N__56904),
            .I(N__56886));
    Span4Mux_h I__12632 (
            .O(N__56901),
            .I(N__56883));
    InMux I__12631 (
            .O(N__56900),
            .I(N__56880));
    LocalMux I__12630 (
            .O(N__56895),
            .I(N__56877));
    Span4Mux_h I__12629 (
            .O(N__56892),
            .I(N__56870));
    LocalMux I__12628 (
            .O(N__56889),
            .I(N__56870));
    LocalMux I__12627 (
            .O(N__56886),
            .I(N__56870));
    Span4Mux_v I__12626 (
            .O(N__56883),
            .I(N__56865));
    LocalMux I__12625 (
            .O(N__56880),
            .I(N__56865));
    Span12Mux_v I__12624 (
            .O(N__56877),
            .I(N__56862));
    Span4Mux_h I__12623 (
            .O(N__56870),
            .I(N__56859));
    Odrv4 I__12622 (
            .O(N__56865),
            .I(\ALU.N_126 ));
    Odrv12 I__12621 (
            .O(N__56862),
            .I(\ALU.N_126 ));
    Odrv4 I__12620 (
            .O(N__56859),
            .I(\ALU.N_126 ));
    CascadeMux I__12619 (
            .O(N__56852),
            .I(N__56849));
    InMux I__12618 (
            .O(N__56849),
            .I(N__56846));
    LocalMux I__12617 (
            .O(N__56846),
            .I(\ALU.aluOut_i_12 ));
    CascadeMux I__12616 (
            .O(N__56843),
            .I(N__56840));
    InMux I__12615 (
            .O(N__56840),
            .I(N__56836));
    CascadeMux I__12614 (
            .O(N__56839),
            .I(N__56833));
    LocalMux I__12613 (
            .O(N__56836),
            .I(N__56830));
    InMux I__12612 (
            .O(N__56833),
            .I(N__56825));
    Span4Mux_v I__12611 (
            .O(N__56830),
            .I(N__56820));
    InMux I__12610 (
            .O(N__56829),
            .I(N__56815));
    InMux I__12609 (
            .O(N__56828),
            .I(N__56815));
    LocalMux I__12608 (
            .O(N__56825),
            .I(N__56812));
    CascadeMux I__12607 (
            .O(N__56824),
            .I(N__56809));
    CascadeMux I__12606 (
            .O(N__56823),
            .I(N__56806));
    Span4Mux_h I__12605 (
            .O(N__56820),
            .I(N__56799));
    LocalMux I__12604 (
            .O(N__56815),
            .I(N__56799));
    Span4Mux_v I__12603 (
            .O(N__56812),
            .I(N__56796));
    InMux I__12602 (
            .O(N__56809),
            .I(N__56793));
    InMux I__12601 (
            .O(N__56806),
            .I(N__56788));
    InMux I__12600 (
            .O(N__56805),
            .I(N__56788));
    CascadeMux I__12599 (
            .O(N__56804),
            .I(N__56784));
    Span4Mux_h I__12598 (
            .O(N__56799),
            .I(N__56781));
    Span4Mux_h I__12597 (
            .O(N__56796),
            .I(N__56778));
    LocalMux I__12596 (
            .O(N__56793),
            .I(N__56773));
    LocalMux I__12595 (
            .O(N__56788),
            .I(N__56773));
    InMux I__12594 (
            .O(N__56787),
            .I(N__56768));
    InMux I__12593 (
            .O(N__56784),
            .I(N__56768));
    Odrv4 I__12592 (
            .O(N__56781),
            .I(\ALU.N_125 ));
    Odrv4 I__12591 (
            .O(N__56778),
            .I(\ALU.N_125 ));
    Odrv12 I__12590 (
            .O(N__56773),
            .I(\ALU.N_125 ));
    LocalMux I__12589 (
            .O(N__56768),
            .I(\ALU.N_125 ));
    InMux I__12588 (
            .O(N__56759),
            .I(N__56756));
    LocalMux I__12587 (
            .O(N__56756),
            .I(\ALU.aluOut_i_13 ));
    InMux I__12586 (
            .O(N__56753),
            .I(N__56750));
    LocalMux I__12585 (
            .O(N__56750),
            .I(N__56745));
    InMux I__12584 (
            .O(N__56749),
            .I(N__56742));
    CascadeMux I__12583 (
            .O(N__56748),
            .I(N__56738));
    Span4Mux_v I__12582 (
            .O(N__56745),
            .I(N__56734));
    LocalMux I__12581 (
            .O(N__56742),
            .I(N__56731));
    InMux I__12580 (
            .O(N__56741),
            .I(N__56728));
    InMux I__12579 (
            .O(N__56738),
            .I(N__56723));
    InMux I__12578 (
            .O(N__56737),
            .I(N__56723));
    Span4Mux_h I__12577 (
            .O(N__56734),
            .I(N__56720));
    Span4Mux_h I__12576 (
            .O(N__56731),
            .I(N__56713));
    LocalMux I__12575 (
            .O(N__56728),
            .I(N__56713));
    LocalMux I__12574 (
            .O(N__56723),
            .I(N__56710));
    Sp12to4 I__12573 (
            .O(N__56720),
            .I(N__56707));
    InMux I__12572 (
            .O(N__56719),
            .I(N__56702));
    InMux I__12571 (
            .O(N__56718),
            .I(N__56702));
    Span4Mux_v I__12570 (
            .O(N__56713),
            .I(N__56699));
    Span4Mux_h I__12569 (
            .O(N__56710),
            .I(N__56696));
    Span12Mux_v I__12568 (
            .O(N__56707),
            .I(N__56693));
    LocalMux I__12567 (
            .O(N__56702),
            .I(N__56688));
    Span4Mux_v I__12566 (
            .O(N__56699),
            .I(N__56688));
    Span4Mux_h I__12565 (
            .O(N__56696),
            .I(N__56685));
    Odrv12 I__12564 (
            .O(N__56693),
            .I(\ALU.status_19_13 ));
    Odrv4 I__12563 (
            .O(N__56688),
            .I(\ALU.status_19_13 ));
    Odrv4 I__12562 (
            .O(N__56685),
            .I(\ALU.status_19_13 ));
    CascadeMux I__12561 (
            .O(N__56678),
            .I(N__56675));
    InMux I__12560 (
            .O(N__56675),
            .I(N__56672));
    LocalMux I__12559 (
            .O(N__56672),
            .I(\ALU.aluOut_i_14 ));
    CascadeMux I__12558 (
            .O(N__56669),
            .I(N__56666));
    InMux I__12557 (
            .O(N__56666),
            .I(N__56663));
    LocalMux I__12556 (
            .O(N__56663),
            .I(\ALU.aluOut_i_15 ));
    InMux I__12555 (
            .O(N__56660),
            .I(bfn_23_9_0_));
    InMux I__12554 (
            .O(N__56657),
            .I(N__56651));
    InMux I__12553 (
            .O(N__56656),
            .I(N__56651));
    LocalMux I__12552 (
            .O(N__56651),
            .I(N__56648));
    Span4Mux_v I__12551 (
            .O(N__56648),
            .I(N__56644));
    CascadeMux I__12550 (
            .O(N__56647),
            .I(N__56641));
    Span4Mux_h I__12549 (
            .O(N__56644),
            .I(N__56638));
    InMux I__12548 (
            .O(N__56641),
            .I(N__56635));
    Sp12to4 I__12547 (
            .O(N__56638),
            .I(N__56632));
    LocalMux I__12546 (
            .O(N__56635),
            .I(aluStatus_5));
    Odrv12 I__12545 (
            .O(N__56632),
            .I(aluStatus_5));
    CascadeMux I__12544 (
            .O(N__56627),
            .I(N__56624));
    InMux I__12543 (
            .O(N__56624),
            .I(N__56618));
    CascadeMux I__12542 (
            .O(N__56623),
            .I(N__56615));
    InMux I__12541 (
            .O(N__56622),
            .I(N__56610));
    InMux I__12540 (
            .O(N__56621),
            .I(N__56610));
    LocalMux I__12539 (
            .O(N__56618),
            .I(N__56607));
    InMux I__12538 (
            .O(N__56615),
            .I(N__56604));
    LocalMux I__12537 (
            .O(N__56610),
            .I(N__56600));
    Span4Mux_h I__12536 (
            .O(N__56607),
            .I(N__56595));
    LocalMux I__12535 (
            .O(N__56604),
            .I(N__56595));
    CEMux I__12534 (
            .O(N__56603),
            .I(N__56592));
    Span4Mux_h I__12533 (
            .O(N__56600),
            .I(N__56589));
    Span4Mux_v I__12532 (
            .O(N__56595),
            .I(N__56586));
    LocalMux I__12531 (
            .O(N__56592),
            .I(N__56583));
    Span4Mux_h I__12530 (
            .O(N__56589),
            .I(N__56580));
    Span4Mux_v I__12529 (
            .O(N__56586),
            .I(N__56577));
    Span4Mux_v I__12528 (
            .O(N__56583),
            .I(N__56574));
    Sp12to4 I__12527 (
            .O(N__56580),
            .I(N__56570));
    Span4Mux_h I__12526 (
            .O(N__56577),
            .I(N__56567));
    Span4Mux_v I__12525 (
            .O(N__56574),
            .I(N__56564));
    InMux I__12524 (
            .O(N__56573),
            .I(N__56561));
    Span12Mux_s8_v I__12523 (
            .O(N__56570),
            .I(N__56558));
    Span4Mux_h I__12522 (
            .O(N__56567),
            .I(N__56555));
    Span4Mux_h I__12521 (
            .O(N__56564),
            .I(N__56552));
    LocalMux I__12520 (
            .O(N__56561),
            .I(\ALU.un1_a41_0 ));
    Odrv12 I__12519 (
            .O(N__56558),
            .I(\ALU.un1_a41_0 ));
    Odrv4 I__12518 (
            .O(N__56555),
            .I(\ALU.un1_a41_0 ));
    Odrv4 I__12517 (
            .O(N__56552),
            .I(\ALU.un1_a41_0 ));
    InMux I__12516 (
            .O(N__56543),
            .I(N__56539));
    CascadeMux I__12515 (
            .O(N__56542),
            .I(N__56536));
    LocalMux I__12514 (
            .O(N__56539),
            .I(N__56533));
    InMux I__12513 (
            .O(N__56536),
            .I(N__56529));
    Span4Mux_h I__12512 (
            .O(N__56533),
            .I(N__56526));
    InMux I__12511 (
            .O(N__56532),
            .I(N__56523));
    LocalMux I__12510 (
            .O(N__56529),
            .I(N__56520));
    Span4Mux_h I__12509 (
            .O(N__56526),
            .I(N__56517));
    LocalMux I__12508 (
            .O(N__56523),
            .I(N__56514));
    Span4Mux_v I__12507 (
            .O(N__56520),
            .I(N__56511));
    Span4Mux_v I__12506 (
            .O(N__56517),
            .I(N__56506));
    Span4Mux_v I__12505 (
            .O(N__56514),
            .I(N__56506));
    Sp12to4 I__12504 (
            .O(N__56511),
            .I(N__56503));
    Sp12to4 I__12503 (
            .O(N__56506),
            .I(N__56500));
    Span12Mux_h I__12502 (
            .O(N__56503),
            .I(N__56495));
    Span12Mux_h I__12501 (
            .O(N__56500),
            .I(N__56495));
    Odrv12 I__12500 (
            .O(N__56495),
            .I(\ALU.aZ0Z32 ));
    InMux I__12499 (
            .O(N__56492),
            .I(N__56487));
    InMux I__12498 (
            .O(N__56491),
            .I(N__56482));
    InMux I__12497 (
            .O(N__56490),
            .I(N__56482));
    LocalMux I__12496 (
            .O(N__56487),
            .I(N__56479));
    LocalMux I__12495 (
            .O(N__56482),
            .I(\ALU.N_866 ));
    Odrv12 I__12494 (
            .O(N__56479),
            .I(\ALU.N_866 ));
    InMux I__12493 (
            .O(N__56474),
            .I(N__56469));
    InMux I__12492 (
            .O(N__56473),
            .I(N__56466));
    CascadeMux I__12491 (
            .O(N__56472),
            .I(N__56462));
    LocalMux I__12490 (
            .O(N__56469),
            .I(N__56459));
    LocalMux I__12489 (
            .O(N__56466),
            .I(N__56456));
    InMux I__12488 (
            .O(N__56465),
            .I(N__56453));
    InMux I__12487 (
            .O(N__56462),
            .I(N__56450));
    Span4Mux_h I__12486 (
            .O(N__56459),
            .I(N__56445));
    Span4Mux_h I__12485 (
            .O(N__56456),
            .I(N__56445));
    LocalMux I__12484 (
            .O(N__56453),
            .I(N__56442));
    LocalMux I__12483 (
            .O(N__56450),
            .I(N__56439));
    Sp12to4 I__12482 (
            .O(N__56445),
            .I(N__56434));
    Span12Mux_h I__12481 (
            .O(N__56442),
            .I(N__56434));
    Span4Mux_h I__12480 (
            .O(N__56439),
            .I(N__56431));
    Odrv12 I__12479 (
            .O(N__56434),
            .I(\ALU.N_967 ));
    Odrv4 I__12478 (
            .O(N__56431),
            .I(\ALU.N_967 ));
    CascadeMux I__12477 (
            .O(N__56426),
            .I(N__56423));
    InMux I__12476 (
            .O(N__56423),
            .I(N__56420));
    LocalMux I__12475 (
            .O(N__56420),
            .I(\ALU.aluOut_i_3 ));
    InMux I__12474 (
            .O(N__56417),
            .I(N__56410));
    InMux I__12473 (
            .O(N__56416),
            .I(N__56407));
    InMux I__12472 (
            .O(N__56415),
            .I(N__56402));
    InMux I__12471 (
            .O(N__56414),
            .I(N__56402));
    InMux I__12470 (
            .O(N__56413),
            .I(N__56398));
    LocalMux I__12469 (
            .O(N__56410),
            .I(N__56395));
    LocalMux I__12468 (
            .O(N__56407),
            .I(N__56391));
    LocalMux I__12467 (
            .O(N__56402),
            .I(N__56388));
    InMux I__12466 (
            .O(N__56401),
            .I(N__56385));
    LocalMux I__12465 (
            .O(N__56398),
            .I(N__56382));
    Span4Mux_v I__12464 (
            .O(N__56395),
            .I(N__56379));
    InMux I__12463 (
            .O(N__56394),
            .I(N__56374));
    Span4Mux_h I__12462 (
            .O(N__56391),
            .I(N__56371));
    Span4Mux_h I__12461 (
            .O(N__56388),
            .I(N__56366));
    LocalMux I__12460 (
            .O(N__56385),
            .I(N__56366));
    Span4Mux_v I__12459 (
            .O(N__56382),
            .I(N__56361));
    Span4Mux_h I__12458 (
            .O(N__56379),
            .I(N__56361));
    InMux I__12457 (
            .O(N__56378),
            .I(N__56352));
    InMux I__12456 (
            .O(N__56377),
            .I(N__56352));
    LocalMux I__12455 (
            .O(N__56374),
            .I(N__56347));
    Span4Mux_h I__12454 (
            .O(N__56371),
            .I(N__56347));
    Span4Mux_h I__12453 (
            .O(N__56366),
            .I(N__56342));
    Span4Mux_h I__12452 (
            .O(N__56361),
            .I(N__56339));
    InMux I__12451 (
            .O(N__56360),
            .I(N__56336));
    InMux I__12450 (
            .O(N__56359),
            .I(N__56329));
    InMux I__12449 (
            .O(N__56358),
            .I(N__56329));
    InMux I__12448 (
            .O(N__56357),
            .I(N__56329));
    LocalMux I__12447 (
            .O(N__56352),
            .I(N__56321));
    Span4Mux_h I__12446 (
            .O(N__56347),
            .I(N__56321));
    InMux I__12445 (
            .O(N__56346),
            .I(N__56316));
    InMux I__12444 (
            .O(N__56345),
            .I(N__56316));
    Span4Mux_v I__12443 (
            .O(N__56342),
            .I(N__56313));
    Span4Mux_h I__12442 (
            .O(N__56339),
            .I(N__56306));
    LocalMux I__12441 (
            .O(N__56336),
            .I(N__56306));
    LocalMux I__12440 (
            .O(N__56329),
            .I(N__56306));
    InMux I__12439 (
            .O(N__56328),
            .I(N__56303));
    InMux I__12438 (
            .O(N__56327),
            .I(N__56298));
    InMux I__12437 (
            .O(N__56326),
            .I(N__56298));
    Odrv4 I__12436 (
            .O(N__56321),
            .I(\ALU.status_19_3 ));
    LocalMux I__12435 (
            .O(N__56316),
            .I(\ALU.status_19_3 ));
    Odrv4 I__12434 (
            .O(N__56313),
            .I(\ALU.status_19_3 ));
    Odrv4 I__12433 (
            .O(N__56306),
            .I(\ALU.status_19_3 ));
    LocalMux I__12432 (
            .O(N__56303),
            .I(\ALU.status_19_3 ));
    LocalMux I__12431 (
            .O(N__56298),
            .I(\ALU.status_19_3 ));
    CascadeMux I__12430 (
            .O(N__56285),
            .I(N__56282));
    InMux I__12429 (
            .O(N__56282),
            .I(N__56279));
    LocalMux I__12428 (
            .O(N__56279),
            .I(\ALU.aluOut_i_4 ));
    InMux I__12427 (
            .O(N__56276),
            .I(N__56273));
    LocalMux I__12426 (
            .O(N__56273),
            .I(N__56269));
    CascadeMux I__12425 (
            .O(N__56272),
            .I(N__56263));
    Span4Mux_h I__12424 (
            .O(N__56269),
            .I(N__56260));
    CascadeMux I__12423 (
            .O(N__56268),
            .I(N__56256));
    InMux I__12422 (
            .O(N__56267),
            .I(N__56253));
    InMux I__12421 (
            .O(N__56266),
            .I(N__56250));
    InMux I__12420 (
            .O(N__56263),
            .I(N__56247));
    Span4Mux_v I__12419 (
            .O(N__56260),
            .I(N__56244));
    InMux I__12418 (
            .O(N__56259),
            .I(N__56241));
    InMux I__12417 (
            .O(N__56256),
            .I(N__56236));
    LocalMux I__12416 (
            .O(N__56253),
            .I(N__56233));
    LocalMux I__12415 (
            .O(N__56250),
            .I(N__56230));
    LocalMux I__12414 (
            .O(N__56247),
            .I(N__56225));
    Sp12to4 I__12413 (
            .O(N__56244),
            .I(N__56218));
    LocalMux I__12412 (
            .O(N__56241),
            .I(N__56218));
    InMux I__12411 (
            .O(N__56240),
            .I(N__56213));
    InMux I__12410 (
            .O(N__56239),
            .I(N__56213));
    LocalMux I__12409 (
            .O(N__56236),
            .I(N__56206));
    Span4Mux_v I__12408 (
            .O(N__56233),
            .I(N__56206));
    Span4Mux_h I__12407 (
            .O(N__56230),
            .I(N__56206));
    CascadeMux I__12406 (
            .O(N__56229),
            .I(N__56203));
    CascadeMux I__12405 (
            .O(N__56228),
            .I(N__56197));
    Span4Mux_v I__12404 (
            .O(N__56225),
            .I(N__56193));
    InMux I__12403 (
            .O(N__56224),
            .I(N__56188));
    InMux I__12402 (
            .O(N__56223),
            .I(N__56188));
    Span12Mux_h I__12401 (
            .O(N__56218),
            .I(N__56185));
    LocalMux I__12400 (
            .O(N__56213),
            .I(N__56182));
    Span4Mux_h I__12399 (
            .O(N__56206),
            .I(N__56179));
    InMux I__12398 (
            .O(N__56203),
            .I(N__56168));
    InMux I__12397 (
            .O(N__56202),
            .I(N__56168));
    InMux I__12396 (
            .O(N__56201),
            .I(N__56168));
    InMux I__12395 (
            .O(N__56200),
            .I(N__56168));
    InMux I__12394 (
            .O(N__56197),
            .I(N__56168));
    InMux I__12393 (
            .O(N__56196),
            .I(N__56165));
    Odrv4 I__12392 (
            .O(N__56193),
            .I(\ALU.status_19_4 ));
    LocalMux I__12391 (
            .O(N__56188),
            .I(\ALU.status_19_4 ));
    Odrv12 I__12390 (
            .O(N__56185),
            .I(\ALU.status_19_4 ));
    Odrv4 I__12389 (
            .O(N__56182),
            .I(\ALU.status_19_4 ));
    Odrv4 I__12388 (
            .O(N__56179),
            .I(\ALU.status_19_4 ));
    LocalMux I__12387 (
            .O(N__56168),
            .I(\ALU.status_19_4 ));
    LocalMux I__12386 (
            .O(N__56165),
            .I(\ALU.status_19_4 ));
    CascadeMux I__12385 (
            .O(N__56150),
            .I(N__56147));
    InMux I__12384 (
            .O(N__56147),
            .I(N__56144));
    LocalMux I__12383 (
            .O(N__56144),
            .I(\ALU.aluOut_i_5 ));
    CascadeMux I__12382 (
            .O(N__56141),
            .I(N__56138));
    InMux I__12381 (
            .O(N__56138),
            .I(N__56135));
    LocalMux I__12380 (
            .O(N__56135),
            .I(N__56132));
    Span4Mux_v I__12379 (
            .O(N__56132),
            .I(N__56127));
    InMux I__12378 (
            .O(N__56131),
            .I(N__56124));
    CascadeMux I__12377 (
            .O(N__56130),
            .I(N__56121));
    Span4Mux_v I__12376 (
            .O(N__56127),
            .I(N__56117));
    LocalMux I__12375 (
            .O(N__56124),
            .I(N__56112));
    InMux I__12374 (
            .O(N__56121),
            .I(N__56109));
    InMux I__12373 (
            .O(N__56120),
            .I(N__56106));
    Span4Mux_h I__12372 (
            .O(N__56117),
            .I(N__56103));
    InMux I__12371 (
            .O(N__56116),
            .I(N__56100));
    InMux I__12370 (
            .O(N__56115),
            .I(N__56097));
    Span4Mux_v I__12369 (
            .O(N__56112),
            .I(N__56093));
    LocalMux I__12368 (
            .O(N__56109),
            .I(N__56090));
    LocalMux I__12367 (
            .O(N__56106),
            .I(N__56087));
    Span4Mux_h I__12366 (
            .O(N__56103),
            .I(N__56083));
    LocalMux I__12365 (
            .O(N__56100),
            .I(N__56079));
    LocalMux I__12364 (
            .O(N__56097),
            .I(N__56073));
    CascadeMux I__12363 (
            .O(N__56096),
            .I(N__56070));
    Span4Mux_v I__12362 (
            .O(N__56093),
            .I(N__56065));
    Span4Mux_v I__12361 (
            .O(N__56090),
            .I(N__56060));
    Span4Mux_v I__12360 (
            .O(N__56087),
            .I(N__56060));
    InMux I__12359 (
            .O(N__56086),
            .I(N__56057));
    Span4Mux_v I__12358 (
            .O(N__56083),
            .I(N__56054));
    InMux I__12357 (
            .O(N__56082),
            .I(N__56051));
    Span4Mux_v I__12356 (
            .O(N__56079),
            .I(N__56048));
    InMux I__12355 (
            .O(N__56078),
            .I(N__56043));
    InMux I__12354 (
            .O(N__56077),
            .I(N__56043));
    InMux I__12353 (
            .O(N__56076),
            .I(N__56040));
    Span4Mux_h I__12352 (
            .O(N__56073),
            .I(N__56037));
    InMux I__12351 (
            .O(N__56070),
            .I(N__56032));
    InMux I__12350 (
            .O(N__56069),
            .I(N__56032));
    InMux I__12349 (
            .O(N__56068),
            .I(N__56029));
    Sp12to4 I__12348 (
            .O(N__56065),
            .I(N__56022));
    Sp12to4 I__12347 (
            .O(N__56060),
            .I(N__56022));
    LocalMux I__12346 (
            .O(N__56057),
            .I(N__56022));
    Odrv4 I__12345 (
            .O(N__56054),
            .I(\ALU.status_19_5 ));
    LocalMux I__12344 (
            .O(N__56051),
            .I(\ALU.status_19_5 ));
    Odrv4 I__12343 (
            .O(N__56048),
            .I(\ALU.status_19_5 ));
    LocalMux I__12342 (
            .O(N__56043),
            .I(\ALU.status_19_5 ));
    LocalMux I__12341 (
            .O(N__56040),
            .I(\ALU.status_19_5 ));
    Odrv4 I__12340 (
            .O(N__56037),
            .I(\ALU.status_19_5 ));
    LocalMux I__12339 (
            .O(N__56032),
            .I(\ALU.status_19_5 ));
    LocalMux I__12338 (
            .O(N__56029),
            .I(\ALU.status_19_5 ));
    Odrv12 I__12337 (
            .O(N__56022),
            .I(\ALU.status_19_5 ));
    CascadeMux I__12336 (
            .O(N__56003),
            .I(N__56000));
    InMux I__12335 (
            .O(N__56000),
            .I(N__55997));
    LocalMux I__12334 (
            .O(N__55997),
            .I(\ALU.aluOut_i_6 ));
    InMux I__12333 (
            .O(N__55994),
            .I(N__55986));
    InMux I__12332 (
            .O(N__55993),
            .I(N__55979));
    InMux I__12331 (
            .O(N__55992),
            .I(N__55979));
    InMux I__12330 (
            .O(N__55991),
            .I(N__55976));
    CascadeMux I__12329 (
            .O(N__55990),
            .I(N__55973));
    InMux I__12328 (
            .O(N__55989),
            .I(N__55970));
    LocalMux I__12327 (
            .O(N__55986),
            .I(N__55967));
    InMux I__12326 (
            .O(N__55985),
            .I(N__55964));
    CascadeMux I__12325 (
            .O(N__55984),
            .I(N__55961));
    LocalMux I__12324 (
            .O(N__55979),
            .I(N__55954));
    LocalMux I__12323 (
            .O(N__55976),
            .I(N__55950));
    InMux I__12322 (
            .O(N__55973),
            .I(N__55946));
    LocalMux I__12321 (
            .O(N__55970),
            .I(N__55941));
    Span4Mux_v I__12320 (
            .O(N__55967),
            .I(N__55941));
    LocalMux I__12319 (
            .O(N__55964),
            .I(N__55938));
    InMux I__12318 (
            .O(N__55961),
            .I(N__55931));
    InMux I__12317 (
            .O(N__55960),
            .I(N__55931));
    InMux I__12316 (
            .O(N__55959),
            .I(N__55931));
    InMux I__12315 (
            .O(N__55958),
            .I(N__55928));
    InMux I__12314 (
            .O(N__55957),
            .I(N__55925));
    Span4Mux_h I__12313 (
            .O(N__55954),
            .I(N__55922));
    InMux I__12312 (
            .O(N__55953),
            .I(N__55919));
    Span4Mux_v I__12311 (
            .O(N__55950),
            .I(N__55916));
    InMux I__12310 (
            .O(N__55949),
            .I(N__55913));
    LocalMux I__12309 (
            .O(N__55946),
            .I(N__55904));
    Span4Mux_h I__12308 (
            .O(N__55941),
            .I(N__55904));
    Span4Mux_v I__12307 (
            .O(N__55938),
            .I(N__55904));
    LocalMux I__12306 (
            .O(N__55931),
            .I(N__55904));
    LocalMux I__12305 (
            .O(N__55928),
            .I(N__55901));
    LocalMux I__12304 (
            .O(N__55925),
            .I(N__55898));
    Span4Mux_h I__12303 (
            .O(N__55922),
            .I(N__55893));
    LocalMux I__12302 (
            .O(N__55919),
            .I(N__55893));
    Span4Mux_h I__12301 (
            .O(N__55916),
            .I(N__55888));
    LocalMux I__12300 (
            .O(N__55913),
            .I(N__55888));
    Span4Mux_h I__12299 (
            .O(N__55904),
            .I(N__55882));
    Span4Mux_v I__12298 (
            .O(N__55901),
            .I(N__55879));
    Span4Mux_v I__12297 (
            .O(N__55898),
            .I(N__55876));
    Span4Mux_h I__12296 (
            .O(N__55893),
            .I(N__55872));
    Span4Mux_v I__12295 (
            .O(N__55888),
            .I(N__55869));
    InMux I__12294 (
            .O(N__55887),
            .I(N__55862));
    InMux I__12293 (
            .O(N__55886),
            .I(N__55862));
    InMux I__12292 (
            .O(N__55885),
            .I(N__55862));
    Span4Mux_h I__12291 (
            .O(N__55882),
            .I(N__55859));
    Span4Mux_v I__12290 (
            .O(N__55879),
            .I(N__55854));
    Span4Mux_h I__12289 (
            .O(N__55876),
            .I(N__55854));
    InMux I__12288 (
            .O(N__55875),
            .I(N__55851));
    Span4Mux_v I__12287 (
            .O(N__55872),
            .I(N__55848));
    Odrv4 I__12286 (
            .O(N__55869),
            .I(\ALU.status_19_6 ));
    LocalMux I__12285 (
            .O(N__55862),
            .I(\ALU.status_19_6 ));
    Odrv4 I__12284 (
            .O(N__55859),
            .I(\ALU.status_19_6 ));
    Odrv4 I__12283 (
            .O(N__55854),
            .I(\ALU.status_19_6 ));
    LocalMux I__12282 (
            .O(N__55851),
            .I(\ALU.status_19_6 ));
    Odrv4 I__12281 (
            .O(N__55848),
            .I(\ALU.status_19_6 ));
    CascadeMux I__12280 (
            .O(N__55835),
            .I(N__55832));
    InMux I__12279 (
            .O(N__55832),
            .I(N__55829));
    LocalMux I__12278 (
            .O(N__55829),
            .I(N__55826));
    Odrv4 I__12277 (
            .O(N__55826),
            .I(\ALU.aluOut_i_7 ));
    CascadeMux I__12276 (
            .O(N__55823),
            .I(N__55818));
    InMux I__12275 (
            .O(N__55822),
            .I(N__55813));
    InMux I__12274 (
            .O(N__55821),
            .I(N__55808));
    InMux I__12273 (
            .O(N__55818),
            .I(N__55805));
    InMux I__12272 (
            .O(N__55817),
            .I(N__55802));
    CascadeMux I__12271 (
            .O(N__55816),
            .I(N__55796));
    LocalMux I__12270 (
            .O(N__55813),
            .I(N__55793));
    InMux I__12269 (
            .O(N__55812),
            .I(N__55788));
    InMux I__12268 (
            .O(N__55811),
            .I(N__55788));
    LocalMux I__12267 (
            .O(N__55808),
            .I(N__55783));
    LocalMux I__12266 (
            .O(N__55805),
            .I(N__55783));
    LocalMux I__12265 (
            .O(N__55802),
            .I(N__55780));
    InMux I__12264 (
            .O(N__55801),
            .I(N__55777));
    InMux I__12263 (
            .O(N__55800),
            .I(N__55772));
    InMux I__12262 (
            .O(N__55799),
            .I(N__55772));
    InMux I__12261 (
            .O(N__55796),
            .I(N__55769));
    Span4Mux_v I__12260 (
            .O(N__55793),
            .I(N__55764));
    LocalMux I__12259 (
            .O(N__55788),
            .I(N__55761));
    Span4Mux_v I__12258 (
            .O(N__55783),
            .I(N__55752));
    Span4Mux_v I__12257 (
            .O(N__55780),
            .I(N__55752));
    LocalMux I__12256 (
            .O(N__55777),
            .I(N__55752));
    LocalMux I__12255 (
            .O(N__55772),
            .I(N__55752));
    LocalMux I__12254 (
            .O(N__55769),
            .I(N__55749));
    InMux I__12253 (
            .O(N__55768),
            .I(N__55746));
    InMux I__12252 (
            .O(N__55767),
            .I(N__55743));
    Sp12to4 I__12251 (
            .O(N__55764),
            .I(N__55740));
    Span4Mux_h I__12250 (
            .O(N__55761),
            .I(N__55737));
    Span4Mux_h I__12249 (
            .O(N__55752),
            .I(N__55734));
    Span4Mux_h I__12248 (
            .O(N__55749),
            .I(N__55727));
    LocalMux I__12247 (
            .O(N__55746),
            .I(N__55727));
    LocalMux I__12246 (
            .O(N__55743),
            .I(N__55727));
    Span12Mux_h I__12245 (
            .O(N__55740),
            .I(N__55721));
    Span4Mux_v I__12244 (
            .O(N__55737),
            .I(N__55716));
    Span4Mux_v I__12243 (
            .O(N__55734),
            .I(N__55716));
    Span4Mux_v I__12242 (
            .O(N__55727),
            .I(N__55713));
    InMux I__12241 (
            .O(N__55726),
            .I(N__55706));
    InMux I__12240 (
            .O(N__55725),
            .I(N__55706));
    InMux I__12239 (
            .O(N__55724),
            .I(N__55706));
    Odrv12 I__12238 (
            .O(N__55721),
            .I(\ALU.status_19_7 ));
    Odrv4 I__12237 (
            .O(N__55716),
            .I(\ALU.status_19_7 ));
    Odrv4 I__12236 (
            .O(N__55713),
            .I(\ALU.status_19_7 ));
    LocalMux I__12235 (
            .O(N__55706),
            .I(\ALU.status_19_7 ));
    CascadeMux I__12234 (
            .O(N__55697),
            .I(N__55694));
    InMux I__12233 (
            .O(N__55694),
            .I(N__55691));
    LocalMux I__12232 (
            .O(N__55691),
            .I(\ALU.aluOut_i_8 ));
    CascadeMux I__12231 (
            .O(N__55688),
            .I(N__55682));
    InMux I__12230 (
            .O(N__55687),
            .I(N__55678));
    CascadeMux I__12229 (
            .O(N__55686),
            .I(N__55675));
    CascadeMux I__12228 (
            .O(N__55685),
            .I(N__55671));
    InMux I__12227 (
            .O(N__55682),
            .I(N__55665));
    InMux I__12226 (
            .O(N__55681),
            .I(N__55665));
    LocalMux I__12225 (
            .O(N__55678),
            .I(N__55662));
    InMux I__12224 (
            .O(N__55675),
            .I(N__55657));
    InMux I__12223 (
            .O(N__55674),
            .I(N__55654));
    InMux I__12222 (
            .O(N__55671),
            .I(N__55651));
    CascadeMux I__12221 (
            .O(N__55670),
            .I(N__55648));
    LocalMux I__12220 (
            .O(N__55665),
            .I(N__55644));
    Span12Mux_s8_v I__12219 (
            .O(N__55662),
            .I(N__55641));
    InMux I__12218 (
            .O(N__55661),
            .I(N__55638));
    InMux I__12217 (
            .O(N__55660),
            .I(N__55635));
    LocalMux I__12216 (
            .O(N__55657),
            .I(N__55628));
    LocalMux I__12215 (
            .O(N__55654),
            .I(N__55628));
    LocalMux I__12214 (
            .O(N__55651),
            .I(N__55628));
    InMux I__12213 (
            .O(N__55648),
            .I(N__55625));
    InMux I__12212 (
            .O(N__55647),
            .I(N__55622));
    Span4Mux_v I__12211 (
            .O(N__55644),
            .I(N__55619));
    Span12Mux_h I__12210 (
            .O(N__55641),
            .I(N__55612));
    LocalMux I__12209 (
            .O(N__55638),
            .I(N__55612));
    LocalMux I__12208 (
            .O(N__55635),
            .I(N__55612));
    Span4Mux_h I__12207 (
            .O(N__55628),
            .I(N__55609));
    LocalMux I__12206 (
            .O(N__55625),
            .I(\ALU.status_19_8 ));
    LocalMux I__12205 (
            .O(N__55622),
            .I(\ALU.status_19_8 ));
    Odrv4 I__12204 (
            .O(N__55619),
            .I(\ALU.status_19_8 ));
    Odrv12 I__12203 (
            .O(N__55612),
            .I(\ALU.status_19_8 ));
    Odrv4 I__12202 (
            .O(N__55609),
            .I(\ALU.status_19_8 ));
    CascadeMux I__12201 (
            .O(N__55598),
            .I(N__55595));
    InMux I__12200 (
            .O(N__55595),
            .I(N__55592));
    LocalMux I__12199 (
            .O(N__55592),
            .I(\ALU.aluOut_i_9 ));
    InMux I__12198 (
            .O(N__55589),
            .I(N__55586));
    LocalMux I__12197 (
            .O(N__55586),
            .I(N__55582));
    InMux I__12196 (
            .O(N__55585),
            .I(N__55579));
    Span4Mux_v I__12195 (
            .O(N__55582),
            .I(N__55573));
    LocalMux I__12194 (
            .O(N__55579),
            .I(N__55570));
    InMux I__12193 (
            .O(N__55578),
            .I(N__55565));
    InMux I__12192 (
            .O(N__55577),
            .I(N__55565));
    InMux I__12191 (
            .O(N__55576),
            .I(N__55562));
    Sp12to4 I__12190 (
            .O(N__55573),
            .I(N__55559));
    Span4Mux_h I__12189 (
            .O(N__55570),
            .I(N__55555));
    LocalMux I__12188 (
            .O(N__55565),
            .I(N__55550));
    LocalMux I__12187 (
            .O(N__55562),
            .I(N__55550));
    Span12Mux_h I__12186 (
            .O(N__55559),
            .I(N__55543));
    InMux I__12185 (
            .O(N__55558),
            .I(N__55540));
    Span4Mux_v I__12184 (
            .O(N__55555),
            .I(N__55535));
    Span4Mux_h I__12183 (
            .O(N__55550),
            .I(N__55535));
    InMux I__12182 (
            .O(N__55549),
            .I(N__55526));
    InMux I__12181 (
            .O(N__55548),
            .I(N__55526));
    InMux I__12180 (
            .O(N__55547),
            .I(N__55526));
    InMux I__12179 (
            .O(N__55546),
            .I(N__55526));
    Odrv12 I__12178 (
            .O(N__55543),
            .I(\ALU.status_19_9 ));
    LocalMux I__12177 (
            .O(N__55540),
            .I(\ALU.status_19_9 ));
    Odrv4 I__12176 (
            .O(N__55535),
            .I(\ALU.status_19_9 ));
    LocalMux I__12175 (
            .O(N__55526),
            .I(\ALU.status_19_9 ));
    CascadeMux I__12174 (
            .O(N__55517),
            .I(N__55514));
    InMux I__12173 (
            .O(N__55514),
            .I(N__55511));
    LocalMux I__12172 (
            .O(N__55511),
            .I(N__55508));
    Odrv4 I__12171 (
            .O(N__55508),
            .I(\ALU.aluOut_i_10 ));
    CascadeMux I__12170 (
            .O(N__55505),
            .I(N__55502));
    InMux I__12169 (
            .O(N__55502),
            .I(N__55499));
    LocalMux I__12168 (
            .O(N__55499),
            .I(N__55496));
    Span4Mux_v I__12167 (
            .O(N__55496),
            .I(N__55493));
    Sp12to4 I__12166 (
            .O(N__55493),
            .I(N__55490));
    Span12Mux_h I__12165 (
            .O(N__55490),
            .I(N__55487));
    Odrv12 I__12164 (
            .O(N__55487),
            .I(\PROM.ROMDATA.m158 ));
    CascadeMux I__12163 (
            .O(N__55484),
            .I(\PROM.ROMDATA.m158_cascade_ ));
    InMux I__12162 (
            .O(N__55481),
            .I(N__55478));
    LocalMux I__12161 (
            .O(N__55478),
            .I(\PROM.ROMDATA.m196_ns ));
    InMux I__12160 (
            .O(N__55475),
            .I(N__55467));
    InMux I__12159 (
            .O(N__55474),
            .I(N__55462));
    InMux I__12158 (
            .O(N__55473),
            .I(N__55457));
    InMux I__12157 (
            .O(N__55472),
            .I(N__55457));
    InMux I__12156 (
            .O(N__55471),
            .I(N__55448));
    InMux I__12155 (
            .O(N__55470),
            .I(N__55445));
    LocalMux I__12154 (
            .O(N__55467),
            .I(N__55441));
    InMux I__12153 (
            .O(N__55466),
            .I(N__55436));
    InMux I__12152 (
            .O(N__55465),
            .I(N__55436));
    LocalMux I__12151 (
            .O(N__55462),
            .I(N__55431));
    LocalMux I__12150 (
            .O(N__55457),
            .I(N__55431));
    InMux I__12149 (
            .O(N__55456),
            .I(N__55424));
    InMux I__12148 (
            .O(N__55455),
            .I(N__55424));
    InMux I__12147 (
            .O(N__55454),
            .I(N__55424));
    InMux I__12146 (
            .O(N__55453),
            .I(N__55418));
    InMux I__12145 (
            .O(N__55452),
            .I(N__55413));
    InMux I__12144 (
            .O(N__55451),
            .I(N__55413));
    LocalMux I__12143 (
            .O(N__55448),
            .I(N__55408));
    LocalMux I__12142 (
            .O(N__55445),
            .I(N__55408));
    InMux I__12141 (
            .O(N__55444),
            .I(N__55405));
    Span4Mux_v I__12140 (
            .O(N__55441),
            .I(N__55400));
    LocalMux I__12139 (
            .O(N__55436),
            .I(N__55400));
    Span4Mux_h I__12138 (
            .O(N__55431),
            .I(N__55396));
    LocalMux I__12137 (
            .O(N__55424),
            .I(N__55393));
    InMux I__12136 (
            .O(N__55423),
            .I(N__55386));
    InMux I__12135 (
            .O(N__55422),
            .I(N__55386));
    InMux I__12134 (
            .O(N__55421),
            .I(N__55386));
    LocalMux I__12133 (
            .O(N__55418),
            .I(N__55381));
    LocalMux I__12132 (
            .O(N__55413),
            .I(N__55381));
    Span4Mux_h I__12131 (
            .O(N__55408),
            .I(N__55376));
    LocalMux I__12130 (
            .O(N__55405),
            .I(N__55376));
    Span4Mux_h I__12129 (
            .O(N__55400),
            .I(N__55373));
    InMux I__12128 (
            .O(N__55399),
            .I(N__55370));
    Span4Mux_h I__12127 (
            .O(N__55396),
            .I(N__55365));
    Span4Mux_h I__12126 (
            .O(N__55393),
            .I(N__55365));
    LocalMux I__12125 (
            .O(N__55386),
            .I(N__55360));
    Span4Mux_v I__12124 (
            .O(N__55381),
            .I(N__55360));
    Span4Mux_h I__12123 (
            .O(N__55376),
            .I(N__55357));
    Span4Mux_h I__12122 (
            .O(N__55373),
            .I(N__55354));
    LocalMux I__12121 (
            .O(N__55370),
            .I(N__55351));
    Span4Mux_v I__12120 (
            .O(N__55365),
            .I(N__55346));
    Span4Mux_h I__12119 (
            .O(N__55360),
            .I(N__55346));
    Span4Mux_h I__12118 (
            .O(N__55357),
            .I(N__55343));
    Odrv4 I__12117 (
            .O(N__55354),
            .I(PROM_ROMDATA_dintern_6ro));
    Odrv12 I__12116 (
            .O(N__55351),
            .I(PROM_ROMDATA_dintern_6ro));
    Odrv4 I__12115 (
            .O(N__55346),
            .I(PROM_ROMDATA_dintern_6ro));
    Odrv4 I__12114 (
            .O(N__55343),
            .I(PROM_ROMDATA_dintern_6ro));
    InMux I__12113 (
            .O(N__55334),
            .I(N__55330));
    InMux I__12112 (
            .O(N__55333),
            .I(N__55327));
    LocalMux I__12111 (
            .O(N__55330),
            .I(N__55324));
    LocalMux I__12110 (
            .O(N__55327),
            .I(N__55321));
    Span4Mux_v I__12109 (
            .O(N__55324),
            .I(N__55318));
    Span12Mux_v I__12108 (
            .O(N__55321),
            .I(N__55315));
    Span4Mux_h I__12107 (
            .O(N__55318),
            .I(N__55312));
    Span12Mux_h I__12106 (
            .O(N__55315),
            .I(N__55309));
    Span4Mux_h I__12105 (
            .O(N__55312),
            .I(N__55306));
    Odrv12 I__12104 (
            .O(N__55309),
            .I(\CONTROL.ctrlOut_4 ));
    Odrv4 I__12103 (
            .O(N__55306),
            .I(\CONTROL.ctrlOut_4 ));
    InMux I__12102 (
            .O(N__55301),
            .I(N__55298));
    LocalMux I__12101 (
            .O(N__55298),
            .I(N__55295));
    Span4Mux_h I__12100 (
            .O(N__55295),
            .I(N__55291));
    InMux I__12099 (
            .O(N__55294),
            .I(N__55288));
    Odrv4 I__12098 (
            .O(N__55291),
            .I(\CONTROL.dout_reto_4 ));
    LocalMux I__12097 (
            .O(N__55288),
            .I(\CONTROL.dout_reto_4 ));
    CascadeMux I__12096 (
            .O(N__55283),
            .I(N__55280));
    InMux I__12095 (
            .O(N__55280),
            .I(N__55277));
    LocalMux I__12094 (
            .O(N__55277),
            .I(\ALU.aluOut_i_0 ));
    CascadeMux I__12093 (
            .O(N__55274),
            .I(N__55271));
    InMux I__12092 (
            .O(N__55271),
            .I(N__55268));
    LocalMux I__12091 (
            .O(N__55268),
            .I(\ALU.aluOut_i_1 ));
    CascadeMux I__12090 (
            .O(N__55265),
            .I(N__55262));
    InMux I__12089 (
            .O(N__55262),
            .I(N__55259));
    LocalMux I__12088 (
            .O(N__55259),
            .I(\ALU.aluOut_i_2 ));
    CascadeMux I__12087 (
            .O(N__55256),
            .I(\PROM.ROMDATA.m183_cascade_ ));
    InMux I__12086 (
            .O(N__55253),
            .I(N__55250));
    LocalMux I__12085 (
            .O(N__55250),
            .I(\PROM.ROMDATA.m185_bm ));
    CascadeMux I__12084 (
            .O(N__55247),
            .I(\PROM.ROMDATA.N_525_mux_cascade_ ));
    InMux I__12083 (
            .O(N__55244),
            .I(N__55241));
    LocalMux I__12082 (
            .O(N__55241),
            .I(\PROM.ROMDATA.i4_mux ));
    InMux I__12081 (
            .O(N__55238),
            .I(N__55235));
    LocalMux I__12080 (
            .O(N__55235),
            .I(N__55232));
    Span4Mux_h I__12079 (
            .O(N__55232),
            .I(N__55229));
    Odrv4 I__12078 (
            .O(N__55229),
            .I(\PROM.ROMDATA.m103 ));
    InMux I__12077 (
            .O(N__55226),
            .I(N__55223));
    LocalMux I__12076 (
            .O(N__55223),
            .I(N__55218));
    InMux I__12075 (
            .O(N__55222),
            .I(N__55215));
    InMux I__12074 (
            .O(N__55221),
            .I(N__55212));
    Odrv12 I__12073 (
            .O(N__55218),
            .I(\PROM.ROMDATA.m226 ));
    LocalMux I__12072 (
            .O(N__55215),
            .I(\PROM.ROMDATA.m226 ));
    LocalMux I__12071 (
            .O(N__55212),
            .I(\PROM.ROMDATA.m226 ));
    CascadeMux I__12070 (
            .O(N__55205),
            .I(N__55202));
    InMux I__12069 (
            .O(N__55202),
            .I(N__55199));
    LocalMux I__12068 (
            .O(N__55199),
            .I(\PROM.ROMDATA.m92_am_1 ));
    InMux I__12067 (
            .O(N__55196),
            .I(N__55193));
    LocalMux I__12066 (
            .O(N__55193),
            .I(N__55190));
    Span4Mux_h I__12065 (
            .O(N__55190),
            .I(N__55187));
    Odrv4 I__12064 (
            .O(N__55187),
            .I(\PROM.ROMDATA.m55 ));
    InMux I__12063 (
            .O(N__55184),
            .I(N__55180));
    InMux I__12062 (
            .O(N__55183),
            .I(N__55177));
    LocalMux I__12061 (
            .O(N__55180),
            .I(N__55174));
    LocalMux I__12060 (
            .O(N__55177),
            .I(\CONTROL.programCounter_1_reto_4 ));
    Odrv4 I__12059 (
            .O(N__55174),
            .I(\CONTROL.programCounter_1_reto_4 ));
    InMux I__12058 (
            .O(N__55169),
            .I(N__55164));
    InMux I__12057 (
            .O(N__55168),
            .I(N__55159));
    InMux I__12056 (
            .O(N__55167),
            .I(N__55159));
    LocalMux I__12055 (
            .O(N__55164),
            .I(N__55156));
    LocalMux I__12054 (
            .O(N__55159),
            .I(N__55152));
    Span4Mux_h I__12053 (
            .O(N__55156),
            .I(N__55149));
    InMux I__12052 (
            .O(N__55155),
            .I(N__55146));
    Odrv12 I__12051 (
            .O(N__55152),
            .I(CONTROL_addrstack_reto_4));
    Odrv4 I__12050 (
            .O(N__55149),
            .I(CONTROL_addrstack_reto_4));
    LocalMux I__12049 (
            .O(N__55146),
            .I(CONTROL_addrstack_reto_4));
    InMux I__12048 (
            .O(N__55139),
            .I(N__55134));
    InMux I__12047 (
            .O(N__55138),
            .I(N__55131));
    InMux I__12046 (
            .O(N__55137),
            .I(N__55128));
    LocalMux I__12045 (
            .O(N__55134),
            .I(N__55125));
    LocalMux I__12044 (
            .O(N__55131),
            .I(N__55115));
    LocalMux I__12043 (
            .O(N__55128),
            .I(N__55112));
    Span4Mux_h I__12042 (
            .O(N__55125),
            .I(N__55109));
    InMux I__12041 (
            .O(N__55124),
            .I(N__55104));
    InMux I__12040 (
            .O(N__55123),
            .I(N__55104));
    InMux I__12039 (
            .O(N__55122),
            .I(N__55099));
    InMux I__12038 (
            .O(N__55121),
            .I(N__55099));
    InMux I__12037 (
            .O(N__55120),
            .I(N__55092));
    InMux I__12036 (
            .O(N__55119),
            .I(N__55092));
    InMux I__12035 (
            .O(N__55118),
            .I(N__55092));
    Odrv4 I__12034 (
            .O(N__55115),
            .I(\CONTROL.programCounter11_reto_fast ));
    Odrv4 I__12033 (
            .O(N__55112),
            .I(\CONTROL.programCounter11_reto_fast ));
    Odrv4 I__12032 (
            .O(N__55109),
            .I(\CONTROL.programCounter11_reto_fast ));
    LocalMux I__12031 (
            .O(N__55104),
            .I(\CONTROL.programCounter11_reto_fast ));
    LocalMux I__12030 (
            .O(N__55099),
            .I(\CONTROL.programCounter11_reto_fast ));
    LocalMux I__12029 (
            .O(N__55092),
            .I(\CONTROL.programCounter11_reto_fast ));
    InMux I__12028 (
            .O(N__55079),
            .I(N__55074));
    InMux I__12027 (
            .O(N__55078),
            .I(N__55071));
    InMux I__12026 (
            .O(N__55077),
            .I(N__55068));
    LocalMux I__12025 (
            .O(N__55074),
            .I(N__55065));
    LocalMux I__12024 (
            .O(N__55071),
            .I(N__55059));
    LocalMux I__12023 (
            .O(N__55068),
            .I(N__55059));
    Span4Mux_v I__12022 (
            .O(N__55065),
            .I(N__55050));
    InMux I__12021 (
            .O(N__55064),
            .I(N__55047));
    Span4Mux_v I__12020 (
            .O(N__55059),
            .I(N__55044));
    InMux I__12019 (
            .O(N__55058),
            .I(N__55041));
    InMux I__12018 (
            .O(N__55057),
            .I(N__55036));
    InMux I__12017 (
            .O(N__55056),
            .I(N__55036));
    InMux I__12016 (
            .O(N__55055),
            .I(N__55033));
    InMux I__12015 (
            .O(N__55054),
            .I(N__55028));
    InMux I__12014 (
            .O(N__55053),
            .I(N__55028));
    Odrv4 I__12013 (
            .O(N__55050),
            .I(\CONTROL.un1_programCounter9_reto_fast ));
    LocalMux I__12012 (
            .O(N__55047),
            .I(\CONTROL.un1_programCounter9_reto_fast ));
    Odrv4 I__12011 (
            .O(N__55044),
            .I(\CONTROL.un1_programCounter9_reto_fast ));
    LocalMux I__12010 (
            .O(N__55041),
            .I(\CONTROL.un1_programCounter9_reto_fast ));
    LocalMux I__12009 (
            .O(N__55036),
            .I(\CONTROL.un1_programCounter9_reto_fast ));
    LocalMux I__12008 (
            .O(N__55033),
            .I(\CONTROL.un1_programCounter9_reto_fast ));
    LocalMux I__12007 (
            .O(N__55028),
            .I(\CONTROL.un1_programCounter9_reto_fast ));
    CascadeMux I__12006 (
            .O(N__55013),
            .I(\CONTROL.programCounter_ret_1_RNINC8IZ0Z_4_cascade_ ));
    InMux I__12005 (
            .O(N__55010),
            .I(N__55007));
    LocalMux I__12004 (
            .O(N__55007),
            .I(N__55004));
    Span4Mux_h I__12003 (
            .O(N__55004),
            .I(N__55001));
    Odrv4 I__12002 (
            .O(N__55001),
            .I(\CONTROL.programCounter_ret_19_RNIGQ8JZ0Z_4 ));
    InMux I__12001 (
            .O(N__54998),
            .I(N__54995));
    LocalMux I__12000 (
            .O(N__54995),
            .I(\PROM.ROMDATA.m143 ));
    CascadeMux I__11999 (
            .O(N__54992),
            .I(progRomAddress_4_cascade_));
    InMux I__11998 (
            .O(N__54989),
            .I(N__54986));
    LocalMux I__11997 (
            .O(N__54986),
            .I(N__54983));
    Odrv4 I__11996 (
            .O(N__54983),
            .I(\PROM.ROMDATA.m145 ));
    InMux I__11995 (
            .O(N__54980),
            .I(N__54977));
    LocalMux I__11994 (
            .O(N__54977),
            .I(N__54974));
    Span12Mux_s11_h I__11993 (
            .O(N__54974),
            .I(N__54971));
    Odrv12 I__11992 (
            .O(N__54971),
            .I(\PROM.ROMDATA.m90 ));
    InMux I__11991 (
            .O(N__54968),
            .I(N__54965));
    LocalMux I__11990 (
            .O(N__54965),
            .I(N__54962));
    Span4Mux_h I__11989 (
            .O(N__54962),
            .I(N__54959));
    Odrv4 I__11988 (
            .O(N__54959),
            .I(\PROM.ROMDATA.m92_bm ));
    InMux I__11987 (
            .O(N__54956),
            .I(N__54953));
    LocalMux I__11986 (
            .O(N__54953),
            .I(N__54950));
    Span4Mux_h I__11985 (
            .O(N__54950),
            .I(N__54947));
    Odrv4 I__11984 (
            .O(N__54947),
            .I(\PROM.ROMDATA.m11_am ));
    CascadeMux I__11983 (
            .O(N__54944),
            .I(\PROM.ROMDATA.m19_ns_1_cascade_ ));
    InMux I__11982 (
            .O(N__54941),
            .I(N__54938));
    LocalMux I__11981 (
            .O(N__54938),
            .I(\PROM.ROMDATA.m18_am ));
    InMux I__11980 (
            .O(N__54935),
            .I(N__54932));
    LocalMux I__11979 (
            .O(N__54932),
            .I(N__54929));
    Span4Mux_v I__11978 (
            .O(N__54929),
            .I(N__54926));
    Odrv4 I__11977 (
            .O(N__54926),
            .I(\PROM.ROMDATA.m19_ns ));
    CascadeMux I__11976 (
            .O(N__54923),
            .I(N__54919));
    InMux I__11975 (
            .O(N__54922),
            .I(N__54916));
    InMux I__11974 (
            .O(N__54919),
            .I(N__54913));
    LocalMux I__11973 (
            .O(N__54916),
            .I(N__54908));
    LocalMux I__11972 (
            .O(N__54913),
            .I(N__54908));
    Span4Mux_v I__11971 (
            .O(N__54908),
            .I(N__54905));
    Odrv4 I__11970 (
            .O(N__54905),
            .I(\PROM.ROMDATA.m33 ));
    InMux I__11969 (
            .O(N__54902),
            .I(N__54898));
    InMux I__11968 (
            .O(N__54901),
            .I(N__54895));
    LocalMux I__11967 (
            .O(N__54898),
            .I(\CONTROL.dout_reto_1 ));
    LocalMux I__11966 (
            .O(N__54895),
            .I(\CONTROL.dout_reto_1 ));
    InMux I__11965 (
            .O(N__54890),
            .I(N__54884));
    InMux I__11964 (
            .O(N__54889),
            .I(N__54884));
    LocalMux I__11963 (
            .O(N__54884),
            .I(N__54881));
    Span4Mux_v I__11962 (
            .O(N__54881),
            .I(N__54878));
    Odrv4 I__11961 (
            .O(N__54878),
            .I(\CONTROL.programCounter_1_reto_1 ));
    CascadeMux I__11960 (
            .O(N__54875),
            .I(\CONTROL.programCounter_ret_1_RNIH68IZ0Z_1_cascade_ ));
    InMux I__11959 (
            .O(N__54872),
            .I(N__54869));
    LocalMux I__11958 (
            .O(N__54869),
            .I(\CONTROL.programCounter_ret_19_RNIAK8JZ0Z_1 ));
    CascadeMux I__11957 (
            .O(N__54866),
            .I(progRomAddress_1_cascade_));
    InMux I__11956 (
            .O(N__54863),
            .I(N__54860));
    LocalMux I__11955 (
            .O(N__54860),
            .I(\PROM.ROMDATA.m437_ns ));
    InMux I__11954 (
            .O(N__54857),
            .I(N__54854));
    LocalMux I__11953 (
            .O(N__54854),
            .I(\PROM.ROMDATA.m312_bm ));
    InMux I__11952 (
            .O(N__54851),
            .I(N__54848));
    LocalMux I__11951 (
            .O(N__54848),
            .I(N__54845));
    Span4Mux_h I__11950 (
            .O(N__54845),
            .I(N__54842));
    Span4Mux_h I__11949 (
            .O(N__54842),
            .I(N__54839));
    Odrv4 I__11948 (
            .O(N__54839),
            .I(\PROM.ROMDATA.m312_am ));
    InMux I__11947 (
            .O(N__54836),
            .I(N__54833));
    LocalMux I__11946 (
            .O(N__54833),
            .I(\PROM.ROMDATA.m437_ns_1 ));
    InMux I__11945 (
            .O(N__54830),
            .I(N__54827));
    LocalMux I__11944 (
            .O(N__54827),
            .I(\PROM.ROMDATA.m11_bm ));
    CascadeMux I__11943 (
            .O(N__54824),
            .I(\PROM.ROMDATA.m18_bm_cascade_ ));
    InMux I__11942 (
            .O(N__54821),
            .I(N__54818));
    LocalMux I__11941 (
            .O(N__54818),
            .I(N__54815));
    Span12Mux_v I__11940 (
            .O(N__54815),
            .I(N__54811));
    InMux I__11939 (
            .O(N__54814),
            .I(N__54808));
    Odrv12 I__11938 (
            .O(N__54811),
            .I(\CONTROL.ctrlOut_2 ));
    LocalMux I__11937 (
            .O(N__54808),
            .I(\CONTROL.ctrlOut_2 ));
    InMux I__11936 (
            .O(N__54803),
            .I(N__54799));
    InMux I__11935 (
            .O(N__54802),
            .I(N__54796));
    LocalMux I__11934 (
            .O(N__54799),
            .I(N__54791));
    LocalMux I__11933 (
            .O(N__54796),
            .I(N__54791));
    Span4Mux_h I__11932 (
            .O(N__54791),
            .I(N__54788));
    Span4Mux_v I__11931 (
            .O(N__54788),
            .I(N__54785));
    Odrv4 I__11930 (
            .O(N__54785),
            .I(\CONTROL.dout_reto_2 ));
    InMux I__11929 (
            .O(N__54782),
            .I(N__54779));
    LocalMux I__11928 (
            .O(N__54779),
            .I(N__54776));
    Span12Mux_v I__11927 (
            .O(N__54776),
            .I(N__54773));
    Odrv12 I__11926 (
            .O(N__54773),
            .I(\CONTROL.N_136_0 ));
    InMux I__11925 (
            .O(N__54770),
            .I(N__54767));
    LocalMux I__11924 (
            .O(N__54767),
            .I(N__54763));
    InMux I__11923 (
            .O(N__54766),
            .I(N__54760));
    Span4Mux_v I__11922 (
            .O(N__54763),
            .I(N__54757));
    LocalMux I__11921 (
            .O(N__54760),
            .I(\CONTROL.N_86_0 ));
    Odrv4 I__11920 (
            .O(N__54757),
            .I(\CONTROL.N_86_0 ));
    CascadeMux I__11919 (
            .O(N__54752),
            .I(N__54747));
    InMux I__11918 (
            .O(N__54751),
            .I(N__54741));
    InMux I__11917 (
            .O(N__54750),
            .I(N__54741));
    InMux I__11916 (
            .O(N__54747),
            .I(N__54738));
    InMux I__11915 (
            .O(N__54746),
            .I(N__54735));
    LocalMux I__11914 (
            .O(N__54741),
            .I(N__54732));
    LocalMux I__11913 (
            .O(N__54738),
            .I(N__54729));
    LocalMux I__11912 (
            .O(N__54735),
            .I(N__54726));
    Span4Mux_v I__11911 (
            .O(N__54732),
            .I(N__54723));
    Span4Mux_h I__11910 (
            .O(N__54729),
            .I(N__54720));
    Span4Mux_v I__11909 (
            .O(N__54726),
            .I(N__54716));
    Span4Mux_h I__11908 (
            .O(N__54723),
            .I(N__54711));
    Span4Mux_v I__11907 (
            .O(N__54720),
            .I(N__54711));
    InMux I__11906 (
            .O(N__54719),
            .I(N__54708));
    Span4Mux_h I__11905 (
            .O(N__54716),
            .I(N__54702));
    Span4Mux_h I__11904 (
            .O(N__54711),
            .I(N__54702));
    LocalMux I__11903 (
            .O(N__54708),
            .I(N__54699));
    InMux I__11902 (
            .O(N__54707),
            .I(N__54696));
    Odrv4 I__11901 (
            .O(N__54702),
            .I(\CONTROL.N_98_0 ));
    Odrv4 I__11900 (
            .O(N__54699),
            .I(\CONTROL.N_98_0 ));
    LocalMux I__11899 (
            .O(N__54696),
            .I(\CONTROL.N_98_0 ));
    InMux I__11898 (
            .O(N__54689),
            .I(N__54682));
    InMux I__11897 (
            .O(N__54688),
            .I(N__54674));
    InMux I__11896 (
            .O(N__54687),
            .I(N__54671));
    InMux I__11895 (
            .O(N__54686),
            .I(N__54665));
    InMux I__11894 (
            .O(N__54685),
            .I(N__54662));
    LocalMux I__11893 (
            .O(N__54682),
            .I(N__54648));
    InMux I__11892 (
            .O(N__54681),
            .I(N__54641));
    InMux I__11891 (
            .O(N__54680),
            .I(N__54641));
    InMux I__11890 (
            .O(N__54679),
            .I(N__54641));
    InMux I__11889 (
            .O(N__54678),
            .I(N__54636));
    InMux I__11888 (
            .O(N__54677),
            .I(N__54636));
    LocalMux I__11887 (
            .O(N__54674),
            .I(N__54627));
    LocalMux I__11886 (
            .O(N__54671),
            .I(N__54627));
    InMux I__11885 (
            .O(N__54670),
            .I(N__54620));
    InMux I__11884 (
            .O(N__54669),
            .I(N__54620));
    InMux I__11883 (
            .O(N__54668),
            .I(N__54620));
    LocalMux I__11882 (
            .O(N__54665),
            .I(N__54615));
    LocalMux I__11881 (
            .O(N__54662),
            .I(N__54615));
    InMux I__11880 (
            .O(N__54661),
            .I(N__54612));
    InMux I__11879 (
            .O(N__54660),
            .I(N__54609));
    InMux I__11878 (
            .O(N__54659),
            .I(N__54602));
    InMux I__11877 (
            .O(N__54658),
            .I(N__54602));
    InMux I__11876 (
            .O(N__54657),
            .I(N__54602));
    InMux I__11875 (
            .O(N__54656),
            .I(N__54599));
    InMux I__11874 (
            .O(N__54655),
            .I(N__54596));
    InMux I__11873 (
            .O(N__54654),
            .I(N__54593));
    InMux I__11872 (
            .O(N__54653),
            .I(N__54588));
    InMux I__11871 (
            .O(N__54652),
            .I(N__54588));
    CascadeMux I__11870 (
            .O(N__54651),
            .I(N__54576));
    Span4Mux_v I__11869 (
            .O(N__54648),
            .I(N__54563));
    LocalMux I__11868 (
            .O(N__54641),
            .I(N__54563));
    LocalMux I__11867 (
            .O(N__54636),
            .I(N__54560));
    InMux I__11866 (
            .O(N__54635),
            .I(N__54553));
    InMux I__11865 (
            .O(N__54634),
            .I(N__54553));
    InMux I__11864 (
            .O(N__54633),
            .I(N__54553));
    InMux I__11863 (
            .O(N__54632),
            .I(N__54550));
    Span4Mux_h I__11862 (
            .O(N__54627),
            .I(N__54545));
    LocalMux I__11861 (
            .O(N__54620),
            .I(N__54545));
    Span4Mux_h I__11860 (
            .O(N__54615),
            .I(N__54536));
    LocalMux I__11859 (
            .O(N__54612),
            .I(N__54531));
    LocalMux I__11858 (
            .O(N__54609),
            .I(N__54531));
    LocalMux I__11857 (
            .O(N__54602),
            .I(N__54528));
    LocalMux I__11856 (
            .O(N__54599),
            .I(N__54519));
    LocalMux I__11855 (
            .O(N__54596),
            .I(N__54519));
    LocalMux I__11854 (
            .O(N__54593),
            .I(N__54519));
    LocalMux I__11853 (
            .O(N__54588),
            .I(N__54519));
    InMux I__11852 (
            .O(N__54587),
            .I(N__54514));
    InMux I__11851 (
            .O(N__54586),
            .I(N__54514));
    InMux I__11850 (
            .O(N__54585),
            .I(N__54511));
    InMux I__11849 (
            .O(N__54584),
            .I(N__54506));
    InMux I__11848 (
            .O(N__54583),
            .I(N__54506));
    InMux I__11847 (
            .O(N__54582),
            .I(N__54501));
    InMux I__11846 (
            .O(N__54581),
            .I(N__54501));
    InMux I__11845 (
            .O(N__54580),
            .I(N__54494));
    InMux I__11844 (
            .O(N__54579),
            .I(N__54494));
    InMux I__11843 (
            .O(N__54576),
            .I(N__54494));
    InMux I__11842 (
            .O(N__54575),
            .I(N__54491));
    InMux I__11841 (
            .O(N__54574),
            .I(N__54486));
    InMux I__11840 (
            .O(N__54573),
            .I(N__54486));
    InMux I__11839 (
            .O(N__54572),
            .I(N__54477));
    InMux I__11838 (
            .O(N__54571),
            .I(N__54477));
    InMux I__11837 (
            .O(N__54570),
            .I(N__54477));
    InMux I__11836 (
            .O(N__54569),
            .I(N__54477));
    InMux I__11835 (
            .O(N__54568),
            .I(N__54474));
    Span4Mux_h I__11834 (
            .O(N__54563),
            .I(N__54469));
    Span4Mux_v I__11833 (
            .O(N__54560),
            .I(N__54469));
    LocalMux I__11832 (
            .O(N__54553),
            .I(N__54466));
    LocalMux I__11831 (
            .O(N__54550),
            .I(N__54461));
    Span4Mux_h I__11830 (
            .O(N__54545),
            .I(N__54461));
    InMux I__11829 (
            .O(N__54544),
            .I(N__54458));
    InMux I__11828 (
            .O(N__54543),
            .I(N__54453));
    InMux I__11827 (
            .O(N__54542),
            .I(N__54453));
    InMux I__11826 (
            .O(N__54541),
            .I(N__54446));
    InMux I__11825 (
            .O(N__54540),
            .I(N__54446));
    InMux I__11824 (
            .O(N__54539),
            .I(N__54446));
    Span4Mux_v I__11823 (
            .O(N__54536),
            .I(N__54435));
    Span4Mux_v I__11822 (
            .O(N__54531),
            .I(N__54435));
    Span4Mux_h I__11821 (
            .O(N__54528),
            .I(N__54435));
    Span4Mux_v I__11820 (
            .O(N__54519),
            .I(N__54435));
    LocalMux I__11819 (
            .O(N__54514),
            .I(N__54435));
    LocalMux I__11818 (
            .O(N__54511),
            .I(N__54426));
    LocalMux I__11817 (
            .O(N__54506),
            .I(N__54426));
    LocalMux I__11816 (
            .O(N__54501),
            .I(N__54426));
    LocalMux I__11815 (
            .O(N__54494),
            .I(N__54426));
    LocalMux I__11814 (
            .O(N__54491),
            .I(controlWord_4));
    LocalMux I__11813 (
            .O(N__54486),
            .I(controlWord_4));
    LocalMux I__11812 (
            .O(N__54477),
            .I(controlWord_4));
    LocalMux I__11811 (
            .O(N__54474),
            .I(controlWord_4));
    Odrv4 I__11810 (
            .O(N__54469),
            .I(controlWord_4));
    Odrv4 I__11809 (
            .O(N__54466),
            .I(controlWord_4));
    Odrv4 I__11808 (
            .O(N__54461),
            .I(controlWord_4));
    LocalMux I__11807 (
            .O(N__54458),
            .I(controlWord_4));
    LocalMux I__11806 (
            .O(N__54453),
            .I(controlWord_4));
    LocalMux I__11805 (
            .O(N__54446),
            .I(controlWord_4));
    Odrv4 I__11804 (
            .O(N__54435),
            .I(controlWord_4));
    Odrv4 I__11803 (
            .O(N__54426),
            .I(controlWord_4));
    InMux I__11802 (
            .O(N__54401),
            .I(N__54398));
    LocalMux I__11801 (
            .O(N__54398),
            .I(\PROM.ROMDATA.m320_am ));
    InMux I__11800 (
            .O(N__54395),
            .I(N__54392));
    LocalMux I__11799 (
            .O(N__54392),
            .I(\PROM.ROMDATA.m150 ));
    CascadeMux I__11798 (
            .O(N__54389),
            .I(N__54386));
    InMux I__11797 (
            .O(N__54386),
            .I(N__54383));
    LocalMux I__11796 (
            .O(N__54383),
            .I(N__54380));
    Span12Mux_v I__11795 (
            .O(N__54380),
            .I(N__54377));
    Odrv12 I__11794 (
            .O(N__54377),
            .I(\PROM.ROMDATA.N_558_mux ));
    CascadeMux I__11793 (
            .O(N__54374),
            .I(\PROM.ROMDATA.m49_cascade_ ));
    InMux I__11792 (
            .O(N__54371),
            .I(N__54368));
    LocalMux I__11791 (
            .O(N__54368),
            .I(\PROM.ROMDATA.m229_1 ));
    CascadeMux I__11790 (
            .O(N__54365),
            .I(\PROM.ROMDATA.m228_bm_cascade_ ));
    InMux I__11789 (
            .O(N__54362),
            .I(N__54359));
    LocalMux I__11788 (
            .O(N__54359),
            .I(N__54352));
    InMux I__11787 (
            .O(N__54358),
            .I(N__54343));
    InMux I__11786 (
            .O(N__54357),
            .I(N__54343));
    InMux I__11785 (
            .O(N__54356),
            .I(N__54343));
    InMux I__11784 (
            .O(N__54355),
            .I(N__54343));
    Span4Mux_h I__11783 (
            .O(N__54352),
            .I(N__54338));
    LocalMux I__11782 (
            .O(N__54343),
            .I(N__54338));
    Span4Mux_h I__11781 (
            .O(N__54338),
            .I(N__54335));
    Span4Mux_h I__11780 (
            .O(N__54335),
            .I(N__54332));
    Odrv4 I__11779 (
            .O(N__54332),
            .I(\PROM.ROMDATA.m229 ));
    InMux I__11778 (
            .O(N__54329),
            .I(N__54323));
    InMux I__11777 (
            .O(N__54328),
            .I(N__54323));
    LocalMux I__11776 (
            .O(N__54323),
            .I(N__54320));
    Odrv12 I__11775 (
            .O(N__54320),
            .I(\ALU.dZ0Z_15 ));
    InMux I__11774 (
            .O(N__54317),
            .I(N__54314));
    LocalMux I__11773 (
            .O(N__54314),
            .I(N__54311));
    Odrv12 I__11772 (
            .O(N__54311),
            .I(\ALU.dout_6_ns_1_15 ));
    CascadeMux I__11771 (
            .O(N__54308),
            .I(N__54305));
    InMux I__11770 (
            .O(N__54305),
            .I(N__54300));
    InMux I__11769 (
            .O(N__54304),
            .I(N__54289));
    InMux I__11768 (
            .O(N__54303),
            .I(N__54286));
    LocalMux I__11767 (
            .O(N__54300),
            .I(N__54281));
    InMux I__11766 (
            .O(N__54299),
            .I(N__54276));
    InMux I__11765 (
            .O(N__54298),
            .I(N__54276));
    InMux I__11764 (
            .O(N__54297),
            .I(N__54271));
    InMux I__11763 (
            .O(N__54296),
            .I(N__54271));
    InMux I__11762 (
            .O(N__54295),
            .I(N__54266));
    InMux I__11761 (
            .O(N__54294),
            .I(N__54266));
    InMux I__11760 (
            .O(N__54293),
            .I(N__54261));
    InMux I__11759 (
            .O(N__54292),
            .I(N__54261));
    LocalMux I__11758 (
            .O(N__54289),
            .I(N__54258));
    LocalMux I__11757 (
            .O(N__54286),
            .I(N__54255));
    InMux I__11756 (
            .O(N__54285),
            .I(N__54250));
    InMux I__11755 (
            .O(N__54284),
            .I(N__54250));
    Span4Mux_h I__11754 (
            .O(N__54281),
            .I(N__54244));
    LocalMux I__11753 (
            .O(N__54276),
            .I(N__54244));
    LocalMux I__11752 (
            .O(N__54271),
            .I(N__54237));
    LocalMux I__11751 (
            .O(N__54266),
            .I(N__54237));
    LocalMux I__11750 (
            .O(N__54261),
            .I(N__54237));
    Span4Mux_h I__11749 (
            .O(N__54258),
            .I(N__54231));
    Span4Mux_h I__11748 (
            .O(N__54255),
            .I(N__54228));
    LocalMux I__11747 (
            .O(N__54250),
            .I(N__54225));
    InMux I__11746 (
            .O(N__54249),
            .I(N__54222));
    Span4Mux_h I__11745 (
            .O(N__54244),
            .I(N__54217));
    Span4Mux_h I__11744 (
            .O(N__54237),
            .I(N__54217));
    InMux I__11743 (
            .O(N__54236),
            .I(N__54212));
    InMux I__11742 (
            .O(N__54235),
            .I(N__54212));
    InMux I__11741 (
            .O(N__54234),
            .I(N__54209));
    Odrv4 I__11740 (
            .O(N__54231),
            .I(aluOperand1_1_rep2));
    Odrv4 I__11739 (
            .O(N__54228),
            .I(aluOperand1_1_rep2));
    Odrv4 I__11738 (
            .O(N__54225),
            .I(aluOperand1_1_rep2));
    LocalMux I__11737 (
            .O(N__54222),
            .I(aluOperand1_1_rep2));
    Odrv4 I__11736 (
            .O(N__54217),
            .I(aluOperand1_1_rep2));
    LocalMux I__11735 (
            .O(N__54212),
            .I(aluOperand1_1_rep2));
    LocalMux I__11734 (
            .O(N__54209),
            .I(aluOperand1_1_rep2));
    InMux I__11733 (
            .O(N__54194),
            .I(N__54191));
    LocalMux I__11732 (
            .O(N__54191),
            .I(N__54188));
    Span12Mux_v I__11731 (
            .O(N__54188),
            .I(N__54183));
    InMux I__11730 (
            .O(N__54187),
            .I(N__54178));
    InMux I__11729 (
            .O(N__54186),
            .I(N__54178));
    Span12Mux_v I__11728 (
            .O(N__54183),
            .I(N__54175));
    LocalMux I__11727 (
            .O(N__54178),
            .I(N__54172));
    Span12Mux_h I__11726 (
            .O(N__54175),
            .I(N__54169));
    Span4Mux_v I__11725 (
            .O(N__54172),
            .I(N__54166));
    Odrv12 I__11724 (
            .O(N__54169),
            .I(h_15));
    Odrv4 I__11723 (
            .O(N__54166),
            .I(h_15));
    InMux I__11722 (
            .O(N__54161),
            .I(N__54158));
    LocalMux I__11721 (
            .O(N__54158),
            .I(N__54155));
    Span4Mux_h I__11720 (
            .O(N__54155),
            .I(N__54152));
    Span4Mux_h I__11719 (
            .O(N__54152),
            .I(N__54149));
    Odrv4 I__11718 (
            .O(N__54149),
            .I(\ALU.N_1100 ));
    CascadeMux I__11717 (
            .O(N__54146),
            .I(\ALU.N_1148_cascade_ ));
    InMux I__11716 (
            .O(N__54143),
            .I(N__54135));
    InMux I__11715 (
            .O(N__54142),
            .I(N__54131));
    InMux I__11714 (
            .O(N__54141),
            .I(N__54125));
    InMux I__11713 (
            .O(N__54140),
            .I(N__54122));
    InMux I__11712 (
            .O(N__54139),
            .I(N__54119));
    InMux I__11711 (
            .O(N__54138),
            .I(N__54115));
    LocalMux I__11710 (
            .O(N__54135),
            .I(N__54107));
    InMux I__11709 (
            .O(N__54134),
            .I(N__54104));
    LocalMux I__11708 (
            .O(N__54131),
            .I(N__54101));
    InMux I__11707 (
            .O(N__54130),
            .I(N__54098));
    InMux I__11706 (
            .O(N__54129),
            .I(N__54093));
    InMux I__11705 (
            .O(N__54128),
            .I(N__54093));
    LocalMux I__11704 (
            .O(N__54125),
            .I(N__54090));
    LocalMux I__11703 (
            .O(N__54122),
            .I(N__54085));
    LocalMux I__11702 (
            .O(N__54119),
            .I(N__54085));
    InMux I__11701 (
            .O(N__54118),
            .I(N__54082));
    LocalMux I__11700 (
            .O(N__54115),
            .I(N__54079));
    InMux I__11699 (
            .O(N__54114),
            .I(N__54074));
    InMux I__11698 (
            .O(N__54113),
            .I(N__54074));
    InMux I__11697 (
            .O(N__54112),
            .I(N__54069));
    InMux I__11696 (
            .O(N__54111),
            .I(N__54069));
    InMux I__11695 (
            .O(N__54110),
            .I(N__54066));
    Span4Mux_h I__11694 (
            .O(N__54107),
            .I(N__54063));
    LocalMux I__11693 (
            .O(N__54104),
            .I(N__54056));
    Span4Mux_v I__11692 (
            .O(N__54101),
            .I(N__54047));
    LocalMux I__11691 (
            .O(N__54098),
            .I(N__54047));
    LocalMux I__11690 (
            .O(N__54093),
            .I(N__54047));
    Span4Mux_h I__11689 (
            .O(N__54090),
            .I(N__54047));
    Span4Mux_h I__11688 (
            .O(N__54085),
            .I(N__54042));
    LocalMux I__11687 (
            .O(N__54082),
            .I(N__54042));
    Span4Mux_v I__11686 (
            .O(N__54079),
            .I(N__54034));
    LocalMux I__11685 (
            .O(N__54074),
            .I(N__54034));
    LocalMux I__11684 (
            .O(N__54069),
            .I(N__54034));
    LocalMux I__11683 (
            .O(N__54066),
            .I(N__54029));
    Span4Mux_v I__11682 (
            .O(N__54063),
            .I(N__54029));
    InMux I__11681 (
            .O(N__54062),
            .I(N__54022));
    InMux I__11680 (
            .O(N__54061),
            .I(N__54022));
    InMux I__11679 (
            .O(N__54060),
            .I(N__54022));
    InMux I__11678 (
            .O(N__54059),
            .I(N__54019));
    Span4Mux_v I__11677 (
            .O(N__54056),
            .I(N__54012));
    Span4Mux_h I__11676 (
            .O(N__54047),
            .I(N__54012));
    Span4Mux_h I__11675 (
            .O(N__54042),
            .I(N__54012));
    InMux I__11674 (
            .O(N__54041),
            .I(N__54009));
    Span4Mux_h I__11673 (
            .O(N__54034),
            .I(N__54006));
    Span4Mux_v I__11672 (
            .O(N__54029),
            .I(N__54001));
    LocalMux I__11671 (
            .O(N__54022),
            .I(N__54001));
    LocalMux I__11670 (
            .O(N__54019),
            .I(aluOperand1_0));
    Odrv4 I__11669 (
            .O(N__54012),
            .I(aluOperand1_0));
    LocalMux I__11668 (
            .O(N__54009),
            .I(aluOperand1_0));
    Odrv4 I__11667 (
            .O(N__54006),
            .I(aluOperand1_0));
    Odrv4 I__11666 (
            .O(N__54001),
            .I(aluOperand1_0));
    InMux I__11665 (
            .O(N__53990),
            .I(N__53987));
    LocalMux I__11664 (
            .O(N__53987),
            .I(\ALU.N_1260 ));
    InMux I__11663 (
            .O(N__53984),
            .I(N__53981));
    LocalMux I__11662 (
            .O(N__53981),
            .I(N__53978));
    Span4Mux_h I__11661 (
            .O(N__53978),
            .I(N__53975));
    Span4Mux_h I__11660 (
            .O(N__53975),
            .I(N__53972));
    Odrv4 I__11659 (
            .O(N__53972),
            .I(\ALU.N_1212 ));
    CascadeMux I__11658 (
            .O(N__53969),
            .I(N__53958));
    InMux I__11657 (
            .O(N__53968),
            .I(N__53953));
    InMux I__11656 (
            .O(N__53967),
            .I(N__53946));
    InMux I__11655 (
            .O(N__53966),
            .I(N__53946));
    InMux I__11654 (
            .O(N__53965),
            .I(N__53943));
    InMux I__11653 (
            .O(N__53964),
            .I(N__53931));
    InMux I__11652 (
            .O(N__53963),
            .I(N__53931));
    InMux I__11651 (
            .O(N__53962),
            .I(N__53924));
    InMux I__11650 (
            .O(N__53961),
            .I(N__53924));
    InMux I__11649 (
            .O(N__53958),
            .I(N__53924));
    InMux I__11648 (
            .O(N__53957),
            .I(N__53919));
    InMux I__11647 (
            .O(N__53956),
            .I(N__53919));
    LocalMux I__11646 (
            .O(N__53953),
            .I(N__53916));
    InMux I__11645 (
            .O(N__53952),
            .I(N__53911));
    InMux I__11644 (
            .O(N__53951),
            .I(N__53911));
    LocalMux I__11643 (
            .O(N__53946),
            .I(N__53904));
    LocalMux I__11642 (
            .O(N__53943),
            .I(N__53904));
    InMux I__11641 (
            .O(N__53942),
            .I(N__53899));
    InMux I__11640 (
            .O(N__53941),
            .I(N__53899));
    CascadeMux I__11639 (
            .O(N__53940),
            .I(N__53895));
    InMux I__11638 (
            .O(N__53939),
            .I(N__53890));
    InMux I__11637 (
            .O(N__53938),
            .I(N__53890));
    InMux I__11636 (
            .O(N__53937),
            .I(N__53882));
    InMux I__11635 (
            .O(N__53936),
            .I(N__53882));
    LocalMux I__11634 (
            .O(N__53931),
            .I(N__53879));
    LocalMux I__11633 (
            .O(N__53924),
            .I(N__53876));
    LocalMux I__11632 (
            .O(N__53919),
            .I(N__53873));
    Span4Mux_v I__11631 (
            .O(N__53916),
            .I(N__53870));
    LocalMux I__11630 (
            .O(N__53911),
            .I(N__53867));
    InMux I__11629 (
            .O(N__53910),
            .I(N__53862));
    InMux I__11628 (
            .O(N__53909),
            .I(N__53862));
    Span4Mux_h I__11627 (
            .O(N__53904),
            .I(N__53856));
    LocalMux I__11626 (
            .O(N__53899),
            .I(N__53853));
    InMux I__11625 (
            .O(N__53898),
            .I(N__53848));
    InMux I__11624 (
            .O(N__53895),
            .I(N__53848));
    LocalMux I__11623 (
            .O(N__53890),
            .I(N__53845));
    InMux I__11622 (
            .O(N__53889),
            .I(N__53842));
    InMux I__11621 (
            .O(N__53888),
            .I(N__53837));
    InMux I__11620 (
            .O(N__53887),
            .I(N__53837));
    LocalMux I__11619 (
            .O(N__53882),
            .I(N__53828));
    Span4Mux_v I__11618 (
            .O(N__53879),
            .I(N__53828));
    Span4Mux_h I__11617 (
            .O(N__53876),
            .I(N__53828));
    Span4Mux_v I__11616 (
            .O(N__53873),
            .I(N__53828));
    Span4Mux_h I__11615 (
            .O(N__53870),
            .I(N__53823));
    Span4Mux_v I__11614 (
            .O(N__53867),
            .I(N__53823));
    LocalMux I__11613 (
            .O(N__53862),
            .I(N__53820));
    InMux I__11612 (
            .O(N__53861),
            .I(N__53817));
    InMux I__11611 (
            .O(N__53860),
            .I(N__53812));
    InMux I__11610 (
            .O(N__53859),
            .I(N__53812));
    Span4Mux_h I__11609 (
            .O(N__53856),
            .I(N__53805));
    Span4Mux_h I__11608 (
            .O(N__53853),
            .I(N__53805));
    LocalMux I__11607 (
            .O(N__53848),
            .I(N__53805));
    Span4Mux_h I__11606 (
            .O(N__53845),
            .I(N__53796));
    LocalMux I__11605 (
            .O(N__53842),
            .I(N__53796));
    LocalMux I__11604 (
            .O(N__53837),
            .I(N__53796));
    Span4Mux_h I__11603 (
            .O(N__53828),
            .I(N__53796));
    Odrv4 I__11602 (
            .O(N__53823),
            .I(aluOperand2_0));
    Odrv12 I__11601 (
            .O(N__53820),
            .I(aluOperand2_0));
    LocalMux I__11600 (
            .O(N__53817),
            .I(aluOperand2_0));
    LocalMux I__11599 (
            .O(N__53812),
            .I(aluOperand2_0));
    Odrv4 I__11598 (
            .O(N__53805),
            .I(aluOperand2_0));
    Odrv4 I__11597 (
            .O(N__53796),
            .I(aluOperand2_0));
    InMux I__11596 (
            .O(N__53783),
            .I(N__53780));
    LocalMux I__11595 (
            .O(N__53780),
            .I(N__53777));
    Span4Mux_v I__11594 (
            .O(N__53777),
            .I(N__53774));
    Sp12to4 I__11593 (
            .O(N__53774),
            .I(N__53771));
    Span12Mux_h I__11592 (
            .O(N__53771),
            .I(N__53768));
    Odrv12 I__11591 (
            .O(N__53768),
            .I(\ALU.combOperand2_d_bmZ0Z_15 ));
    CascadeMux I__11590 (
            .O(N__53765),
            .I(\ALU.c_RNI8VV95Z0Z_15_cascade_ ));
    InMux I__11589 (
            .O(N__53762),
            .I(N__53759));
    LocalMux I__11588 (
            .O(N__53759),
            .I(N__53754));
    InMux I__11587 (
            .O(N__53758),
            .I(N__53749));
    InMux I__11586 (
            .O(N__53757),
            .I(N__53749));
    Odrv4 I__11585 (
            .O(N__53754),
            .I(\ALU.c_RNIJTKD7Z0Z_15 ));
    LocalMux I__11584 (
            .O(N__53749),
            .I(\ALU.c_RNIJTKD7Z0Z_15 ));
    CascadeMux I__11583 (
            .O(N__53744),
            .I(\PROM.ROMDATA.m320_bm_cascade_ ));
    InMux I__11582 (
            .O(N__53741),
            .I(N__53738));
    LocalMux I__11581 (
            .O(N__53738),
            .I(\PROM.ROMDATA.m410_am ));
    CascadeMux I__11580 (
            .O(N__53735),
            .I(\PROM.ROMDATA.m413_am_cascade_ ));
    CascadeMux I__11579 (
            .O(N__53732),
            .I(\ALU.status_e_0_RNO_0Z0Z_2_cascade_ ));
    CascadeMux I__11578 (
            .O(N__53729),
            .I(\ALU.N_570_cascade_ ));
    InMux I__11577 (
            .O(N__53726),
            .I(N__53723));
    LocalMux I__11576 (
            .O(N__53723),
            .I(\ALU.status_e_0_RNO_1Z0Z_2 ));
    InMux I__11575 (
            .O(N__53720),
            .I(N__53714));
    InMux I__11574 (
            .O(N__53719),
            .I(N__53709));
    InMux I__11573 (
            .O(N__53718),
            .I(N__53709));
    CascadeMux I__11572 (
            .O(N__53717),
            .I(N__53706));
    LocalMux I__11571 (
            .O(N__53714),
            .I(N__53701));
    LocalMux I__11570 (
            .O(N__53709),
            .I(N__53698));
    InMux I__11569 (
            .O(N__53706),
            .I(N__53691));
    InMux I__11568 (
            .O(N__53705),
            .I(N__53691));
    InMux I__11567 (
            .O(N__53704),
            .I(N__53691));
    Span4Mux_v I__11566 (
            .O(N__53701),
            .I(N__53682));
    Span4Mux_v I__11565 (
            .O(N__53698),
            .I(N__53682));
    LocalMux I__11564 (
            .O(N__53691),
            .I(N__53682));
    InMux I__11563 (
            .O(N__53690),
            .I(N__53677));
    InMux I__11562 (
            .O(N__53689),
            .I(N__53677));
    Span4Mux_v I__11561 (
            .O(N__53682),
            .I(N__53674));
    LocalMux I__11560 (
            .O(N__53677),
            .I(aluStatus_2));
    Odrv4 I__11559 (
            .O(N__53674),
            .I(aluStatus_2));
    InMux I__11558 (
            .O(N__53669),
            .I(N__53663));
    InMux I__11557 (
            .O(N__53668),
            .I(N__53658));
    InMux I__11556 (
            .O(N__53667),
            .I(N__53653));
    InMux I__11555 (
            .O(N__53666),
            .I(N__53653));
    LocalMux I__11554 (
            .O(N__53663),
            .I(N__53650));
    InMux I__11553 (
            .O(N__53662),
            .I(N__53645));
    InMux I__11552 (
            .O(N__53661),
            .I(N__53645));
    LocalMux I__11551 (
            .O(N__53658),
            .I(N__53642));
    LocalMux I__11550 (
            .O(N__53653),
            .I(N__53639));
    Span4Mux_h I__11549 (
            .O(N__53650),
            .I(N__53636));
    LocalMux I__11548 (
            .O(N__53645),
            .I(PROM_ROMDATA_dintern_9ro));
    Odrv12 I__11547 (
            .O(N__53642),
            .I(PROM_ROMDATA_dintern_9ro));
    Odrv4 I__11546 (
            .O(N__53639),
            .I(PROM_ROMDATA_dintern_9ro));
    Odrv4 I__11545 (
            .O(N__53636),
            .I(PROM_ROMDATA_dintern_9ro));
    InMux I__11544 (
            .O(N__53627),
            .I(N__53624));
    LocalMux I__11543 (
            .O(N__53624),
            .I(N__53621));
    Span4Mux_v I__11542 (
            .O(N__53621),
            .I(N__53618));
    Span4Mux_h I__11541 (
            .O(N__53618),
            .I(N__53615));
    Odrv4 I__11540 (
            .O(N__53615),
            .I(\CONTROL.g3Z0Z_0 ));
    InMux I__11539 (
            .O(N__53612),
            .I(N__53608));
    InMux I__11538 (
            .O(N__53611),
            .I(N__53605));
    LocalMux I__11537 (
            .O(N__53608),
            .I(N__53602));
    LocalMux I__11536 (
            .O(N__53605),
            .I(N__53599));
    Span12Mux_h I__11535 (
            .O(N__53602),
            .I(N__53596));
    Span4Mux_v I__11534 (
            .O(N__53599),
            .I(N__53593));
    Odrv12 I__11533 (
            .O(N__53596),
            .I(\ALU.bZ0Z_15 ));
    Odrv4 I__11532 (
            .O(N__53593),
            .I(\ALU.bZ0Z_15 ));
    InMux I__11531 (
            .O(N__53588),
            .I(N__53585));
    LocalMux I__11530 (
            .O(N__53585),
            .I(N__53580));
    InMux I__11529 (
            .O(N__53584),
            .I(N__53575));
    InMux I__11528 (
            .O(N__53583),
            .I(N__53575));
    Span4Mux_v I__11527 (
            .O(N__53580),
            .I(N__53567));
    LocalMux I__11526 (
            .O(N__53575),
            .I(N__53564));
    InMux I__11525 (
            .O(N__53574),
            .I(N__53561));
    InMux I__11524 (
            .O(N__53573),
            .I(N__53558));
    InMux I__11523 (
            .O(N__53572),
            .I(N__53555));
    InMux I__11522 (
            .O(N__53571),
            .I(N__53550));
    InMux I__11521 (
            .O(N__53570),
            .I(N__53550));
    Span4Mux_h I__11520 (
            .O(N__53567),
            .I(N__53545));
    Span4Mux_v I__11519 (
            .O(N__53564),
            .I(N__53545));
    LocalMux I__11518 (
            .O(N__53561),
            .I(aluOperand2_fast_2));
    LocalMux I__11517 (
            .O(N__53558),
            .I(aluOperand2_fast_2));
    LocalMux I__11516 (
            .O(N__53555),
            .I(aluOperand2_fast_2));
    LocalMux I__11515 (
            .O(N__53550),
            .I(aluOperand2_fast_2));
    Odrv4 I__11514 (
            .O(N__53545),
            .I(aluOperand2_fast_2));
    CascadeMux I__11513 (
            .O(N__53534),
            .I(N__53531));
    InMux I__11512 (
            .O(N__53531),
            .I(N__53527));
    CascadeMux I__11511 (
            .O(N__53530),
            .I(N__53524));
    LocalMux I__11510 (
            .O(N__53527),
            .I(N__53521));
    InMux I__11509 (
            .O(N__53524),
            .I(N__53518));
    Span4Mux_h I__11508 (
            .O(N__53521),
            .I(N__53514));
    LocalMux I__11507 (
            .O(N__53518),
            .I(N__53511));
    CascadeMux I__11506 (
            .O(N__53517),
            .I(N__53508));
    Span4Mux_v I__11505 (
            .O(N__53514),
            .I(N__53505));
    Span4Mux_v I__11504 (
            .O(N__53511),
            .I(N__53502));
    InMux I__11503 (
            .O(N__53508),
            .I(N__53499));
    Sp12to4 I__11502 (
            .O(N__53505),
            .I(N__53496));
    Sp12to4 I__11501 (
            .O(N__53502),
            .I(N__53493));
    LocalMux I__11500 (
            .O(N__53499),
            .I(N__53490));
    Span12Mux_v I__11499 (
            .O(N__53496),
            .I(N__53485));
    Span12Mux_h I__11498 (
            .O(N__53493),
            .I(N__53485));
    Odrv4 I__11497 (
            .O(N__53490),
            .I(f_15));
    Odrv12 I__11496 (
            .O(N__53485),
            .I(f_15));
    InMux I__11495 (
            .O(N__53480),
            .I(N__53474));
    InMux I__11494 (
            .O(N__53479),
            .I(N__53471));
    InMux I__11493 (
            .O(N__53478),
            .I(N__53468));
    InMux I__11492 (
            .O(N__53477),
            .I(N__53463));
    LocalMux I__11491 (
            .O(N__53474),
            .I(N__53458));
    LocalMux I__11490 (
            .O(N__53471),
            .I(N__53458));
    LocalMux I__11489 (
            .O(N__53468),
            .I(N__53455));
    InMux I__11488 (
            .O(N__53467),
            .I(N__53450));
    InMux I__11487 (
            .O(N__53466),
            .I(N__53450));
    LocalMux I__11486 (
            .O(N__53463),
            .I(N__53445));
    Span4Mux_v I__11485 (
            .O(N__53458),
            .I(N__53445));
    Odrv12 I__11484 (
            .O(N__53455),
            .I(aluOperand2_fast_1));
    LocalMux I__11483 (
            .O(N__53450),
            .I(aluOperand2_fast_1));
    Odrv4 I__11482 (
            .O(N__53445),
            .I(aluOperand2_fast_1));
    CascadeMux I__11481 (
            .O(N__53438),
            .I(\ALU.operand2_6_ns_1_15_cascade_ ));
    InMux I__11480 (
            .O(N__53435),
            .I(N__53431));
    InMux I__11479 (
            .O(N__53434),
            .I(N__53426));
    LocalMux I__11478 (
            .O(N__53431),
            .I(N__53422));
    InMux I__11477 (
            .O(N__53430),
            .I(N__53417));
    InMux I__11476 (
            .O(N__53429),
            .I(N__53417));
    LocalMux I__11475 (
            .O(N__53426),
            .I(N__53414));
    InMux I__11474 (
            .O(N__53425),
            .I(N__53411));
    Span4Mux_h I__11473 (
            .O(N__53422),
            .I(N__53407));
    LocalMux I__11472 (
            .O(N__53417),
            .I(N__53402));
    Span4Mux_h I__11471 (
            .O(N__53414),
            .I(N__53395));
    LocalMux I__11470 (
            .O(N__53411),
            .I(N__53395));
    InMux I__11469 (
            .O(N__53410),
            .I(N__53392));
    Span4Mux_h I__11468 (
            .O(N__53407),
            .I(N__53389));
    InMux I__11467 (
            .O(N__53406),
            .I(N__53384));
    InMux I__11466 (
            .O(N__53405),
            .I(N__53384));
    Span4Mux_h I__11465 (
            .O(N__53402),
            .I(N__53381));
    InMux I__11464 (
            .O(N__53401),
            .I(N__53376));
    InMux I__11463 (
            .O(N__53400),
            .I(N__53376));
    Odrv4 I__11462 (
            .O(N__53395),
            .I(aluOperand2_1_rep1));
    LocalMux I__11461 (
            .O(N__53392),
            .I(aluOperand2_1_rep1));
    Odrv4 I__11460 (
            .O(N__53389),
            .I(aluOperand2_1_rep1));
    LocalMux I__11459 (
            .O(N__53384),
            .I(aluOperand2_1_rep1));
    Odrv4 I__11458 (
            .O(N__53381),
            .I(aluOperand2_1_rep1));
    LocalMux I__11457 (
            .O(N__53376),
            .I(aluOperand2_1_rep1));
    CascadeMux I__11456 (
            .O(N__53363),
            .I(\ALU.status_14_0_0_cascade_ ));
    CascadeMux I__11455 (
            .O(N__53360),
            .I(N__53357));
    InMux I__11454 (
            .O(N__53357),
            .I(N__53354));
    LocalMux I__11453 (
            .O(N__53354),
            .I(N__53351));
    Span4Mux_v I__11452 (
            .O(N__53351),
            .I(N__53348));
    Odrv4 I__11451 (
            .O(N__53348),
            .I(\ALU.status_14_5_0 ));
    CascadeMux I__11450 (
            .O(N__53345),
            .I(\ALU.status_14_7_0_cascade_ ));
    InMux I__11449 (
            .O(N__53342),
            .I(N__53339));
    LocalMux I__11448 (
            .O(N__53339),
            .I(N__53336));
    Odrv4 I__11447 (
            .O(N__53336),
            .I(\ALU.status_14_13_0 ));
    InMux I__11446 (
            .O(N__53333),
            .I(N__53329));
    InMux I__11445 (
            .O(N__53332),
            .I(N__53326));
    LocalMux I__11444 (
            .O(N__53329),
            .I(N__53323));
    LocalMux I__11443 (
            .O(N__53326),
            .I(N__53320));
    Span4Mux_h I__11442 (
            .O(N__53323),
            .I(N__53317));
    Span4Mux_v I__11441 (
            .O(N__53320),
            .I(N__53314));
    Odrv4 I__11440 (
            .O(N__53317),
            .I(\ALU.N_979 ));
    Odrv4 I__11439 (
            .O(N__53314),
            .I(\ALU.N_979 ));
    CascadeMux I__11438 (
            .O(N__53309),
            .I(\ALU.N_979_cascade_ ));
    InMux I__11437 (
            .O(N__53306),
            .I(N__53285));
    InMux I__11436 (
            .O(N__53305),
            .I(N__53282));
    InMux I__11435 (
            .O(N__53304),
            .I(N__53275));
    InMux I__11434 (
            .O(N__53303),
            .I(N__53275));
    InMux I__11433 (
            .O(N__53302),
            .I(N__53275));
    CascadeMux I__11432 (
            .O(N__53301),
            .I(N__53272));
    InMux I__11431 (
            .O(N__53300),
            .I(N__53267));
    InMux I__11430 (
            .O(N__53299),
            .I(N__53267));
    InMux I__11429 (
            .O(N__53298),
            .I(N__53264));
    InMux I__11428 (
            .O(N__53297),
            .I(N__53259));
    InMux I__11427 (
            .O(N__53296),
            .I(N__53259));
    InMux I__11426 (
            .O(N__53295),
            .I(N__53250));
    InMux I__11425 (
            .O(N__53294),
            .I(N__53250));
    InMux I__11424 (
            .O(N__53293),
            .I(N__53250));
    InMux I__11423 (
            .O(N__53292),
            .I(N__53250));
    CascadeMux I__11422 (
            .O(N__53291),
            .I(N__53246));
    InMux I__11421 (
            .O(N__53290),
            .I(N__53242));
    InMux I__11420 (
            .O(N__53289),
            .I(N__53239));
    CascadeMux I__11419 (
            .O(N__53288),
            .I(N__53234));
    LocalMux I__11418 (
            .O(N__53285),
            .I(N__53226));
    LocalMux I__11417 (
            .O(N__53282),
            .I(N__53226));
    LocalMux I__11416 (
            .O(N__53275),
            .I(N__53223));
    InMux I__11415 (
            .O(N__53272),
            .I(N__53220));
    LocalMux I__11414 (
            .O(N__53267),
            .I(N__53217));
    LocalMux I__11413 (
            .O(N__53264),
            .I(N__53209));
    LocalMux I__11412 (
            .O(N__53259),
            .I(N__53209));
    LocalMux I__11411 (
            .O(N__53250),
            .I(N__53209));
    CascadeMux I__11410 (
            .O(N__53249),
            .I(N__53206));
    InMux I__11409 (
            .O(N__53246),
            .I(N__53201));
    InMux I__11408 (
            .O(N__53245),
            .I(N__53198));
    LocalMux I__11407 (
            .O(N__53242),
            .I(N__53195));
    LocalMux I__11406 (
            .O(N__53239),
            .I(N__53192));
    InMux I__11405 (
            .O(N__53238),
            .I(N__53187));
    InMux I__11404 (
            .O(N__53237),
            .I(N__53187));
    InMux I__11403 (
            .O(N__53234),
            .I(N__53184));
    InMux I__11402 (
            .O(N__53233),
            .I(N__53181));
    InMux I__11401 (
            .O(N__53232),
            .I(N__53178));
    InMux I__11400 (
            .O(N__53231),
            .I(N__53174));
    Span4Mux_v I__11399 (
            .O(N__53226),
            .I(N__53171));
    Span4Mux_v I__11398 (
            .O(N__53223),
            .I(N__53166));
    LocalMux I__11397 (
            .O(N__53220),
            .I(N__53166));
    Span4Mux_v I__11396 (
            .O(N__53217),
            .I(N__53162));
    InMux I__11395 (
            .O(N__53216),
            .I(N__53158));
    Span4Mux_v I__11394 (
            .O(N__53209),
            .I(N__53155));
    InMux I__11393 (
            .O(N__53206),
            .I(N__53152));
    InMux I__11392 (
            .O(N__53205),
            .I(N__53147));
    InMux I__11391 (
            .O(N__53204),
            .I(N__53147));
    LocalMux I__11390 (
            .O(N__53201),
            .I(N__53141));
    LocalMux I__11389 (
            .O(N__53198),
            .I(N__53138));
    Span4Mux_h I__11388 (
            .O(N__53195),
            .I(N__53133));
    Span4Mux_h I__11387 (
            .O(N__53192),
            .I(N__53133));
    LocalMux I__11386 (
            .O(N__53187),
            .I(N__53130));
    LocalMux I__11385 (
            .O(N__53184),
            .I(N__53127));
    LocalMux I__11384 (
            .O(N__53181),
            .I(N__53122));
    LocalMux I__11383 (
            .O(N__53178),
            .I(N__53122));
    InMux I__11382 (
            .O(N__53177),
            .I(N__53119));
    LocalMux I__11381 (
            .O(N__53174),
            .I(N__53112));
    Span4Mux_h I__11380 (
            .O(N__53171),
            .I(N__53112));
    Span4Mux_v I__11379 (
            .O(N__53166),
            .I(N__53112));
    InMux I__11378 (
            .O(N__53165),
            .I(N__53109));
    Span4Mux_h I__11377 (
            .O(N__53162),
            .I(N__53106));
    InMux I__11376 (
            .O(N__53161),
            .I(N__53103));
    LocalMux I__11375 (
            .O(N__53158),
            .I(N__53094));
    Span4Mux_h I__11374 (
            .O(N__53155),
            .I(N__53094));
    LocalMux I__11373 (
            .O(N__53152),
            .I(N__53094));
    LocalMux I__11372 (
            .O(N__53147),
            .I(N__53094));
    InMux I__11371 (
            .O(N__53146),
            .I(N__53089));
    InMux I__11370 (
            .O(N__53145),
            .I(N__53089));
    InMux I__11369 (
            .O(N__53144),
            .I(N__53086));
    Span4Mux_h I__11368 (
            .O(N__53141),
            .I(N__53079));
    Span4Mux_h I__11367 (
            .O(N__53138),
            .I(N__53079));
    Span4Mux_v I__11366 (
            .O(N__53133),
            .I(N__53079));
    Span4Mux_h I__11365 (
            .O(N__53130),
            .I(N__53072));
    Span4Mux_v I__11364 (
            .O(N__53127),
            .I(N__53072));
    Span4Mux_h I__11363 (
            .O(N__53122),
            .I(N__53072));
    LocalMux I__11362 (
            .O(N__53119),
            .I(N__53067));
    Sp12to4 I__11361 (
            .O(N__53112),
            .I(N__53067));
    LocalMux I__11360 (
            .O(N__53109),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    Odrv4 I__11359 (
            .O(N__53106),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    LocalMux I__11358 (
            .O(N__53103),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    Odrv4 I__11357 (
            .O(N__53094),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    LocalMux I__11356 (
            .O(N__53089),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    LocalMux I__11355 (
            .O(N__53086),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    Odrv4 I__11354 (
            .O(N__53079),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    Odrv4 I__11353 (
            .O(N__53072),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    Odrv12 I__11352 (
            .O(N__53067),
            .I(\ALU.combOperand2_a0_0Z0Z_6 ));
    InMux I__11351 (
            .O(N__53048),
            .I(N__53045));
    LocalMux I__11350 (
            .O(N__53045),
            .I(N__53042));
    Span4Mux_v I__11349 (
            .O(N__53042),
            .I(N__53039));
    Odrv4 I__11348 (
            .O(N__53039),
            .I(\ALU.status_RNO_22Z0Z_0 ));
    InMux I__11347 (
            .O(N__53036),
            .I(N__53033));
    LocalMux I__11346 (
            .O(N__53033),
            .I(\ALU.status_14_6_0 ));
    InMux I__11345 (
            .O(N__53030),
            .I(N__53027));
    LocalMux I__11344 (
            .O(N__53027),
            .I(N__53024));
    Sp12to4 I__11343 (
            .O(N__53024),
            .I(N__53021));
    Span12Mux_v I__11342 (
            .O(N__53021),
            .I(N__53018));
    Span12Mux_h I__11341 (
            .O(N__53018),
            .I(N__53015));
    Odrv12 I__11340 (
            .O(N__53015),
            .I(\ALU.status_17_I_21_c_RNOZ0 ));
    InMux I__11339 (
            .O(N__53012),
            .I(N__53003));
    InMux I__11338 (
            .O(N__53011),
            .I(N__53000));
    InMux I__11337 (
            .O(N__53010),
            .I(N__52997));
    InMux I__11336 (
            .O(N__53009),
            .I(N__52994));
    InMux I__11335 (
            .O(N__53008),
            .I(N__52991));
    InMux I__11334 (
            .O(N__53007),
            .I(N__52988));
    InMux I__11333 (
            .O(N__53006),
            .I(N__52984));
    LocalMux I__11332 (
            .O(N__53003),
            .I(N__52981));
    LocalMux I__11331 (
            .O(N__53000),
            .I(N__52974));
    LocalMux I__11330 (
            .O(N__52997),
            .I(N__52974));
    LocalMux I__11329 (
            .O(N__52994),
            .I(N__52974));
    LocalMux I__11328 (
            .O(N__52991),
            .I(N__52971));
    LocalMux I__11327 (
            .O(N__52988),
            .I(N__52968));
    InMux I__11326 (
            .O(N__52987),
            .I(N__52965));
    LocalMux I__11325 (
            .O(N__52984),
            .I(N__52958));
    Span4Mux_h I__11324 (
            .O(N__52981),
            .I(N__52958));
    Span4Mux_v I__11323 (
            .O(N__52974),
            .I(N__52958));
    Span4Mux_h I__11322 (
            .O(N__52971),
            .I(N__52953));
    Span4Mux_h I__11321 (
            .O(N__52968),
            .I(N__52953));
    LocalMux I__11320 (
            .O(N__52965),
            .I(N__52950));
    Span4Mux_h I__11319 (
            .O(N__52958),
            .I(N__52947));
    Span4Mux_h I__11318 (
            .O(N__52953),
            .I(N__52942));
    Span4Mux_h I__11317 (
            .O(N__52950),
            .I(N__52942));
    Odrv4 I__11316 (
            .O(N__52947),
            .I(\ALU.mult_15 ));
    Odrv4 I__11315 (
            .O(N__52942),
            .I(\ALU.mult_15 ));
    InMux I__11314 (
            .O(N__52937),
            .I(N__52928));
    InMux I__11313 (
            .O(N__52936),
            .I(N__52925));
    InMux I__11312 (
            .O(N__52935),
            .I(N__52922));
    InMux I__11311 (
            .O(N__52934),
            .I(N__52919));
    InMux I__11310 (
            .O(N__52933),
            .I(N__52916));
    InMux I__11309 (
            .O(N__52932),
            .I(N__52913));
    InMux I__11308 (
            .O(N__52931),
            .I(N__52910));
    LocalMux I__11307 (
            .O(N__52928),
            .I(N__52905));
    LocalMux I__11306 (
            .O(N__52925),
            .I(N__52905));
    LocalMux I__11305 (
            .O(N__52922),
            .I(N__52902));
    LocalMux I__11304 (
            .O(N__52919),
            .I(\ALU.a_15_1_15 ));
    LocalMux I__11303 (
            .O(N__52916),
            .I(\ALU.a_15_1_15 ));
    LocalMux I__11302 (
            .O(N__52913),
            .I(\ALU.a_15_1_15 ));
    LocalMux I__11301 (
            .O(N__52910),
            .I(\ALU.a_15_1_15 ));
    Odrv4 I__11300 (
            .O(N__52905),
            .I(\ALU.a_15_1_15 ));
    Odrv4 I__11299 (
            .O(N__52902),
            .I(\ALU.a_15_1_15 ));
    CascadeMux I__11298 (
            .O(N__52889),
            .I(N__52886));
    InMux I__11297 (
            .O(N__52886),
            .I(N__52883));
    LocalMux I__11296 (
            .O(N__52883),
            .I(N__52880));
    Span4Mux_v I__11295 (
            .O(N__52880),
            .I(N__52875));
    InMux I__11294 (
            .O(N__52879),
            .I(N__52872));
    InMux I__11293 (
            .O(N__52878),
            .I(N__52867));
    Span4Mux_h I__11292 (
            .O(N__52875),
            .I(N__52863));
    LocalMux I__11291 (
            .O(N__52872),
            .I(N__52860));
    InMux I__11290 (
            .O(N__52871),
            .I(N__52857));
    InMux I__11289 (
            .O(N__52870),
            .I(N__52853));
    LocalMux I__11288 (
            .O(N__52867),
            .I(N__52850));
    InMux I__11287 (
            .O(N__52866),
            .I(N__52847));
    Span4Mux_v I__11286 (
            .O(N__52863),
            .I(N__52844));
    Span4Mux_v I__11285 (
            .O(N__52860),
            .I(N__52839));
    LocalMux I__11284 (
            .O(N__52857),
            .I(N__52839));
    InMux I__11283 (
            .O(N__52856),
            .I(N__52836));
    LocalMux I__11282 (
            .O(N__52853),
            .I(N__52833));
    Span4Mux_v I__11281 (
            .O(N__52850),
            .I(N__52830));
    LocalMux I__11280 (
            .O(N__52847),
            .I(N__52825));
    Span4Mux_h I__11279 (
            .O(N__52844),
            .I(N__52825));
    Span4Mux_h I__11278 (
            .O(N__52839),
            .I(N__52822));
    LocalMux I__11277 (
            .O(N__52836),
            .I(N__52813));
    Span4Mux_v I__11276 (
            .O(N__52833),
            .I(N__52813));
    Span4Mux_v I__11275 (
            .O(N__52830),
            .I(N__52813));
    Span4Mux_v I__11274 (
            .O(N__52825),
            .I(N__52813));
    Odrv4 I__11273 (
            .O(N__52822),
            .I(\ALU.a_15_m1_9 ));
    Odrv4 I__11272 (
            .O(N__52813),
            .I(\ALU.a_15_m1_9 ));
    InMux I__11271 (
            .O(N__52808),
            .I(N__52802));
    CascadeMux I__11270 (
            .O(N__52807),
            .I(N__52798));
    InMux I__11269 (
            .O(N__52806),
            .I(N__52795));
    InMux I__11268 (
            .O(N__52805),
            .I(N__52792));
    LocalMux I__11267 (
            .O(N__52802),
            .I(N__52789));
    InMux I__11266 (
            .O(N__52801),
            .I(N__52783));
    InMux I__11265 (
            .O(N__52798),
            .I(N__52780));
    LocalMux I__11264 (
            .O(N__52795),
            .I(N__52777));
    LocalMux I__11263 (
            .O(N__52792),
            .I(N__52772));
    Span4Mux_v I__11262 (
            .O(N__52789),
            .I(N__52772));
    InMux I__11261 (
            .O(N__52788),
            .I(N__52769));
    InMux I__11260 (
            .O(N__52787),
            .I(N__52766));
    InMux I__11259 (
            .O(N__52786),
            .I(N__52763));
    LocalMux I__11258 (
            .O(N__52783),
            .I(N__52754));
    LocalMux I__11257 (
            .O(N__52780),
            .I(N__52754));
    Span4Mux_v I__11256 (
            .O(N__52777),
            .I(N__52754));
    Span4Mux_h I__11255 (
            .O(N__52772),
            .I(N__52754));
    LocalMux I__11254 (
            .O(N__52769),
            .I(\ALU.mult_546_c_RNIJOT4JZ0Z8 ));
    LocalMux I__11253 (
            .O(N__52766),
            .I(\ALU.mult_546_c_RNIJOT4JZ0Z8 ));
    LocalMux I__11252 (
            .O(N__52763),
            .I(\ALU.mult_546_c_RNIJOT4JZ0Z8 ));
    Odrv4 I__11251 (
            .O(N__52754),
            .I(\ALU.mult_546_c_RNIJOT4JZ0Z8 ));
    InMux I__11250 (
            .O(N__52745),
            .I(N__52741));
    InMux I__11249 (
            .O(N__52744),
            .I(N__52738));
    LocalMux I__11248 (
            .O(N__52741),
            .I(N__52735));
    LocalMux I__11247 (
            .O(N__52738),
            .I(N__52732));
    Span4Mux_v I__11246 (
            .O(N__52735),
            .I(N__52729));
    Span4Mux_v I__11245 (
            .O(N__52732),
            .I(N__52726));
    Span4Mux_h I__11244 (
            .O(N__52729),
            .I(N__52723));
    Span4Mux_h I__11243 (
            .O(N__52726),
            .I(N__52720));
    Span4Mux_h I__11242 (
            .O(N__52723),
            .I(N__52717));
    Span4Mux_v I__11241 (
            .O(N__52720),
            .I(N__52714));
    Odrv4 I__11240 (
            .O(N__52717),
            .I(\ALU.dZ0Z_9 ));
    Odrv4 I__11239 (
            .O(N__52714),
            .I(\ALU.dZ0Z_9 ));
    InMux I__11238 (
            .O(N__52709),
            .I(N__52706));
    LocalMux I__11237 (
            .O(N__52706),
            .I(N__52702));
    InMux I__11236 (
            .O(N__52705),
            .I(N__52699));
    Span4Mux_v I__11235 (
            .O(N__52702),
            .I(N__52696));
    LocalMux I__11234 (
            .O(N__52699),
            .I(\ALU.N_835 ));
    Odrv4 I__11233 (
            .O(N__52696),
            .I(\ALU.N_835 ));
    CascadeMux I__11232 (
            .O(N__52691),
            .I(\ALU.d_RNIPFFDD1_0Z0Z_6_cascade_ ));
    CascadeMux I__11231 (
            .O(N__52688),
            .I(\ALU.N_863_cascade_ ));
    InMux I__11230 (
            .O(N__52685),
            .I(N__52680));
    InMux I__11229 (
            .O(N__52684),
            .I(N__52675));
    InMux I__11228 (
            .O(N__52683),
            .I(N__52672));
    LocalMux I__11227 (
            .O(N__52680),
            .I(N__52669));
    InMux I__11226 (
            .O(N__52679),
            .I(N__52666));
    InMux I__11225 (
            .O(N__52678),
            .I(N__52663));
    LocalMux I__11224 (
            .O(N__52675),
            .I(N__52660));
    LocalMux I__11223 (
            .O(N__52672),
            .I(N__52657));
    Span12Mux_h I__11222 (
            .O(N__52669),
            .I(N__52654));
    LocalMux I__11221 (
            .O(N__52666),
            .I(N__52645));
    LocalMux I__11220 (
            .O(N__52663),
            .I(N__52645));
    Span12Mux_v I__11219 (
            .O(N__52660),
            .I(N__52645));
    Span12Mux_h I__11218 (
            .O(N__52657),
            .I(N__52645));
    Odrv12 I__11217 (
            .O(N__52654),
            .I(\ALU.d_RNIN3H0DZ0Z_3 ));
    Odrv12 I__11216 (
            .O(N__52645),
            .I(\ALU.d_RNIN3H0DZ0Z_3 ));
    CascadeMux I__11215 (
            .O(N__52640),
            .I(\ALU.d_RNIGPBNB6Z0Z_2_cascade_ ));
    InMux I__11214 (
            .O(N__52637),
            .I(N__52632));
    CascadeMux I__11213 (
            .O(N__52636),
            .I(N__52629));
    InMux I__11212 (
            .O(N__52635),
            .I(N__52624));
    LocalMux I__11211 (
            .O(N__52632),
            .I(N__52620));
    InMux I__11210 (
            .O(N__52629),
            .I(N__52616));
    InMux I__11209 (
            .O(N__52628),
            .I(N__52613));
    InMux I__11208 (
            .O(N__52627),
            .I(N__52609));
    LocalMux I__11207 (
            .O(N__52624),
            .I(N__52606));
    InMux I__11206 (
            .O(N__52623),
            .I(N__52603));
    Span4Mux_h I__11205 (
            .O(N__52620),
            .I(N__52600));
    InMux I__11204 (
            .O(N__52619),
            .I(N__52597));
    LocalMux I__11203 (
            .O(N__52616),
            .I(N__52592));
    LocalMux I__11202 (
            .O(N__52613),
            .I(N__52592));
    InMux I__11201 (
            .O(N__52612),
            .I(N__52589));
    LocalMux I__11200 (
            .O(N__52609),
            .I(N__52586));
    Span4Mux_h I__11199 (
            .O(N__52606),
            .I(N__52583));
    LocalMux I__11198 (
            .O(N__52603),
            .I(N__52580));
    Span4Mux_h I__11197 (
            .O(N__52600),
            .I(N__52577));
    LocalMux I__11196 (
            .O(N__52597),
            .I(N__52572));
    Span4Mux_v I__11195 (
            .O(N__52592),
            .I(N__52572));
    LocalMux I__11194 (
            .O(N__52589),
            .I(N__52565));
    Span4Mux_h I__11193 (
            .O(N__52586),
            .I(N__52565));
    Span4Mux_v I__11192 (
            .O(N__52583),
            .I(N__52565));
    Span4Mux_h I__11191 (
            .O(N__52580),
            .I(N__52562));
    Span4Mux_h I__11190 (
            .O(N__52577),
            .I(N__52559));
    Span4Mux_h I__11189 (
            .O(N__52572),
            .I(N__52556));
    Sp12to4 I__11188 (
            .O(N__52565),
            .I(N__52553));
    Span4Mux_h I__11187 (
            .O(N__52562),
            .I(N__52548));
    Span4Mux_v I__11186 (
            .O(N__52559),
            .I(N__52548));
    Odrv4 I__11185 (
            .O(N__52556),
            .I(\ALU.a_15_m0_5 ));
    Odrv12 I__11184 (
            .O(N__52553),
            .I(\ALU.a_15_m0_5 ));
    Odrv4 I__11183 (
            .O(N__52548),
            .I(\ALU.a_15_m0_5 ));
    IoInMux I__11182 (
            .O(N__52541),
            .I(N__52538));
    LocalMux I__11181 (
            .O(N__52538),
            .I(N__52535));
    IoSpan4Mux I__11180 (
            .O(N__52535),
            .I(N__52532));
    IoSpan4Mux I__11179 (
            .O(N__52532),
            .I(N__52528));
    IoInMux I__11178 (
            .O(N__52531),
            .I(N__52524));
    Span4Mux_s2_h I__11177 (
            .O(N__52528),
            .I(N__52521));
    InMux I__11176 (
            .O(N__52527),
            .I(N__52518));
    LocalMux I__11175 (
            .O(N__52524),
            .I(N__52515));
    Sp12to4 I__11174 (
            .O(N__52521),
            .I(N__52510));
    LocalMux I__11173 (
            .O(N__52518),
            .I(N__52510));
    Span12Mux_s8_h I__11172 (
            .O(N__52515),
            .I(N__52507));
    Span12Mux_h I__11171 (
            .O(N__52510),
            .I(N__52504));
    Odrv12 I__11170 (
            .O(N__52507),
            .I(bus_5));
    Odrv12 I__11169 (
            .O(N__52504),
            .I(bus_5));
    InMux I__11168 (
            .O(N__52499),
            .I(N__52496));
    LocalMux I__11167 (
            .O(N__52496),
            .I(\ALU.c_RNINGV0T2Z0Z_15 ));
    InMux I__11166 (
            .O(N__52493),
            .I(N__52490));
    LocalMux I__11165 (
            .O(N__52490),
            .I(\ALU.d_RNIPFFDD1Z0Z_6 ));
    CascadeMux I__11164 (
            .O(N__52487),
            .I(N__52484));
    InMux I__11163 (
            .O(N__52484),
            .I(N__52481));
    LocalMux I__11162 (
            .O(N__52481),
            .I(N__52478));
    Span4Mux_h I__11161 (
            .O(N__52478),
            .I(N__52474));
    InMux I__11160 (
            .O(N__52477),
            .I(N__52471));
    Span4Mux_h I__11159 (
            .O(N__52474),
            .I(N__52468));
    LocalMux I__11158 (
            .O(N__52471),
            .I(N__52465));
    Span4Mux_v I__11157 (
            .O(N__52468),
            .I(N__52462));
    Span4Mux_h I__11156 (
            .O(N__52465),
            .I(N__52459));
    Span4Mux_v I__11155 (
            .O(N__52462),
            .I(N__52456));
    Odrv4 I__11154 (
            .O(N__52459),
            .I(\ALU.eZ0Z_13 ));
    Odrv4 I__11153 (
            .O(N__52456),
            .I(\ALU.eZ0Z_13 ));
    CascadeMux I__11152 (
            .O(N__52451),
            .I(N__52448));
    InMux I__11151 (
            .O(N__52448),
            .I(N__52444));
    InMux I__11150 (
            .O(N__52447),
            .I(N__52441));
    LocalMux I__11149 (
            .O(N__52444),
            .I(N__52438));
    LocalMux I__11148 (
            .O(N__52441),
            .I(N__52435));
    Span4Mux_h I__11147 (
            .O(N__52438),
            .I(N__52432));
    Span4Mux_h I__11146 (
            .O(N__52435),
            .I(N__52429));
    Span4Mux_h I__11145 (
            .O(N__52432),
            .I(N__52426));
    Span4Mux_h I__11144 (
            .O(N__52429),
            .I(N__52423));
    Sp12to4 I__11143 (
            .O(N__52426),
            .I(N__52420));
    Span4Mux_v I__11142 (
            .O(N__52423),
            .I(N__52417));
    Odrv12 I__11141 (
            .O(N__52420),
            .I(\ALU.eZ0Z_14 ));
    Odrv4 I__11140 (
            .O(N__52417),
            .I(\ALU.eZ0Z_14 ));
    InMux I__11139 (
            .O(N__52412),
            .I(N__52407));
    InMux I__11138 (
            .O(N__52411),
            .I(N__52404));
    InMux I__11137 (
            .O(N__52410),
            .I(N__52401));
    LocalMux I__11136 (
            .O(N__52407),
            .I(N__52398));
    LocalMux I__11135 (
            .O(N__52404),
            .I(N__52395));
    LocalMux I__11134 (
            .O(N__52401),
            .I(N__52392));
    Span4Mux_h I__11133 (
            .O(N__52398),
            .I(N__52389));
    Span4Mux_v I__11132 (
            .O(N__52395),
            .I(N__52386));
    Span4Mux_v I__11131 (
            .O(N__52392),
            .I(N__52383));
    Span4Mux_h I__11130 (
            .O(N__52389),
            .I(N__52380));
    Span4Mux_h I__11129 (
            .O(N__52386),
            .I(N__52375));
    Span4Mux_v I__11128 (
            .O(N__52383),
            .I(N__52375));
    Span4Mux_h I__11127 (
            .O(N__52380),
            .I(N__52372));
    Span4Mux_h I__11126 (
            .O(N__52375),
            .I(N__52369));
    Span4Mux_v I__11125 (
            .O(N__52372),
            .I(N__52366));
    Span4Mux_h I__11124 (
            .O(N__52369),
            .I(N__52363));
    Odrv4 I__11123 (
            .O(N__52366),
            .I(g_12));
    Odrv4 I__11122 (
            .O(N__52363),
            .I(g_12));
    InMux I__11121 (
            .O(N__52358),
            .I(N__52354));
    CascadeMux I__11120 (
            .O(N__52357),
            .I(N__52351));
    LocalMux I__11119 (
            .O(N__52354),
            .I(N__52347));
    InMux I__11118 (
            .O(N__52351),
            .I(N__52344));
    InMux I__11117 (
            .O(N__52350),
            .I(N__52341));
    Span4Mux_v I__11116 (
            .O(N__52347),
            .I(N__52338));
    LocalMux I__11115 (
            .O(N__52344),
            .I(N__52335));
    LocalMux I__11114 (
            .O(N__52341),
            .I(N__52332));
    Span4Mux_h I__11113 (
            .O(N__52338),
            .I(N__52329));
    Sp12to4 I__11112 (
            .O(N__52335),
            .I(N__52326));
    Span4Mux_v I__11111 (
            .O(N__52332),
            .I(N__52323));
    Span4Mux_h I__11110 (
            .O(N__52329),
            .I(N__52320));
    Span12Mux_v I__11109 (
            .O(N__52326),
            .I(N__52315));
    Sp12to4 I__11108 (
            .O(N__52323),
            .I(N__52315));
    Sp12to4 I__11107 (
            .O(N__52320),
            .I(N__52312));
    Span12Mux_h I__11106 (
            .O(N__52315),
            .I(N__52307));
    Span12Mux_s10_h I__11105 (
            .O(N__52312),
            .I(N__52307));
    Odrv12 I__11104 (
            .O(N__52307),
            .I(g_13));
    InMux I__11103 (
            .O(N__52304),
            .I(N__52301));
    LocalMux I__11102 (
            .O(N__52301),
            .I(N__52298));
    Span4Mux_v I__11101 (
            .O(N__52298),
            .I(N__52295));
    Span4Mux_h I__11100 (
            .O(N__52295),
            .I(N__52292));
    Span4Mux_h I__11099 (
            .O(N__52292),
            .I(N__52288));
    InMux I__11098 (
            .O(N__52291),
            .I(N__52285));
    Span4Mux_h I__11097 (
            .O(N__52288),
            .I(N__52281));
    LocalMux I__11096 (
            .O(N__52285),
            .I(N__52278));
    InMux I__11095 (
            .O(N__52284),
            .I(N__52275));
    Span4Mux_v I__11094 (
            .O(N__52281),
            .I(N__52270));
    Span4Mux_h I__11093 (
            .O(N__52278),
            .I(N__52270));
    LocalMux I__11092 (
            .O(N__52275),
            .I(N__52267));
    Span4Mux_h I__11091 (
            .O(N__52270),
            .I(N__52264));
    Span4Mux_h I__11090 (
            .O(N__52267),
            .I(N__52261));
    Span4Mux_h I__11089 (
            .O(N__52264),
            .I(N__52258));
    Span4Mux_v I__11088 (
            .O(N__52261),
            .I(N__52255));
    Span4Mux_v I__11087 (
            .O(N__52258),
            .I(N__52252));
    Odrv4 I__11086 (
            .O(N__52255),
            .I(g_14));
    Odrv4 I__11085 (
            .O(N__52252),
            .I(g_14));
    CascadeMux I__11084 (
            .O(N__52247),
            .I(N__52242));
    CascadeMux I__11083 (
            .O(N__52246),
            .I(N__52237));
    CascadeMux I__11082 (
            .O(N__52245),
            .I(N__52233));
    InMux I__11081 (
            .O(N__52242),
            .I(N__52230));
    InMux I__11080 (
            .O(N__52241),
            .I(N__52227));
    InMux I__11079 (
            .O(N__52240),
            .I(N__52224));
    InMux I__11078 (
            .O(N__52237),
            .I(N__52220));
    InMux I__11077 (
            .O(N__52236),
            .I(N__52217));
    InMux I__11076 (
            .O(N__52233),
            .I(N__52214));
    LocalMux I__11075 (
            .O(N__52230),
            .I(N__52211));
    LocalMux I__11074 (
            .O(N__52227),
            .I(N__52206));
    LocalMux I__11073 (
            .O(N__52224),
            .I(N__52206));
    InMux I__11072 (
            .O(N__52223),
            .I(N__52202));
    LocalMux I__11071 (
            .O(N__52220),
            .I(N__52199));
    LocalMux I__11070 (
            .O(N__52217),
            .I(N__52196));
    LocalMux I__11069 (
            .O(N__52214),
            .I(N__52189));
    Span4Mux_h I__11068 (
            .O(N__52211),
            .I(N__52189));
    Span4Mux_v I__11067 (
            .O(N__52206),
            .I(N__52189));
    InMux I__11066 (
            .O(N__52205),
            .I(N__52186));
    LocalMux I__11065 (
            .O(N__52202),
            .I(N__52183));
    Span4Mux_h I__11064 (
            .O(N__52199),
            .I(N__52178));
    Span4Mux_v I__11063 (
            .O(N__52196),
            .I(N__52178));
    Span4Mux_h I__11062 (
            .O(N__52189),
            .I(N__52175));
    LocalMux I__11061 (
            .O(N__52186),
            .I(\ALU.a_15_ns_1_1 ));
    Odrv4 I__11060 (
            .O(N__52183),
            .I(\ALU.a_15_ns_1_1 ));
    Odrv4 I__11059 (
            .O(N__52178),
            .I(\ALU.a_15_ns_1_1 ));
    Odrv4 I__11058 (
            .O(N__52175),
            .I(\ALU.a_15_ns_1_1 ));
    InMux I__11057 (
            .O(N__52166),
            .I(N__52162));
    InMux I__11056 (
            .O(N__52165),
            .I(N__52159));
    LocalMux I__11055 (
            .O(N__52162),
            .I(N__52156));
    LocalMux I__11054 (
            .O(N__52159),
            .I(N__52153));
    Span4Mux_v I__11053 (
            .O(N__52156),
            .I(N__52150));
    Span4Mux_v I__11052 (
            .O(N__52153),
            .I(N__52147));
    Span4Mux_h I__11051 (
            .O(N__52150),
            .I(N__52144));
    Span4Mux_h I__11050 (
            .O(N__52147),
            .I(N__52141));
    Span4Mux_h I__11049 (
            .O(N__52144),
            .I(N__52138));
    Span4Mux_h I__11048 (
            .O(N__52141),
            .I(N__52135));
    Span4Mux_v I__11047 (
            .O(N__52138),
            .I(N__52132));
    Span4Mux_h I__11046 (
            .O(N__52135),
            .I(N__52129));
    Odrv4 I__11045 (
            .O(N__52132),
            .I(\ALU.dZ0Z_1 ));
    Odrv4 I__11044 (
            .O(N__52129),
            .I(\ALU.dZ0Z_1 ));
    InMux I__11043 (
            .O(N__52124),
            .I(N__52119));
    InMux I__11042 (
            .O(N__52123),
            .I(N__52114));
    InMux I__11041 (
            .O(N__52122),
            .I(N__52111));
    LocalMux I__11040 (
            .O(N__52119),
            .I(N__52108));
    InMux I__11039 (
            .O(N__52118),
            .I(N__52105));
    InMux I__11038 (
            .O(N__52117),
            .I(N__52102));
    LocalMux I__11037 (
            .O(N__52114),
            .I(N__52097));
    LocalMux I__11036 (
            .O(N__52111),
            .I(N__52097));
    Span4Mux_v I__11035 (
            .O(N__52108),
            .I(N__52093));
    LocalMux I__11034 (
            .O(N__52105),
            .I(N__52090));
    LocalMux I__11033 (
            .O(N__52102),
            .I(N__52087));
    Span4Mux_v I__11032 (
            .O(N__52097),
            .I(N__52084));
    InMux I__11031 (
            .O(N__52096),
            .I(N__52081));
    Span4Mux_h I__11030 (
            .O(N__52093),
            .I(N__52077));
    Span4Mux_v I__11029 (
            .O(N__52090),
            .I(N__52072));
    Span4Mux_v I__11028 (
            .O(N__52087),
            .I(N__52072));
    Sp12to4 I__11027 (
            .O(N__52084),
            .I(N__52067));
    LocalMux I__11026 (
            .O(N__52081),
            .I(N__52067));
    InMux I__11025 (
            .O(N__52080),
            .I(N__52064));
    Odrv4 I__11024 (
            .O(N__52077),
            .I(\ALU.d_RNINUGCF4Z0Z_0 ));
    Odrv4 I__11023 (
            .O(N__52072),
            .I(\ALU.d_RNINUGCF4Z0Z_0 ));
    Odrv12 I__11022 (
            .O(N__52067),
            .I(\ALU.d_RNINUGCF4Z0Z_0 ));
    LocalMux I__11021 (
            .O(N__52064),
            .I(\ALU.d_RNINUGCF4Z0Z_0 ));
    InMux I__11020 (
            .O(N__52055),
            .I(N__52046));
    InMux I__11019 (
            .O(N__52054),
            .I(N__52043));
    InMux I__11018 (
            .O(N__52053),
            .I(N__52040));
    InMux I__11017 (
            .O(N__52052),
            .I(N__52037));
    InMux I__11016 (
            .O(N__52051),
            .I(N__52034));
    InMux I__11015 (
            .O(N__52050),
            .I(N__52030));
    InMux I__11014 (
            .O(N__52049),
            .I(N__52027));
    LocalMux I__11013 (
            .O(N__52046),
            .I(N__52024));
    LocalMux I__11012 (
            .O(N__52043),
            .I(N__52021));
    LocalMux I__11011 (
            .O(N__52040),
            .I(N__52014));
    LocalMux I__11010 (
            .O(N__52037),
            .I(N__52014));
    LocalMux I__11009 (
            .O(N__52034),
            .I(N__52014));
    InMux I__11008 (
            .O(N__52033),
            .I(N__52011));
    LocalMux I__11007 (
            .O(N__52030),
            .I(N__52008));
    LocalMux I__11006 (
            .O(N__52027),
            .I(N__52005));
    Span4Mux_h I__11005 (
            .O(N__52024),
            .I(N__52002));
    Span4Mux_v I__11004 (
            .O(N__52021),
            .I(N__51999));
    Span4Mux_v I__11003 (
            .O(N__52014),
            .I(N__51996));
    LocalMux I__11002 (
            .O(N__52011),
            .I(N__51989));
    Span4Mux_h I__11001 (
            .O(N__52008),
            .I(N__51989));
    Span4Mux_v I__11000 (
            .O(N__52005),
            .I(N__51989));
    Span4Mux_v I__10999 (
            .O(N__52002),
            .I(N__51986));
    Span4Mux_v I__10998 (
            .O(N__51999),
            .I(N__51981));
    Span4Mux_v I__10997 (
            .O(N__51996),
            .I(N__51981));
    Span4Mux_v I__10996 (
            .O(N__51989),
            .I(N__51978));
    Odrv4 I__10995 (
            .O(N__51986),
            .I(\ALU.rshift_0 ));
    Odrv4 I__10994 (
            .O(N__51981),
            .I(\ALU.rshift_0 ));
    Odrv4 I__10993 (
            .O(N__51978),
            .I(\ALU.rshift_0 ));
    InMux I__10992 (
            .O(N__51971),
            .I(N__51968));
    LocalMux I__10991 (
            .O(N__51968),
            .I(N__51964));
    InMux I__10990 (
            .O(N__51967),
            .I(N__51961));
    Span4Mux_v I__10989 (
            .O(N__51964),
            .I(N__51958));
    LocalMux I__10988 (
            .O(N__51961),
            .I(N__51955));
    Span4Mux_h I__10987 (
            .O(N__51958),
            .I(N__51952));
    Span4Mux_v I__10986 (
            .O(N__51955),
            .I(N__51949));
    Span4Mux_h I__10985 (
            .O(N__51952),
            .I(N__51946));
    Span4Mux_h I__10984 (
            .O(N__51949),
            .I(N__51941));
    Span4Mux_v I__10983 (
            .O(N__51946),
            .I(N__51941));
    Odrv4 I__10982 (
            .O(N__51941),
            .I(\ALU.dZ0Z_0 ));
    CascadeMux I__10981 (
            .O(N__51938),
            .I(N__51934));
    InMux I__10980 (
            .O(N__51937),
            .I(N__51926));
    InMux I__10979 (
            .O(N__51934),
            .I(N__51923));
    CascadeMux I__10978 (
            .O(N__51933),
            .I(N__51920));
    InMux I__10977 (
            .O(N__51932),
            .I(N__51917));
    InMux I__10976 (
            .O(N__51931),
            .I(N__51914));
    InMux I__10975 (
            .O(N__51930),
            .I(N__51911));
    InMux I__10974 (
            .O(N__51929),
            .I(N__51908));
    LocalMux I__10973 (
            .O(N__51926),
            .I(N__51905));
    LocalMux I__10972 (
            .O(N__51923),
            .I(N__51901));
    InMux I__10971 (
            .O(N__51920),
            .I(N__51898));
    LocalMux I__10970 (
            .O(N__51917),
            .I(N__51893));
    LocalMux I__10969 (
            .O(N__51914),
            .I(N__51893));
    LocalMux I__10968 (
            .O(N__51911),
            .I(N__51886));
    LocalMux I__10967 (
            .O(N__51908),
            .I(N__51886));
    Span4Mux_v I__10966 (
            .O(N__51905),
            .I(N__51886));
    InMux I__10965 (
            .O(N__51904),
            .I(N__51883));
    Span4Mux_h I__10964 (
            .O(N__51901),
            .I(N__51880));
    LocalMux I__10963 (
            .O(N__51898),
            .I(N__51875));
    Span4Mux_v I__10962 (
            .O(N__51893),
            .I(N__51875));
    Span4Mux_v I__10961 (
            .O(N__51886),
            .I(N__51872));
    LocalMux I__10960 (
            .O(N__51883),
            .I(\ALU.a_15_m0_7 ));
    Odrv4 I__10959 (
            .O(N__51880),
            .I(\ALU.a_15_m0_7 ));
    Odrv4 I__10958 (
            .O(N__51875),
            .I(\ALU.a_15_m0_7 ));
    Odrv4 I__10957 (
            .O(N__51872),
            .I(\ALU.a_15_m0_7 ));
    CascadeMux I__10956 (
            .O(N__51863),
            .I(N__51859));
    InMux I__10955 (
            .O(N__51862),
            .I(N__51854));
    InMux I__10954 (
            .O(N__51859),
            .I(N__51848));
    InMux I__10953 (
            .O(N__51858),
            .I(N__51845));
    InMux I__10952 (
            .O(N__51857),
            .I(N__51842));
    LocalMux I__10951 (
            .O(N__51854),
            .I(N__51839));
    InMux I__10950 (
            .O(N__51853),
            .I(N__51836));
    InMux I__10949 (
            .O(N__51852),
            .I(N__51833));
    InMux I__10948 (
            .O(N__51851),
            .I(N__51830));
    LocalMux I__10947 (
            .O(N__51848),
            .I(N__51827));
    LocalMux I__10946 (
            .O(N__51845),
            .I(N__51824));
    LocalMux I__10945 (
            .O(N__51842),
            .I(N__51819));
    Span4Mux_v I__10944 (
            .O(N__51839),
            .I(N__51819));
    LocalMux I__10943 (
            .O(N__51836),
            .I(\ALU.mult_492_c_RNIGN2JECZ0 ));
    LocalMux I__10942 (
            .O(N__51833),
            .I(\ALU.mult_492_c_RNIGN2JECZ0 ));
    LocalMux I__10941 (
            .O(N__51830),
            .I(\ALU.mult_492_c_RNIGN2JECZ0 ));
    Odrv4 I__10940 (
            .O(N__51827),
            .I(\ALU.mult_492_c_RNIGN2JECZ0 ));
    Odrv4 I__10939 (
            .O(N__51824),
            .I(\ALU.mult_492_c_RNIGN2JECZ0 ));
    Odrv4 I__10938 (
            .O(N__51819),
            .I(\ALU.mult_492_c_RNIGN2JECZ0 ));
    InMux I__10937 (
            .O(N__51806),
            .I(N__51802));
    InMux I__10936 (
            .O(N__51805),
            .I(N__51799));
    LocalMux I__10935 (
            .O(N__51802),
            .I(N__51794));
    LocalMux I__10934 (
            .O(N__51799),
            .I(N__51794));
    Span4Mux_v I__10933 (
            .O(N__51794),
            .I(N__51791));
    Odrv4 I__10932 (
            .O(N__51791),
            .I(\ALU.dZ0Z_7 ));
    CascadeMux I__10931 (
            .O(N__51788),
            .I(N__51785));
    InMux I__10930 (
            .O(N__51785),
            .I(N__51780));
    InMux I__10929 (
            .O(N__51784),
            .I(N__51772));
    InMux I__10928 (
            .O(N__51783),
            .I(N__51769));
    LocalMux I__10927 (
            .O(N__51780),
            .I(N__51766));
    InMux I__10926 (
            .O(N__51779),
            .I(N__51763));
    InMux I__10925 (
            .O(N__51778),
            .I(N__51760));
    InMux I__10924 (
            .O(N__51777),
            .I(N__51757));
    InMux I__10923 (
            .O(N__51776),
            .I(N__51754));
    InMux I__10922 (
            .O(N__51775),
            .I(N__51751));
    LocalMux I__10921 (
            .O(N__51772),
            .I(N__51748));
    LocalMux I__10920 (
            .O(N__51769),
            .I(N__51743));
    Span4Mux_h I__10919 (
            .O(N__51766),
            .I(N__51743));
    LocalMux I__10918 (
            .O(N__51763),
            .I(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ));
    LocalMux I__10917 (
            .O(N__51760),
            .I(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ));
    LocalMux I__10916 (
            .O(N__51757),
            .I(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ));
    LocalMux I__10915 (
            .O(N__51754),
            .I(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ));
    LocalMux I__10914 (
            .O(N__51751),
            .I(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ));
    Odrv4 I__10913 (
            .O(N__51748),
            .I(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ));
    Odrv4 I__10912 (
            .O(N__51743),
            .I(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ));
    CascadeMux I__10911 (
            .O(N__51728),
            .I(N__51724));
    InMux I__10910 (
            .O(N__51727),
            .I(N__51717));
    InMux I__10909 (
            .O(N__51724),
            .I(N__51714));
    CascadeMux I__10908 (
            .O(N__51723),
            .I(N__51711));
    CascadeMux I__10907 (
            .O(N__51722),
            .I(N__51708));
    CascadeMux I__10906 (
            .O(N__51721),
            .I(N__51705));
    CascadeMux I__10905 (
            .O(N__51720),
            .I(N__51700));
    LocalMux I__10904 (
            .O(N__51717),
            .I(N__51695));
    LocalMux I__10903 (
            .O(N__51714),
            .I(N__51695));
    InMux I__10902 (
            .O(N__51711),
            .I(N__51692));
    InMux I__10901 (
            .O(N__51708),
            .I(N__51689));
    InMux I__10900 (
            .O(N__51705),
            .I(N__51686));
    InMux I__10899 (
            .O(N__51704),
            .I(N__51683));
    InMux I__10898 (
            .O(N__51703),
            .I(N__51680));
    InMux I__10897 (
            .O(N__51700),
            .I(N__51677));
    Span4Mux_v I__10896 (
            .O(N__51695),
            .I(N__51674));
    LocalMux I__10895 (
            .O(N__51692),
            .I(N__51669));
    LocalMux I__10894 (
            .O(N__51689),
            .I(N__51669));
    LocalMux I__10893 (
            .O(N__51686),
            .I(N__51660));
    LocalMux I__10892 (
            .O(N__51683),
            .I(N__51660));
    LocalMux I__10891 (
            .O(N__51680),
            .I(N__51660));
    LocalMux I__10890 (
            .O(N__51677),
            .I(N__51660));
    Span4Mux_v I__10889 (
            .O(N__51674),
            .I(N__51657));
    Span4Mux_v I__10888 (
            .O(N__51669),
            .I(N__51654));
    Span12Mux_v I__10887 (
            .O(N__51660),
            .I(N__51649));
    Sp12to4 I__10886 (
            .O(N__51657),
            .I(N__51649));
    Span4Mux_h I__10885 (
            .O(N__51654),
            .I(N__51646));
    Span12Mux_s11_h I__10884 (
            .O(N__51649),
            .I(N__51643));
    Odrv4 I__10883 (
            .O(N__51646),
            .I(\ALU.a_15_m3_sZ0Z_13 ));
    Odrv12 I__10882 (
            .O(N__51643),
            .I(\ALU.a_15_m3_sZ0Z_13 ));
    InMux I__10881 (
            .O(N__51638),
            .I(N__51629));
    InMux I__10880 (
            .O(N__51637),
            .I(N__51626));
    InMux I__10879 (
            .O(N__51636),
            .I(N__51623));
    InMux I__10878 (
            .O(N__51635),
            .I(N__51620));
    InMux I__10877 (
            .O(N__51634),
            .I(N__51617));
    InMux I__10876 (
            .O(N__51633),
            .I(N__51614));
    InMux I__10875 (
            .O(N__51632),
            .I(N__51611));
    LocalMux I__10874 (
            .O(N__51629),
            .I(N__51608));
    LocalMux I__10873 (
            .O(N__51626),
            .I(N__51605));
    LocalMux I__10872 (
            .O(N__51623),
            .I(N__51602));
    LocalMux I__10871 (
            .O(N__51620),
            .I(\ALU.mult_495_c_RNIKOB51JZ0 ));
    LocalMux I__10870 (
            .O(N__51617),
            .I(\ALU.mult_495_c_RNIKOB51JZ0 ));
    LocalMux I__10869 (
            .O(N__51614),
            .I(\ALU.mult_495_c_RNIKOB51JZ0 ));
    LocalMux I__10868 (
            .O(N__51611),
            .I(\ALU.mult_495_c_RNIKOB51JZ0 ));
    Odrv4 I__10867 (
            .O(N__51608),
            .I(\ALU.mult_495_c_RNIKOB51JZ0 ));
    Odrv4 I__10866 (
            .O(N__51605),
            .I(\ALU.mult_495_c_RNIKOB51JZ0 ));
    Odrv12 I__10865 (
            .O(N__51602),
            .I(\ALU.mult_495_c_RNIKOB51JZ0 ));
    InMux I__10864 (
            .O(N__51587),
            .I(N__51584));
    LocalMux I__10863 (
            .O(N__51584),
            .I(N__51581));
    Span4Mux_h I__10862 (
            .O(N__51581),
            .I(N__51577));
    InMux I__10861 (
            .O(N__51580),
            .I(N__51574));
    Span4Mux_h I__10860 (
            .O(N__51577),
            .I(N__51571));
    LocalMux I__10859 (
            .O(N__51574),
            .I(N__51568));
    Span4Mux_h I__10858 (
            .O(N__51571),
            .I(N__51565));
    Span12Mux_h I__10857 (
            .O(N__51568),
            .I(N__51562));
    Span4Mux_v I__10856 (
            .O(N__51565),
            .I(N__51559));
    Odrv12 I__10855 (
            .O(N__51562),
            .I(\ALU.dZ0Z_8 ));
    Odrv4 I__10854 (
            .O(N__51559),
            .I(\ALU.dZ0Z_8 ));
    CascadeMux I__10853 (
            .O(N__51554),
            .I(\ALU.c_RNIV5AOKZ0Z_13_cascade_ ));
    CascadeMux I__10852 (
            .O(N__51551),
            .I(\ALU.c_RNIO5N04A_0Z0Z_13_cascade_ ));
    InMux I__10851 (
            .O(N__51548),
            .I(N__51545));
    LocalMux I__10850 (
            .O(N__51545),
            .I(N__51542));
    Span4Mux_v I__10849 (
            .O(N__51542),
            .I(N__51538));
    InMux I__10848 (
            .O(N__51541),
            .I(N__51535));
    Span4Mux_v I__10847 (
            .O(N__51538),
            .I(N__51532));
    LocalMux I__10846 (
            .O(N__51535),
            .I(N__51529));
    Sp12to4 I__10845 (
            .O(N__51532),
            .I(N__51526));
    Span4Mux_v I__10844 (
            .O(N__51529),
            .I(N__51523));
    Span12Mux_h I__10843 (
            .O(N__51526),
            .I(N__51520));
    Odrv4 I__10842 (
            .O(N__51523),
            .I(\ALU.bZ0Z_13 ));
    Odrv12 I__10841 (
            .O(N__51520),
            .I(\ALU.bZ0Z_13 ));
    InMux I__10840 (
            .O(N__51515),
            .I(N__51512));
    LocalMux I__10839 (
            .O(N__51512),
            .I(\ALU.c_RNIV5AOKZ0Z_13 ));
    CascadeMux I__10838 (
            .O(N__51509),
            .I(N__51506));
    InMux I__10837 (
            .O(N__51506),
            .I(N__51503));
    LocalMux I__10836 (
            .O(N__51503),
            .I(N__51499));
    InMux I__10835 (
            .O(N__51502),
            .I(N__51496));
    Odrv4 I__10834 (
            .O(N__51499),
            .I(\ALU.d_RNIRFBHE9Z0Z_0 ));
    LocalMux I__10833 (
            .O(N__51496),
            .I(\ALU.d_RNIRFBHE9Z0Z_0 ));
    InMux I__10832 (
            .O(N__51491),
            .I(N__51487));
    InMux I__10831 (
            .O(N__51490),
            .I(N__51484));
    LocalMux I__10830 (
            .O(N__51487),
            .I(N__51481));
    LocalMux I__10829 (
            .O(N__51484),
            .I(N__51478));
    Span4Mux_h I__10828 (
            .O(N__51481),
            .I(N__51475));
    Span12Mux_v I__10827 (
            .O(N__51478),
            .I(N__51472));
    Span4Mux_v I__10826 (
            .O(N__51475),
            .I(N__51469));
    Span12Mux_h I__10825 (
            .O(N__51472),
            .I(N__51466));
    Odrv4 I__10824 (
            .O(N__51469),
            .I(\ALU.log_1_4 ));
    Odrv12 I__10823 (
            .O(N__51466),
            .I(\ALU.log_1_4 ));
    CascadeMux I__10822 (
            .O(N__51461),
            .I(\ALU.N_16_0_cascade_ ));
    InMux I__10821 (
            .O(N__51458),
            .I(N__51455));
    LocalMux I__10820 (
            .O(N__51455),
            .I(N__51452));
    Span4Mux_h I__10819 (
            .O(N__51452),
            .I(N__51449));
    Span4Mux_h I__10818 (
            .O(N__51449),
            .I(N__51446));
    Odrv4 I__10817 (
            .O(N__51446),
            .I(\ALU.status_8_8_0 ));
    InMux I__10816 (
            .O(N__51443),
            .I(N__51440));
    LocalMux I__10815 (
            .O(N__51440),
            .I(\ALU.log_1_9 ));
    InMux I__10814 (
            .O(N__51437),
            .I(N__51434));
    LocalMux I__10813 (
            .O(N__51434),
            .I(N__51431));
    Span4Mux_h I__10812 (
            .O(N__51431),
            .I(N__51428));
    Span4Mux_v I__10811 (
            .O(N__51428),
            .I(N__51425));
    Odrv4 I__10810 (
            .O(N__51425),
            .I(\ALU.d_RNI7KS2IZ0Z_9 ));
    CascadeMux I__10809 (
            .O(N__51422),
            .I(N__51418));
    CascadeMux I__10808 (
            .O(N__51421),
            .I(N__51415));
    InMux I__10807 (
            .O(N__51418),
            .I(N__51412));
    InMux I__10806 (
            .O(N__51415),
            .I(N__51409));
    LocalMux I__10805 (
            .O(N__51412),
            .I(N__51406));
    LocalMux I__10804 (
            .O(N__51409),
            .I(N__51403));
    Span4Mux_h I__10803 (
            .O(N__51406),
            .I(N__51400));
    Span4Mux_v I__10802 (
            .O(N__51403),
            .I(N__51397));
    Span4Mux_h I__10801 (
            .O(N__51400),
            .I(N__51394));
    Span4Mux_h I__10800 (
            .O(N__51397),
            .I(N__51391));
    Span4Mux_v I__10799 (
            .O(N__51394),
            .I(N__51388));
    Span4Mux_h I__10798 (
            .O(N__51391),
            .I(N__51385));
    Span4Mux_h I__10797 (
            .O(N__51388),
            .I(N__51382));
    Odrv4 I__10796 (
            .O(N__51385),
            .I(\ALU.eZ0Z_12 ));
    Odrv4 I__10795 (
            .O(N__51382),
            .I(\ALU.eZ0Z_12 ));
    CascadeMux I__10794 (
            .O(N__51377),
            .I(\PROM.ROMDATA.m58_cascade_ ));
    InMux I__10793 (
            .O(N__51374),
            .I(N__51371));
    LocalMux I__10792 (
            .O(N__51371),
            .I(\PROM.ROMDATA.m64_am ));
    InMux I__10791 (
            .O(N__51368),
            .I(N__51365));
    LocalMux I__10790 (
            .O(N__51365),
            .I(N__51362));
    Odrv4 I__10789 (
            .O(N__51362),
            .I(\PROM.ROMDATA.m45 ));
    InMux I__10788 (
            .O(N__51359),
            .I(N__51356));
    LocalMux I__10787 (
            .O(N__51356),
            .I(N__51353));
    Span4Mux_h I__10786 (
            .O(N__51353),
            .I(N__51350));
    Span4Mux_v I__10785 (
            .O(N__51350),
            .I(N__51347));
    Odrv4 I__10784 (
            .O(N__51347),
            .I(\ALU.log_1_7 ));
    InMux I__10783 (
            .O(N__51344),
            .I(N__51341));
    LocalMux I__10782 (
            .O(N__51341),
            .I(N__51338));
    Span4Mux_h I__10781 (
            .O(N__51338),
            .I(N__51335));
    Span4Mux_h I__10780 (
            .O(N__51335),
            .I(N__51331));
    InMux I__10779 (
            .O(N__51334),
            .I(N__51328));
    Odrv4 I__10778 (
            .O(N__51331),
            .I(\ALU.log_1_5 ));
    LocalMux I__10777 (
            .O(N__51328),
            .I(\ALU.log_1_5 ));
    CascadeMux I__10776 (
            .O(N__51323),
            .I(N__51319));
    InMux I__10775 (
            .O(N__51322),
            .I(N__51316));
    InMux I__10774 (
            .O(N__51319),
            .I(N__51313));
    LocalMux I__10773 (
            .O(N__51316),
            .I(N__51310));
    LocalMux I__10772 (
            .O(N__51313),
            .I(N__51307));
    Span4Mux_v I__10771 (
            .O(N__51310),
            .I(N__51304));
    Span4Mux_h I__10770 (
            .O(N__51307),
            .I(N__51301));
    Odrv4 I__10769 (
            .O(N__51304),
            .I(\ALU.log_1_11 ));
    Odrv4 I__10768 (
            .O(N__51301),
            .I(\ALU.log_1_11 ));
    InMux I__10767 (
            .O(N__51296),
            .I(N__51292));
    InMux I__10766 (
            .O(N__51295),
            .I(N__51289));
    LocalMux I__10765 (
            .O(N__51292),
            .I(N__51286));
    LocalMux I__10764 (
            .O(N__51289),
            .I(N__51283));
    Span4Mux_v I__10763 (
            .O(N__51286),
            .I(N__51280));
    Span4Mux_v I__10762 (
            .O(N__51283),
            .I(N__51277));
    Span4Mux_v I__10761 (
            .O(N__51280),
            .I(N__51272));
    Span4Mux_v I__10760 (
            .O(N__51277),
            .I(N__51272));
    Sp12to4 I__10759 (
            .O(N__51272),
            .I(N__51269));
    Span12Mux_h I__10758 (
            .O(N__51269),
            .I(N__51266));
    Odrv12 I__10757 (
            .O(N__51266),
            .I(\ALU.log_1_10 ));
    InMux I__10756 (
            .O(N__51263),
            .I(N__51259));
    InMux I__10755 (
            .O(N__51262),
            .I(N__51256));
    LocalMux I__10754 (
            .O(N__51259),
            .I(N__51253));
    LocalMux I__10753 (
            .O(N__51256),
            .I(N__51248));
    Span12Mux_v I__10752 (
            .O(N__51253),
            .I(N__51248));
    Span12Mux_h I__10751 (
            .O(N__51248),
            .I(N__51245));
    Odrv12 I__10750 (
            .O(N__51245),
            .I(\ALU.N_22_0 ));
    InMux I__10749 (
            .O(N__51242),
            .I(N__51239));
    LocalMux I__10748 (
            .O(N__51239),
            .I(N__51235));
    InMux I__10747 (
            .O(N__51238),
            .I(N__51232));
    Span4Mux_h I__10746 (
            .O(N__51235),
            .I(N__51229));
    LocalMux I__10745 (
            .O(N__51232),
            .I(N__51226));
    Span4Mux_v I__10744 (
            .O(N__51229),
            .I(N__51223));
    Span4Mux_v I__10743 (
            .O(N__51226),
            .I(N__51220));
    Span4Mux_h I__10742 (
            .O(N__51223),
            .I(N__51217));
    Span4Mux_h I__10741 (
            .O(N__51220),
            .I(N__51214));
    Span4Mux_v I__10740 (
            .O(N__51217),
            .I(N__51211));
    Odrv4 I__10739 (
            .O(N__51214),
            .I(\ALU.N_20_0 ));
    Odrv4 I__10738 (
            .O(N__51211),
            .I(\ALU.N_20_0 ));
    CascadeMux I__10737 (
            .O(N__51206),
            .I(\ALU.status_8_10_0_cascade_ ));
    InMux I__10736 (
            .O(N__51203),
            .I(N__51200));
    LocalMux I__10735 (
            .O(N__51200),
            .I(N__51197));
    Span4Mux_h I__10734 (
            .O(N__51197),
            .I(N__51194));
    Span4Mux_h I__10733 (
            .O(N__51194),
            .I(N__51191));
    Odrv4 I__10732 (
            .O(N__51191),
            .I(\ALU.status_8_13_0 ));
    InMux I__10731 (
            .O(N__51188),
            .I(N__51185));
    LocalMux I__10730 (
            .O(N__51185),
            .I(\ALU.status_8_3_1_0 ));
    CascadeMux I__10729 (
            .O(N__51182),
            .I(\ALU.log_1_15_cascade_ ));
    InMux I__10728 (
            .O(N__51179),
            .I(N__51176));
    LocalMux I__10727 (
            .O(N__51176),
            .I(\ALU.status_8_13_1_0 ));
    CascadeMux I__10726 (
            .O(N__51173),
            .I(\PROM.ROMDATA.m191_cascade_ ));
    InMux I__10725 (
            .O(N__51170),
            .I(N__51167));
    LocalMux I__10724 (
            .O(N__51167),
            .I(\PROM.ROMDATA.m193 ));
    InMux I__10723 (
            .O(N__51164),
            .I(N__51161));
    LocalMux I__10722 (
            .O(N__51161),
            .I(\PROM.ROMDATA.m195_bm ));
    InMux I__10721 (
            .O(N__51158),
            .I(N__51155));
    LocalMux I__10720 (
            .O(N__51155),
            .I(N__51152));
    Span4Mux_v I__10719 (
            .O(N__51152),
            .I(N__51149));
    Span4Mux_h I__10718 (
            .O(N__51149),
            .I(N__51145));
    InMux I__10717 (
            .O(N__51148),
            .I(N__51142));
    Span4Mux_h I__10716 (
            .O(N__51145),
            .I(N__51139));
    LocalMux I__10715 (
            .O(N__51142),
            .I(N__51136));
    Span4Mux_v I__10714 (
            .O(N__51139),
            .I(N__51133));
    Span4Mux_h I__10713 (
            .O(N__51136),
            .I(N__51130));
    Odrv4 I__10712 (
            .O(N__51133),
            .I(\CONTROL.programCounter_1_3 ));
    Odrv4 I__10711 (
            .O(N__51130),
            .I(\CONTROL.programCounter_1_3 ));
    InMux I__10710 (
            .O(N__51125),
            .I(N__51122));
    LocalMux I__10709 (
            .O(N__51122),
            .I(N__51118));
    InMux I__10708 (
            .O(N__51121),
            .I(N__51115));
    Span4Mux_h I__10707 (
            .O(N__51118),
            .I(N__51110));
    LocalMux I__10706 (
            .O(N__51115),
            .I(N__51110));
    Odrv4 I__10705 (
            .O(N__51110),
            .I(\CONTROL.programCounter_1_reto_3 ));
    InMux I__10704 (
            .O(N__51107),
            .I(N__51104));
    LocalMux I__10703 (
            .O(N__51104),
            .I(N__51101));
    Odrv12 I__10702 (
            .O(N__51101),
            .I(\PROM.ROMDATA.m92_am ));
    CascadeMux I__10701 (
            .O(N__51098),
            .I(\PROM.ROMDATA.m62_cascade_ ));
    InMux I__10700 (
            .O(N__51095),
            .I(N__51092));
    LocalMux I__10699 (
            .O(N__51092),
            .I(N__51089));
    Odrv4 I__10698 (
            .O(N__51089),
            .I(\PROM.ROMDATA.m53_am ));
    CascadeMux I__10697 (
            .O(N__51086),
            .I(N__51083));
    InMux I__10696 (
            .O(N__51083),
            .I(N__51080));
    LocalMux I__10695 (
            .O(N__51080),
            .I(N__51077));
    Odrv4 I__10694 (
            .O(N__51077),
            .I(\PROM.ROMDATA.m53_bm ));
    InMux I__10693 (
            .O(N__51074),
            .I(N__51071));
    LocalMux I__10692 (
            .O(N__51071),
            .I(\PROM.ROMDATA.m64_bm ));
    CascadeMux I__10691 (
            .O(N__51068),
            .I(\PROM.ROMDATA.m65_ns_1_cascade_ ));
    InMux I__10690 (
            .O(N__51065),
            .I(N__51059));
    InMux I__10689 (
            .O(N__51064),
            .I(N__51059));
    LocalMux I__10688 (
            .O(N__51059),
            .I(N__51056));
    Span4Mux_h I__10687 (
            .O(N__51056),
            .I(N__51053));
    Odrv4 I__10686 (
            .O(N__51053),
            .I(m65_ns));
    CascadeMux I__10685 (
            .O(N__51050),
            .I(\PROM.ROMDATA.m80_am_cascade_ ));
    InMux I__10684 (
            .O(N__51047),
            .I(N__51044));
    LocalMux I__10683 (
            .O(N__51044),
            .I(N__51041));
    Span4Mux_v I__10682 (
            .O(N__51041),
            .I(N__51038));
    Odrv4 I__10681 (
            .O(N__51038),
            .I(\PROM.ROMDATA.m93_ns_1 ));
    InMux I__10680 (
            .O(N__51035),
            .I(N__51032));
    LocalMux I__10679 (
            .O(N__51032),
            .I(\CONTROL.programCounter_ret_1_RNIJ88IZ0Z_2 ));
    InMux I__10678 (
            .O(N__51029),
            .I(N__51026));
    LocalMux I__10677 (
            .O(N__51026),
            .I(\CONTROL.programCounter_ret_19_RNICM8JZ0Z_2 ));
    CascadeMux I__10676 (
            .O(N__51023),
            .I(progRomAddress_2_cascade_));
    InMux I__10675 (
            .O(N__51020),
            .I(N__51017));
    LocalMux I__10674 (
            .O(N__51017),
            .I(N__51014));
    Span4Mux_v I__10673 (
            .O(N__51014),
            .I(N__51011));
    Odrv4 I__10672 (
            .O(N__51011),
            .I(\PROM.ROMDATA.m195_am ));
    CascadeMux I__10671 (
            .O(N__51008),
            .I(\PROM.ROMDATA.m196_ns_1_cascade_ ));
    InMux I__10670 (
            .O(N__51005),
            .I(N__51002));
    LocalMux I__10669 (
            .O(N__51002),
            .I(N__50999));
    Odrv4 I__10668 (
            .O(N__50999),
            .I(\PROM.ROMDATA.m179 ));
    InMux I__10667 (
            .O(N__50996),
            .I(N__50993));
    LocalMux I__10666 (
            .O(N__50993),
            .I(\PROM.ROMDATA.m185_am ));
    InMux I__10665 (
            .O(N__50990),
            .I(N__50987));
    LocalMux I__10664 (
            .O(N__50987),
            .I(N__50983));
    InMux I__10663 (
            .O(N__50986),
            .I(N__50980));
    Span4Mux_h I__10662 (
            .O(N__50983),
            .I(N__50977));
    LocalMux I__10661 (
            .O(N__50980),
            .I(N__50974));
    Odrv4 I__10660 (
            .O(N__50977),
            .I(\CONTROL.dout_reto_0 ));
    Odrv4 I__10659 (
            .O(N__50974),
            .I(\CONTROL.dout_reto_0 ));
    InMux I__10658 (
            .O(N__50969),
            .I(N__50966));
    LocalMux I__10657 (
            .O(N__50966),
            .I(N__50963));
    Span4Mux_h I__10656 (
            .O(N__50963),
            .I(N__50959));
    InMux I__10655 (
            .O(N__50962),
            .I(N__50956));
    Sp12to4 I__10654 (
            .O(N__50959),
            .I(N__50952));
    LocalMux I__10653 (
            .O(N__50956),
            .I(N__50949));
    InMux I__10652 (
            .O(N__50955),
            .I(N__50944));
    Span12Mux_v I__10651 (
            .O(N__50952),
            .I(N__50941));
    Span4Mux_h I__10650 (
            .O(N__50949),
            .I(N__50938));
    InMux I__10649 (
            .O(N__50948),
            .I(N__50935));
    InMux I__10648 (
            .O(N__50947),
            .I(N__50932));
    LocalMux I__10647 (
            .O(N__50944),
            .I(CONTROL_addrstack_reto_0));
    Odrv12 I__10646 (
            .O(N__50941),
            .I(CONTROL_addrstack_reto_0));
    Odrv4 I__10645 (
            .O(N__50938),
            .I(CONTROL_addrstack_reto_0));
    LocalMux I__10644 (
            .O(N__50935),
            .I(CONTROL_addrstack_reto_0));
    LocalMux I__10643 (
            .O(N__50932),
            .I(CONTROL_addrstack_reto_0));
    CascadeMux I__10642 (
            .O(N__50921),
            .I(N__50918));
    InMux I__10641 (
            .O(N__50918),
            .I(N__50915));
    LocalMux I__10640 (
            .O(N__50915),
            .I(N__50912));
    Span4Mux_v I__10639 (
            .O(N__50912),
            .I(N__50909));
    Odrv4 I__10638 (
            .O(N__50909),
            .I(\PROM.ROMDATA.m248_ns_1 ));
    InMux I__10637 (
            .O(N__50906),
            .I(N__50900));
    InMux I__10636 (
            .O(N__50905),
            .I(N__50893));
    InMux I__10635 (
            .O(N__50904),
            .I(N__50893));
    InMux I__10634 (
            .O(N__50903),
            .I(N__50890));
    LocalMux I__10633 (
            .O(N__50900),
            .I(N__50887));
    InMux I__10632 (
            .O(N__50899),
            .I(N__50884));
    InMux I__10631 (
            .O(N__50898),
            .I(N__50881));
    LocalMux I__10630 (
            .O(N__50893),
            .I(N__50876));
    LocalMux I__10629 (
            .O(N__50890),
            .I(N__50876));
    Span4Mux_v I__10628 (
            .O(N__50887),
            .I(N__50873));
    LocalMux I__10627 (
            .O(N__50884),
            .I(N__50866));
    LocalMux I__10626 (
            .O(N__50881),
            .I(N__50866));
    Span4Mux_h I__10625 (
            .O(N__50876),
            .I(N__50863));
    Span4Mux_h I__10624 (
            .O(N__50873),
            .I(N__50860));
    InMux I__10623 (
            .O(N__50872),
            .I(N__50855));
    InMux I__10622 (
            .O(N__50871),
            .I(N__50855));
    Span4Mux_v I__10621 (
            .O(N__50866),
            .I(N__50850));
    Span4Mux_h I__10620 (
            .O(N__50863),
            .I(N__50850));
    Odrv4 I__10619 (
            .O(N__50860),
            .I(\CONTROL.incrementZ0Z_0 ));
    LocalMux I__10618 (
            .O(N__50855),
            .I(\CONTROL.incrementZ0Z_0 ));
    Odrv4 I__10617 (
            .O(N__50850),
            .I(\CONTROL.incrementZ0Z_0 ));
    CascadeMux I__10616 (
            .O(N__50843),
            .I(N__50838));
    CascadeMux I__10615 (
            .O(N__50842),
            .I(N__50831));
    InMux I__10614 (
            .O(N__50841),
            .I(N__50827));
    InMux I__10613 (
            .O(N__50838),
            .I(N__50822));
    InMux I__10612 (
            .O(N__50837),
            .I(N__50822));
    InMux I__10611 (
            .O(N__50836),
            .I(N__50819));
    InMux I__10610 (
            .O(N__50835),
            .I(N__50816));
    InMux I__10609 (
            .O(N__50834),
            .I(N__50813));
    InMux I__10608 (
            .O(N__50831),
            .I(N__50808));
    InMux I__10607 (
            .O(N__50830),
            .I(N__50808));
    LocalMux I__10606 (
            .O(N__50827),
            .I(N__50805));
    LocalMux I__10605 (
            .O(N__50822),
            .I(N__50800));
    LocalMux I__10604 (
            .O(N__50819),
            .I(N__50800));
    LocalMux I__10603 (
            .O(N__50816),
            .I(N__50797));
    LocalMux I__10602 (
            .O(N__50813),
            .I(N__50794));
    LocalMux I__10601 (
            .O(N__50808),
            .I(N__50791));
    Span4Mux_v I__10600 (
            .O(N__50805),
            .I(N__50788));
    Span4Mux_v I__10599 (
            .O(N__50800),
            .I(N__50785));
    Span4Mux_v I__10598 (
            .O(N__50797),
            .I(N__50782));
    Span4Mux_h I__10597 (
            .O(N__50794),
            .I(N__50775));
    Span4Mux_v I__10596 (
            .O(N__50791),
            .I(N__50775));
    Span4Mux_h I__10595 (
            .O(N__50788),
            .I(N__50775));
    Span4Mux_h I__10594 (
            .O(N__50785),
            .I(N__50772));
    Span4Mux_h I__10593 (
            .O(N__50782),
            .I(N__50767));
    Span4Mux_v I__10592 (
            .O(N__50775),
            .I(N__50767));
    Span4Mux_h I__10591 (
            .O(N__50772),
            .I(N__50764));
    Odrv4 I__10590 (
            .O(N__50767),
            .I(\CONTROL.incrementZ0Z_1 ));
    Odrv4 I__10589 (
            .O(N__50764),
            .I(\CONTROL.incrementZ0Z_1 ));
    InMux I__10588 (
            .O(N__50759),
            .I(N__50756));
    LocalMux I__10587 (
            .O(N__50756),
            .I(N__50753));
    Span4Mux_h I__10586 (
            .O(N__50753),
            .I(N__50750));
    Odrv4 I__10585 (
            .O(N__50750),
            .I(\PROM.ROMDATA.m284_1 ));
    InMux I__10584 (
            .O(N__50747),
            .I(N__50744));
    LocalMux I__10583 (
            .O(N__50744),
            .I(\CONTROL.programCounter_ret_19_RNI8I8JZ0Z_0 ));
    InMux I__10582 (
            .O(N__50741),
            .I(N__50738));
    LocalMux I__10581 (
            .O(N__50738),
            .I(\CONTROL.programCounter_ret_1_RNIF48IZ0Z_0 ));
    CascadeMux I__10580 (
            .O(N__50735),
            .I(progRomAddress_0_cascade_));
    CascadeMux I__10579 (
            .O(N__50732),
            .I(\PROM.ROMDATA.m72_cascade_ ));
    InMux I__10578 (
            .O(N__50729),
            .I(N__50726));
    LocalMux I__10577 (
            .O(N__50726),
            .I(\PROM.ROMDATA.m74 ));
    CascadeMux I__10576 (
            .O(N__50723),
            .I(\PROM.ROMDATA.m169_cascade_ ));
    InMux I__10575 (
            .O(N__50720),
            .I(N__50717));
    LocalMux I__10574 (
            .O(N__50717),
            .I(N__50714));
    Span4Mux_h I__10573 (
            .O(N__50714),
            .I(N__50710));
    InMux I__10572 (
            .O(N__50713),
            .I(N__50707));
    Span4Mux_h I__10571 (
            .O(N__50710),
            .I(N__50704));
    LocalMux I__10570 (
            .O(N__50707),
            .I(N__50701));
    Odrv4 I__10569 (
            .O(N__50704),
            .I(\PROM.ROMDATA.m270_am ));
    Odrv12 I__10568 (
            .O(N__50701),
            .I(\PROM.ROMDATA.m270_am ));
    CascadeMux I__10567 (
            .O(N__50696),
            .I(\PROM.ROMDATA.m13_cascade_ ));
    InMux I__10566 (
            .O(N__50693),
            .I(N__50690));
    LocalMux I__10565 (
            .O(N__50690),
            .I(\PROM.ROMDATA.m188 ));
    CascadeMux I__10564 (
            .O(N__50687),
            .I(N__50684));
    InMux I__10563 (
            .O(N__50684),
            .I(N__50681));
    LocalMux I__10562 (
            .O(N__50681),
            .I(\PROM.ROMDATA.m13 ));
    InMux I__10561 (
            .O(N__50678),
            .I(N__50675));
    LocalMux I__10560 (
            .O(N__50675),
            .I(\PROM.ROMDATA.m263 ));
    InMux I__10559 (
            .O(N__50672),
            .I(N__50669));
    LocalMux I__10558 (
            .O(N__50669),
            .I(N__50666));
    Span4Mux_v I__10557 (
            .O(N__50666),
            .I(N__50663));
    Span4Mux_h I__10556 (
            .O(N__50663),
            .I(N__50659));
    InMux I__10555 (
            .O(N__50662),
            .I(N__50656));
    Odrv4 I__10554 (
            .O(N__50659),
            .I(\CONTROL.ctrlOut_1 ));
    LocalMux I__10553 (
            .O(N__50656),
            .I(\CONTROL.ctrlOut_1 ));
    CascadeMux I__10552 (
            .O(N__50651),
            .I(\PROM.ROMDATA.m150_cascade_ ));
    CascadeMux I__10551 (
            .O(N__50648),
            .I(\PROM.ROMDATA.m228_am_cascade_ ));
    CascadeMux I__10550 (
            .O(N__50645),
            .I(N__50642));
    InMux I__10549 (
            .O(N__50642),
            .I(N__50639));
    LocalMux I__10548 (
            .O(N__50639),
            .I(N__50636));
    Odrv4 I__10547 (
            .O(N__50636),
            .I(\PROM.ROMDATA.m25 ));
    InMux I__10546 (
            .O(N__50633),
            .I(N__50630));
    LocalMux I__10545 (
            .O(N__50630),
            .I(N__50627));
    Span4Mux_v I__10544 (
            .O(N__50627),
            .I(N__50624));
    Odrv4 I__10543 (
            .O(N__50624),
            .I(\PROM.ROMDATA.m280 ));
    CascadeMux I__10542 (
            .O(N__50621),
            .I(N__50617));
    InMux I__10541 (
            .O(N__50620),
            .I(N__50612));
    InMux I__10540 (
            .O(N__50617),
            .I(N__50612));
    LocalMux I__10539 (
            .O(N__50612),
            .I(N__50609));
    Span4Mux_v I__10538 (
            .O(N__50609),
            .I(N__50606));
    Span4Mux_h I__10537 (
            .O(N__50606),
            .I(N__50603));
    Span4Mux_h I__10536 (
            .O(N__50603),
            .I(N__50600));
    Span4Mux_h I__10535 (
            .O(N__50600),
            .I(N__50597));
    Span4Mux_v I__10534 (
            .O(N__50597),
            .I(N__50594));
    Odrv4 I__10533 (
            .O(N__50594),
            .I(\PROM.ROMDATA.m438 ));
    InMux I__10532 (
            .O(N__50591),
            .I(N__50587));
    InMux I__10531 (
            .O(N__50590),
            .I(N__50584));
    LocalMux I__10530 (
            .O(N__50587),
            .I(\PROM.ROMDATA.m173 ));
    LocalMux I__10529 (
            .O(N__50584),
            .I(\PROM.ROMDATA.m173 ));
    InMux I__10528 (
            .O(N__50579),
            .I(N__50576));
    LocalMux I__10527 (
            .O(N__50576),
            .I(N__50573));
    Span4Mux_v I__10526 (
            .O(N__50573),
            .I(N__50569));
    InMux I__10525 (
            .O(N__50572),
            .I(N__50566));
    Odrv4 I__10524 (
            .O(N__50569),
            .I(\PROM.ROMDATA.m23 ));
    LocalMux I__10523 (
            .O(N__50566),
            .I(\PROM.ROMDATA.m23 ));
    InMux I__10522 (
            .O(N__50561),
            .I(N__50558));
    LocalMux I__10521 (
            .O(N__50558),
            .I(N__50555));
    Span4Mux_v I__10520 (
            .O(N__50555),
            .I(N__50552));
    Span4Mux_h I__10519 (
            .O(N__50552),
            .I(N__50549));
    Span4Mux_h I__10518 (
            .O(N__50549),
            .I(N__50546));
    Odrv4 I__10517 (
            .O(N__50546),
            .I(PROM_ROMDATA_dintern_31_0__g1));
    CascadeMux I__10516 (
            .O(N__50543),
            .I(N__50538));
    InMux I__10515 (
            .O(N__50542),
            .I(N__50532));
    InMux I__10514 (
            .O(N__50541),
            .I(N__50532));
    InMux I__10513 (
            .O(N__50538),
            .I(N__50527));
    InMux I__10512 (
            .O(N__50537),
            .I(N__50527));
    LocalMux I__10511 (
            .O(N__50532),
            .I(N__50524));
    LocalMux I__10510 (
            .O(N__50527),
            .I(N__50521));
    Odrv4 I__10509 (
            .O(N__50524),
            .I(\ALU.a_15_m2_d_d_sZ0Z_0 ));
    Odrv4 I__10508 (
            .O(N__50521),
            .I(\ALU.a_15_m2_d_d_sZ0Z_0 ));
    CascadeMux I__10507 (
            .O(N__50516),
            .I(bus_15_cascade_));
    InMux I__10506 (
            .O(N__50513),
            .I(N__50507));
    InMux I__10505 (
            .O(N__50512),
            .I(N__50507));
    LocalMux I__10504 (
            .O(N__50507),
            .I(\ALU.c_RNIJI6SHZ0Z_15 ));
    InMux I__10503 (
            .O(N__50504),
            .I(N__50501));
    LocalMux I__10502 (
            .O(N__50501),
            .I(\ALU.c_RNID85GQZ0Z_15 ));
    CascadeMux I__10501 (
            .O(N__50498),
            .I(\PROM.ROMDATA.m248_ns_cascade_ ));
    CascadeMux I__10500 (
            .O(N__50495),
            .I(N__50491));
    CascadeMux I__10499 (
            .O(N__50494),
            .I(N__50488));
    InMux I__10498 (
            .O(N__50491),
            .I(N__50477));
    InMux I__10497 (
            .O(N__50488),
            .I(N__50477));
    InMux I__10496 (
            .O(N__50487),
            .I(N__50477));
    InMux I__10495 (
            .O(N__50486),
            .I(N__50477));
    LocalMux I__10494 (
            .O(N__50477),
            .I(N__50474));
    Span4Mux_v I__10493 (
            .O(N__50474),
            .I(N__50471));
    Span4Mux_h I__10492 (
            .O(N__50471),
            .I(N__50467));
    InMux I__10491 (
            .O(N__50470),
            .I(N__50464));
    Span4Mux_v I__10490 (
            .O(N__50467),
            .I(N__50461));
    LocalMux I__10489 (
            .O(N__50464),
            .I(N__50458));
    Span4Mux_h I__10488 (
            .O(N__50461),
            .I(N__50455));
    Span4Mux_h I__10487 (
            .O(N__50458),
            .I(N__50452));
    Odrv4 I__10486 (
            .O(N__50455),
            .I(\PROM.ROMDATA.m249 ));
    Odrv4 I__10485 (
            .O(N__50452),
            .I(\PROM.ROMDATA.m249 ));
    InMux I__10484 (
            .O(N__50447),
            .I(N__50444));
    LocalMux I__10483 (
            .O(N__50444),
            .I(N__50441));
    Odrv4 I__10482 (
            .O(N__50441),
            .I(\PROM.ROMDATA.m359 ));
    InMux I__10481 (
            .O(N__50438),
            .I(N__50435));
    LocalMux I__10480 (
            .O(N__50435),
            .I(N__50432));
    Span4Mux_v I__10479 (
            .O(N__50432),
            .I(N__50427));
    InMux I__10478 (
            .O(N__50431),
            .I(N__50422));
    InMux I__10477 (
            .O(N__50430),
            .I(N__50422));
    Span4Mux_v I__10476 (
            .O(N__50427),
            .I(N__50417));
    LocalMux I__10475 (
            .O(N__50422),
            .I(N__50417));
    Span4Mux_h I__10474 (
            .O(N__50417),
            .I(N__50414));
    Span4Mux_h I__10473 (
            .O(N__50414),
            .I(N__50411));
    Span4Mux_h I__10472 (
            .O(N__50411),
            .I(N__50408));
    Odrv4 I__10471 (
            .O(N__50408),
            .I(g_8));
    CascadeMux I__10470 (
            .O(N__50405),
            .I(N__50401));
    CascadeMux I__10469 (
            .O(N__50404),
            .I(N__50397));
    InMux I__10468 (
            .O(N__50401),
            .I(N__50394));
    InMux I__10467 (
            .O(N__50400),
            .I(N__50389));
    InMux I__10466 (
            .O(N__50397),
            .I(N__50389));
    LocalMux I__10465 (
            .O(N__50394),
            .I(N__50386));
    LocalMux I__10464 (
            .O(N__50389),
            .I(N__50383));
    Span4Mux_v I__10463 (
            .O(N__50386),
            .I(N__50380));
    Span4Mux_v I__10462 (
            .O(N__50383),
            .I(N__50377));
    Span4Mux_h I__10461 (
            .O(N__50380),
            .I(N__50374));
    Span4Mux_h I__10460 (
            .O(N__50377),
            .I(N__50371));
    Span4Mux_h I__10459 (
            .O(N__50374),
            .I(N__50368));
    Span4Mux_h I__10458 (
            .O(N__50371),
            .I(N__50365));
    Span4Mux_v I__10457 (
            .O(N__50368),
            .I(N__50362));
    Span4Mux_h I__10456 (
            .O(N__50365),
            .I(N__50359));
    Odrv4 I__10455 (
            .O(N__50362),
            .I(g_15));
    Odrv4 I__10454 (
            .O(N__50359),
            .I(g_15));
    CascadeMux I__10453 (
            .O(N__50354),
            .I(\ALU.c_RNID85GQ_0Z0Z_15_cascade_ ));
    InMux I__10452 (
            .O(N__50351),
            .I(N__50348));
    LocalMux I__10451 (
            .O(N__50348),
            .I(N__50345));
    Odrv12 I__10450 (
            .O(N__50345),
            .I(\ALU.c_RNI9DCRE2Z0Z_15 ));
    InMux I__10449 (
            .O(N__50342),
            .I(N__50338));
    InMux I__10448 (
            .O(N__50341),
            .I(N__50334));
    LocalMux I__10447 (
            .O(N__50338),
            .I(N__50331));
    InMux I__10446 (
            .O(N__50337),
            .I(N__50328));
    LocalMux I__10445 (
            .O(N__50334),
            .I(N__50321));
    Span4Mux_v I__10444 (
            .O(N__50331),
            .I(N__50318));
    LocalMux I__10443 (
            .O(N__50328),
            .I(N__50315));
    InMux I__10442 (
            .O(N__50327),
            .I(N__50312));
    InMux I__10441 (
            .O(N__50326),
            .I(N__50309));
    InMux I__10440 (
            .O(N__50325),
            .I(N__50306));
    InMux I__10439 (
            .O(N__50324),
            .I(N__50302));
    Span4Mux_v I__10438 (
            .O(N__50321),
            .I(N__50299));
    Span4Mux_h I__10437 (
            .O(N__50318),
            .I(N__50293));
    Span4Mux_v I__10436 (
            .O(N__50315),
            .I(N__50293));
    LocalMux I__10435 (
            .O(N__50312),
            .I(N__50290));
    LocalMux I__10434 (
            .O(N__50309),
            .I(N__50287));
    LocalMux I__10433 (
            .O(N__50306),
            .I(N__50284));
    InMux I__10432 (
            .O(N__50305),
            .I(N__50281));
    LocalMux I__10431 (
            .O(N__50302),
            .I(N__50277));
    Span4Mux_v I__10430 (
            .O(N__50299),
            .I(N__50274));
    InMux I__10429 (
            .O(N__50298),
            .I(N__50271));
    Span4Mux_h I__10428 (
            .O(N__50293),
            .I(N__50266));
    Span4Mux_v I__10427 (
            .O(N__50290),
            .I(N__50266));
    Span12Mux_h I__10426 (
            .O(N__50287),
            .I(N__50259));
    Sp12to4 I__10425 (
            .O(N__50284),
            .I(N__50259));
    LocalMux I__10424 (
            .O(N__50281),
            .I(N__50259));
    InMux I__10423 (
            .O(N__50280),
            .I(N__50256));
    Odrv12 I__10422 (
            .O(N__50277),
            .I(DROM_ROMDATA_dintern_adflt));
    Odrv4 I__10421 (
            .O(N__50274),
            .I(DROM_ROMDATA_dintern_adflt));
    LocalMux I__10420 (
            .O(N__50271),
            .I(DROM_ROMDATA_dintern_adflt));
    Odrv4 I__10419 (
            .O(N__50266),
            .I(DROM_ROMDATA_dintern_adflt));
    Odrv12 I__10418 (
            .O(N__50259),
            .I(DROM_ROMDATA_dintern_adflt));
    LocalMux I__10417 (
            .O(N__50256),
            .I(DROM_ROMDATA_dintern_adflt));
    CascadeMux I__10416 (
            .O(N__50243),
            .I(N__50240));
    InMux I__10415 (
            .O(N__50240),
            .I(N__50237));
    LocalMux I__10414 (
            .O(N__50237),
            .I(N__50234));
    Span12Mux_v I__10413 (
            .O(N__50234),
            .I(N__50231));
    Span12Mux_h I__10412 (
            .O(N__50231),
            .I(N__50228));
    Odrv12 I__10411 (
            .O(N__50228),
            .I(DROM_ROMDATA_dintern_15ro));
    InMux I__10410 (
            .O(N__50225),
            .I(N__50204));
    InMux I__10409 (
            .O(N__50224),
            .I(N__50204));
    InMux I__10408 (
            .O(N__50223),
            .I(N__50204));
    InMux I__10407 (
            .O(N__50222),
            .I(N__50204));
    InMux I__10406 (
            .O(N__50221),
            .I(N__50194));
    InMux I__10405 (
            .O(N__50220),
            .I(N__50191));
    InMux I__10404 (
            .O(N__50219),
            .I(N__50187));
    InMux I__10403 (
            .O(N__50218),
            .I(N__50183));
    InMux I__10402 (
            .O(N__50217),
            .I(N__50178));
    InMux I__10401 (
            .O(N__50216),
            .I(N__50178));
    InMux I__10400 (
            .O(N__50215),
            .I(N__50175));
    InMux I__10399 (
            .O(N__50214),
            .I(N__50172));
    InMux I__10398 (
            .O(N__50213),
            .I(N__50169));
    LocalMux I__10397 (
            .O(N__50204),
            .I(N__50165));
    InMux I__10396 (
            .O(N__50203),
            .I(N__50158));
    InMux I__10395 (
            .O(N__50202),
            .I(N__50158));
    InMux I__10394 (
            .O(N__50201),
            .I(N__50158));
    CascadeMux I__10393 (
            .O(N__50200),
            .I(N__50149));
    InMux I__10392 (
            .O(N__50199),
            .I(N__50144));
    InMux I__10391 (
            .O(N__50198),
            .I(N__50138));
    InMux I__10390 (
            .O(N__50197),
            .I(N__50138));
    LocalMux I__10389 (
            .O(N__50194),
            .I(N__50133));
    LocalMux I__10388 (
            .O(N__50191),
            .I(N__50133));
    InMux I__10387 (
            .O(N__50190),
            .I(N__50128));
    LocalMux I__10386 (
            .O(N__50187),
            .I(N__50120));
    CascadeMux I__10385 (
            .O(N__50186),
            .I(N__50117));
    LocalMux I__10384 (
            .O(N__50183),
            .I(N__50114));
    LocalMux I__10383 (
            .O(N__50178),
            .I(N__50108));
    LocalMux I__10382 (
            .O(N__50175),
            .I(N__50095));
    LocalMux I__10381 (
            .O(N__50172),
            .I(N__50095));
    LocalMux I__10380 (
            .O(N__50169),
            .I(N__50095));
    InMux I__10379 (
            .O(N__50168),
            .I(N__50092));
    Span4Mux_v I__10378 (
            .O(N__50165),
            .I(N__50087));
    LocalMux I__10377 (
            .O(N__50158),
            .I(N__50087));
    InMux I__10376 (
            .O(N__50157),
            .I(N__50084));
    InMux I__10375 (
            .O(N__50156),
            .I(N__50077));
    InMux I__10374 (
            .O(N__50155),
            .I(N__50077));
    InMux I__10373 (
            .O(N__50154),
            .I(N__50077));
    InMux I__10372 (
            .O(N__50153),
            .I(N__50074));
    InMux I__10371 (
            .O(N__50152),
            .I(N__50071));
    InMux I__10370 (
            .O(N__50149),
            .I(N__50068));
    InMux I__10369 (
            .O(N__50148),
            .I(N__50063));
    InMux I__10368 (
            .O(N__50147),
            .I(N__50063));
    LocalMux I__10367 (
            .O(N__50144),
            .I(N__50060));
    InMux I__10366 (
            .O(N__50143),
            .I(N__50057));
    LocalMux I__10365 (
            .O(N__50138),
            .I(N__50052));
    Span4Mux_h I__10364 (
            .O(N__50133),
            .I(N__50052));
    InMux I__10363 (
            .O(N__50132),
            .I(N__50047));
    InMux I__10362 (
            .O(N__50131),
            .I(N__50047));
    LocalMux I__10361 (
            .O(N__50128),
            .I(N__50044));
    InMux I__10360 (
            .O(N__50127),
            .I(N__50041));
    InMux I__10359 (
            .O(N__50126),
            .I(N__50032));
    InMux I__10358 (
            .O(N__50125),
            .I(N__50032));
    InMux I__10357 (
            .O(N__50124),
            .I(N__50032));
    InMux I__10356 (
            .O(N__50123),
            .I(N__50032));
    Span4Mux_v I__10355 (
            .O(N__50120),
            .I(N__50029));
    InMux I__10354 (
            .O(N__50117),
            .I(N__50026));
    Span12Mux_h I__10353 (
            .O(N__50114),
            .I(N__50023));
    InMux I__10352 (
            .O(N__50113),
            .I(N__50012));
    InMux I__10351 (
            .O(N__50112),
            .I(N__50012));
    InMux I__10350 (
            .O(N__50111),
            .I(N__50012));
    Span4Mux_h I__10349 (
            .O(N__50108),
            .I(N__50000));
    InMux I__10348 (
            .O(N__50107),
            .I(N__49991));
    InMux I__10347 (
            .O(N__50106),
            .I(N__49991));
    InMux I__10346 (
            .O(N__50105),
            .I(N__49991));
    InMux I__10345 (
            .O(N__50104),
            .I(N__49991));
    InMux I__10344 (
            .O(N__50103),
            .I(N__49986));
    InMux I__10343 (
            .O(N__50102),
            .I(N__49986));
    Span4Mux_h I__10342 (
            .O(N__50095),
            .I(N__49979));
    LocalMux I__10341 (
            .O(N__50092),
            .I(N__49979));
    Span4Mux_h I__10340 (
            .O(N__50087),
            .I(N__49979));
    LocalMux I__10339 (
            .O(N__50084),
            .I(N__49974));
    LocalMux I__10338 (
            .O(N__50077),
            .I(N__49974));
    LocalMux I__10337 (
            .O(N__50074),
            .I(N__49969));
    LocalMux I__10336 (
            .O(N__50071),
            .I(N__49969));
    LocalMux I__10335 (
            .O(N__50068),
            .I(N__49956));
    LocalMux I__10334 (
            .O(N__50063),
            .I(N__49956));
    Span4Mux_h I__10333 (
            .O(N__50060),
            .I(N__49956));
    LocalMux I__10332 (
            .O(N__50057),
            .I(N__49956));
    Span4Mux_v I__10331 (
            .O(N__50052),
            .I(N__49956));
    LocalMux I__10330 (
            .O(N__50047),
            .I(N__49956));
    Span4Mux_v I__10329 (
            .O(N__50044),
            .I(N__49949));
    LocalMux I__10328 (
            .O(N__50041),
            .I(N__49949));
    LocalMux I__10327 (
            .O(N__50032),
            .I(N__49949));
    Span4Mux_v I__10326 (
            .O(N__50029),
            .I(N__49939));
    LocalMux I__10325 (
            .O(N__50026),
            .I(N__49934));
    Span12Mux_v I__10324 (
            .O(N__50023),
            .I(N__49934));
    InMux I__10323 (
            .O(N__50022),
            .I(N__49925));
    InMux I__10322 (
            .O(N__50021),
            .I(N__49925));
    InMux I__10321 (
            .O(N__50020),
            .I(N__49925));
    InMux I__10320 (
            .O(N__50019),
            .I(N__49925));
    LocalMux I__10319 (
            .O(N__50012),
            .I(N__49922));
    InMux I__10318 (
            .O(N__50011),
            .I(N__49911));
    InMux I__10317 (
            .O(N__50010),
            .I(N__49911));
    InMux I__10316 (
            .O(N__50009),
            .I(N__49911));
    InMux I__10315 (
            .O(N__50008),
            .I(N__49911));
    InMux I__10314 (
            .O(N__50007),
            .I(N__49911));
    InMux I__10313 (
            .O(N__50006),
            .I(N__49902));
    InMux I__10312 (
            .O(N__50005),
            .I(N__49902));
    InMux I__10311 (
            .O(N__50004),
            .I(N__49902));
    InMux I__10310 (
            .O(N__50003),
            .I(N__49902));
    Span4Mux_v I__10309 (
            .O(N__50000),
            .I(N__49893));
    LocalMux I__10308 (
            .O(N__49991),
            .I(N__49893));
    LocalMux I__10307 (
            .O(N__49986),
            .I(N__49893));
    Span4Mux_h I__10306 (
            .O(N__49979),
            .I(N__49893));
    Span4Mux_h I__10305 (
            .O(N__49974),
            .I(N__49888));
    Span4Mux_v I__10304 (
            .O(N__49969),
            .I(N__49888));
    Span4Mux_v I__10303 (
            .O(N__49956),
            .I(N__49883));
    Span4Mux_h I__10302 (
            .O(N__49949),
            .I(N__49883));
    InMux I__10301 (
            .O(N__49948),
            .I(N__49880));
    InMux I__10300 (
            .O(N__49947),
            .I(N__49867));
    InMux I__10299 (
            .O(N__49946),
            .I(N__49867));
    InMux I__10298 (
            .O(N__49945),
            .I(N__49867));
    InMux I__10297 (
            .O(N__49944),
            .I(N__49867));
    InMux I__10296 (
            .O(N__49943),
            .I(N__49867));
    InMux I__10295 (
            .O(N__49942),
            .I(N__49867));
    Odrv4 I__10294 (
            .O(N__49939),
            .I(busState_1));
    Odrv12 I__10293 (
            .O(N__49934),
            .I(busState_1));
    LocalMux I__10292 (
            .O(N__49925),
            .I(busState_1));
    Odrv12 I__10291 (
            .O(N__49922),
            .I(busState_1));
    LocalMux I__10290 (
            .O(N__49911),
            .I(busState_1));
    LocalMux I__10289 (
            .O(N__49902),
            .I(busState_1));
    Odrv4 I__10288 (
            .O(N__49893),
            .I(busState_1));
    Odrv4 I__10287 (
            .O(N__49888),
            .I(busState_1));
    Odrv4 I__10286 (
            .O(N__49883),
            .I(busState_1));
    LocalMux I__10285 (
            .O(N__49880),
            .I(busState_1));
    LocalMux I__10284 (
            .O(N__49867),
            .I(busState_1));
    CascadeMux I__10283 (
            .O(N__49844),
            .I(N_208_cascade_));
    CascadeMux I__10282 (
            .O(N__49841),
            .I(\ALU.status_19_14_cascade_ ));
    InMux I__10281 (
            .O(N__49838),
            .I(N__49835));
    LocalMux I__10280 (
            .O(N__49835),
            .I(N_208));
    InMux I__10279 (
            .O(N__49832),
            .I(N__49826));
    InMux I__10278 (
            .O(N__49831),
            .I(N__49819));
    InMux I__10277 (
            .O(N__49830),
            .I(N__49819));
    InMux I__10276 (
            .O(N__49829),
            .I(N__49812));
    LocalMux I__10275 (
            .O(N__49826),
            .I(N__49807));
    InMux I__10274 (
            .O(N__49825),
            .I(N__49803));
    CascadeMux I__10273 (
            .O(N__49824),
            .I(N__49799));
    LocalMux I__10272 (
            .O(N__49819),
            .I(N__49794));
    InMux I__10271 (
            .O(N__49818),
            .I(N__49790));
    InMux I__10270 (
            .O(N__49817),
            .I(N__49787));
    InMux I__10269 (
            .O(N__49816),
            .I(N__49780));
    InMux I__10268 (
            .O(N__49815),
            .I(N__49780));
    LocalMux I__10267 (
            .O(N__49812),
            .I(N__49777));
    InMux I__10266 (
            .O(N__49811),
            .I(N__49774));
    InMux I__10265 (
            .O(N__49810),
            .I(N__49771));
    Span4Mux_v I__10264 (
            .O(N__49807),
            .I(N__49768));
    InMux I__10263 (
            .O(N__49806),
            .I(N__49765));
    LocalMux I__10262 (
            .O(N__49803),
            .I(N__49762));
    InMux I__10261 (
            .O(N__49802),
            .I(N__49759));
    InMux I__10260 (
            .O(N__49799),
            .I(N__49755));
    InMux I__10259 (
            .O(N__49798),
            .I(N__49752));
    InMux I__10258 (
            .O(N__49797),
            .I(N__49749));
    Span4Mux_h I__10257 (
            .O(N__49794),
            .I(N__49746));
    InMux I__10256 (
            .O(N__49793),
            .I(N__49743));
    LocalMux I__10255 (
            .O(N__49790),
            .I(N__49739));
    LocalMux I__10254 (
            .O(N__49787),
            .I(N__49736));
    InMux I__10253 (
            .O(N__49786),
            .I(N__49733));
    InMux I__10252 (
            .O(N__49785),
            .I(N__49730));
    LocalMux I__10251 (
            .O(N__49780),
            .I(N__49727));
    Span4Mux_v I__10250 (
            .O(N__49777),
            .I(N__49724));
    LocalMux I__10249 (
            .O(N__49774),
            .I(N__49719));
    LocalMux I__10248 (
            .O(N__49771),
            .I(N__49719));
    Span4Mux_h I__10247 (
            .O(N__49768),
            .I(N__49712));
    LocalMux I__10246 (
            .O(N__49765),
            .I(N__49712));
    Span4Mux_v I__10245 (
            .O(N__49762),
            .I(N__49712));
    LocalMux I__10244 (
            .O(N__49759),
            .I(N__49706));
    InMux I__10243 (
            .O(N__49758),
            .I(N__49703));
    LocalMux I__10242 (
            .O(N__49755),
            .I(N__49700));
    LocalMux I__10241 (
            .O(N__49752),
            .I(N__49697));
    LocalMux I__10240 (
            .O(N__49749),
            .I(N__49690));
    Span4Mux_h I__10239 (
            .O(N__49746),
            .I(N__49690));
    LocalMux I__10238 (
            .O(N__49743),
            .I(N__49690));
    InMux I__10237 (
            .O(N__49742),
            .I(N__49687));
    Span12Mux_v I__10236 (
            .O(N__49739),
            .I(N__49684));
    Span12Mux_h I__10235 (
            .O(N__49736),
            .I(N__49681));
    LocalMux I__10234 (
            .O(N__49733),
            .I(N__49678));
    LocalMux I__10233 (
            .O(N__49730),
            .I(N__49675));
    Span4Mux_v I__10232 (
            .O(N__49727),
            .I(N__49666));
    Span4Mux_v I__10231 (
            .O(N__49724),
            .I(N__49666));
    Span4Mux_v I__10230 (
            .O(N__49719),
            .I(N__49666));
    Span4Mux_h I__10229 (
            .O(N__49712),
            .I(N__49666));
    InMux I__10228 (
            .O(N__49711),
            .I(N__49659));
    InMux I__10227 (
            .O(N__49710),
            .I(N__49659));
    InMux I__10226 (
            .O(N__49709),
            .I(N__49659));
    Span4Mux_h I__10225 (
            .O(N__49706),
            .I(N__49652));
    LocalMux I__10224 (
            .O(N__49703),
            .I(N__49652));
    Span4Mux_h I__10223 (
            .O(N__49700),
            .I(N__49652));
    Span4Mux_h I__10222 (
            .O(N__49697),
            .I(N__49647));
    Span4Mux_h I__10221 (
            .O(N__49690),
            .I(N__49647));
    LocalMux I__10220 (
            .O(N__49687),
            .I(busState_0));
    Odrv12 I__10219 (
            .O(N__49684),
            .I(busState_0));
    Odrv12 I__10218 (
            .O(N__49681),
            .I(busState_0));
    Odrv4 I__10217 (
            .O(N__49678),
            .I(busState_0));
    Odrv4 I__10216 (
            .O(N__49675),
            .I(busState_0));
    Odrv4 I__10215 (
            .O(N__49666),
            .I(busState_0));
    LocalMux I__10214 (
            .O(N__49659),
            .I(busState_0));
    Odrv4 I__10213 (
            .O(N__49652),
            .I(busState_0));
    Odrv4 I__10212 (
            .O(N__49647),
            .I(busState_0));
    CascadeMux I__10211 (
            .O(N__49628),
            .I(N__49625));
    InMux I__10210 (
            .O(N__49625),
            .I(N__49622));
    LocalMux I__10209 (
            .O(N__49622),
            .I(N__49619));
    Span4Mux_v I__10208 (
            .O(N__49619),
            .I(N__49616));
    Span4Mux_v I__10207 (
            .O(N__49616),
            .I(N__49613));
    Span4Mux_h I__10206 (
            .O(N__49613),
            .I(N__49610));
    Odrv4 I__10205 (
            .O(N__49610),
            .I(\CONTROL.bus_7_ns_1_15 ));
    InMux I__10204 (
            .O(N__49607),
            .I(N__49601));
    CascadeMux I__10203 (
            .O(N__49606),
            .I(N__49597));
    InMux I__10202 (
            .O(N__49605),
            .I(N__49589));
    InMux I__10201 (
            .O(N__49604),
            .I(N__49584));
    LocalMux I__10200 (
            .O(N__49601),
            .I(N__49569));
    InMux I__10199 (
            .O(N__49600),
            .I(N__49564));
    InMux I__10198 (
            .O(N__49597),
            .I(N__49564));
    InMux I__10197 (
            .O(N__49596),
            .I(N__49554));
    InMux I__10196 (
            .O(N__49595),
            .I(N__49554));
    InMux I__10195 (
            .O(N__49594),
            .I(N__49554));
    InMux I__10194 (
            .O(N__49593),
            .I(N__49547));
    InMux I__10193 (
            .O(N__49592),
            .I(N__49547));
    LocalMux I__10192 (
            .O(N__49589),
            .I(N__49541));
    InMux I__10191 (
            .O(N__49588),
            .I(N__49538));
    InMux I__10190 (
            .O(N__49587),
            .I(N__49535));
    LocalMux I__10189 (
            .O(N__49584),
            .I(N__49529));
    InMux I__10188 (
            .O(N__49583),
            .I(N__49525));
    CascadeMux I__10187 (
            .O(N__49582),
            .I(N__49520));
    InMux I__10186 (
            .O(N__49581),
            .I(N__49516));
    InMux I__10185 (
            .O(N__49580),
            .I(N__49513));
    CascadeMux I__10184 (
            .O(N__49579),
            .I(N__49509));
    CascadeMux I__10183 (
            .O(N__49578),
            .I(N__49506));
    InMux I__10182 (
            .O(N__49577),
            .I(N__49502));
    InMux I__10181 (
            .O(N__49576),
            .I(N__49496));
    InMux I__10180 (
            .O(N__49575),
            .I(N__49496));
    InMux I__10179 (
            .O(N__49574),
            .I(N__49486));
    InMux I__10178 (
            .O(N__49573),
            .I(N__49486));
    InMux I__10177 (
            .O(N__49572),
            .I(N__49486));
    Span4Mux_v I__10176 (
            .O(N__49569),
            .I(N__49481));
    LocalMux I__10175 (
            .O(N__49564),
            .I(N__49481));
    InMux I__10174 (
            .O(N__49563),
            .I(N__49478));
    InMux I__10173 (
            .O(N__49562),
            .I(N__49475));
    InMux I__10172 (
            .O(N__49561),
            .I(N__49472));
    LocalMux I__10171 (
            .O(N__49554),
            .I(N__49469));
    InMux I__10170 (
            .O(N__49553),
            .I(N__49464));
    InMux I__10169 (
            .O(N__49552),
            .I(N__49464));
    LocalMux I__10168 (
            .O(N__49547),
            .I(N__49461));
    InMux I__10167 (
            .O(N__49546),
            .I(N__49456));
    InMux I__10166 (
            .O(N__49545),
            .I(N__49456));
    InMux I__10165 (
            .O(N__49544),
            .I(N__49453));
    Span4Mux_v I__10164 (
            .O(N__49541),
            .I(N__49450));
    LocalMux I__10163 (
            .O(N__49538),
            .I(N__49445));
    LocalMux I__10162 (
            .O(N__49535),
            .I(N__49445));
    InMux I__10161 (
            .O(N__49534),
            .I(N__49438));
    InMux I__10160 (
            .O(N__49533),
            .I(N__49438));
    InMux I__10159 (
            .O(N__49532),
            .I(N__49438));
    Span4Mux_h I__10158 (
            .O(N__49529),
            .I(N__49435));
    CascadeMux I__10157 (
            .O(N__49528),
            .I(N__49432));
    LocalMux I__10156 (
            .O(N__49525),
            .I(N__49428));
    InMux I__10155 (
            .O(N__49524),
            .I(N__49423));
    InMux I__10154 (
            .O(N__49523),
            .I(N__49423));
    InMux I__10153 (
            .O(N__49520),
            .I(N__49418));
    InMux I__10152 (
            .O(N__49519),
            .I(N__49418));
    LocalMux I__10151 (
            .O(N__49516),
            .I(N__49413));
    LocalMux I__10150 (
            .O(N__49513),
            .I(N__49413));
    InMux I__10149 (
            .O(N__49512),
            .I(N__49408));
    InMux I__10148 (
            .O(N__49509),
            .I(N__49408));
    InMux I__10147 (
            .O(N__49506),
            .I(N__49405));
    CascadeMux I__10146 (
            .O(N__49505),
            .I(N__49402));
    LocalMux I__10145 (
            .O(N__49502),
            .I(N__49399));
    InMux I__10144 (
            .O(N__49501),
            .I(N__49396));
    LocalMux I__10143 (
            .O(N__49496),
            .I(N__49393));
    InMux I__10142 (
            .O(N__49495),
            .I(N__49384));
    InMux I__10141 (
            .O(N__49494),
            .I(N__49384));
    InMux I__10140 (
            .O(N__49493),
            .I(N__49384));
    LocalMux I__10139 (
            .O(N__49486),
            .I(N__49375));
    Span4Mux_h I__10138 (
            .O(N__49481),
            .I(N__49375));
    LocalMux I__10137 (
            .O(N__49478),
            .I(N__49375));
    LocalMux I__10136 (
            .O(N__49475),
            .I(N__49375));
    LocalMux I__10135 (
            .O(N__49472),
            .I(N__49370));
    Span4Mux_v I__10134 (
            .O(N__49469),
            .I(N__49370));
    LocalMux I__10133 (
            .O(N__49464),
            .I(N__49367));
    Span4Mux_v I__10132 (
            .O(N__49461),
            .I(N__49364));
    LocalMux I__10131 (
            .O(N__49456),
            .I(N__49361));
    LocalMux I__10130 (
            .O(N__49453),
            .I(N__49354));
    Span4Mux_v I__10129 (
            .O(N__49450),
            .I(N__49354));
    Span4Mux_h I__10128 (
            .O(N__49445),
            .I(N__49354));
    LocalMux I__10127 (
            .O(N__49438),
            .I(N__49351));
    Span4Mux_v I__10126 (
            .O(N__49435),
            .I(N__49348));
    InMux I__10125 (
            .O(N__49432),
            .I(N__49343));
    InMux I__10124 (
            .O(N__49431),
            .I(N__49343));
    Span4Mux_v I__10123 (
            .O(N__49428),
            .I(N__49334));
    LocalMux I__10122 (
            .O(N__49423),
            .I(N__49334));
    LocalMux I__10121 (
            .O(N__49418),
            .I(N__49331));
    Span4Mux_h I__10120 (
            .O(N__49413),
            .I(N__49324));
    LocalMux I__10119 (
            .O(N__49408),
            .I(N__49324));
    LocalMux I__10118 (
            .O(N__49405),
            .I(N__49324));
    InMux I__10117 (
            .O(N__49402),
            .I(N__49317));
    Span4Mux_v I__10116 (
            .O(N__49399),
            .I(N__49312));
    LocalMux I__10115 (
            .O(N__49396),
            .I(N__49312));
    Span4Mux_v I__10114 (
            .O(N__49393),
            .I(N__49309));
    InMux I__10113 (
            .O(N__49392),
            .I(N__49304));
    InMux I__10112 (
            .O(N__49391),
            .I(N__49304));
    LocalMux I__10111 (
            .O(N__49384),
            .I(N__49295));
    Span4Mux_v I__10110 (
            .O(N__49375),
            .I(N__49295));
    Span4Mux_h I__10109 (
            .O(N__49370),
            .I(N__49295));
    Span4Mux_h I__10108 (
            .O(N__49367),
            .I(N__49295));
    Span4Mux_h I__10107 (
            .O(N__49364),
            .I(N__49286));
    Span4Mux_v I__10106 (
            .O(N__49361),
            .I(N__49286));
    Span4Mux_v I__10105 (
            .O(N__49354),
            .I(N__49286));
    Span4Mux_v I__10104 (
            .O(N__49351),
            .I(N__49286));
    Span4Mux_v I__10103 (
            .O(N__49348),
            .I(N__49281));
    LocalMux I__10102 (
            .O(N__49343),
            .I(N__49281));
    InMux I__10101 (
            .O(N__49342),
            .I(N__49272));
    InMux I__10100 (
            .O(N__49341),
            .I(N__49272));
    InMux I__10099 (
            .O(N__49340),
            .I(N__49272));
    InMux I__10098 (
            .O(N__49339),
            .I(N__49272));
    Span4Mux_v I__10097 (
            .O(N__49334),
            .I(N__49269));
    Span4Mux_v I__10096 (
            .O(N__49331),
            .I(N__49264));
    Span4Mux_h I__10095 (
            .O(N__49324),
            .I(N__49264));
    InMux I__10094 (
            .O(N__49323),
            .I(N__49255));
    InMux I__10093 (
            .O(N__49322),
            .I(N__49255));
    InMux I__10092 (
            .O(N__49321),
            .I(N__49255));
    InMux I__10091 (
            .O(N__49320),
            .I(N__49255));
    LocalMux I__10090 (
            .O(N__49317),
            .I(busState_2));
    Odrv4 I__10089 (
            .O(N__49312),
            .I(busState_2));
    Odrv4 I__10088 (
            .O(N__49309),
            .I(busState_2));
    LocalMux I__10087 (
            .O(N__49304),
            .I(busState_2));
    Odrv4 I__10086 (
            .O(N__49295),
            .I(busState_2));
    Odrv4 I__10085 (
            .O(N__49286),
            .I(busState_2));
    Odrv4 I__10084 (
            .O(N__49281),
            .I(busState_2));
    LocalMux I__10083 (
            .O(N__49272),
            .I(busState_2));
    Odrv4 I__10082 (
            .O(N__49269),
            .I(busState_2));
    Odrv4 I__10081 (
            .O(N__49264),
            .I(busState_2));
    LocalMux I__10080 (
            .O(N__49255),
            .I(busState_2));
    IoInMux I__10079 (
            .O(N__49232),
            .I(N__49229));
    LocalMux I__10078 (
            .O(N__49229),
            .I(N__49226));
    IoSpan4Mux I__10077 (
            .O(N__49226),
            .I(N__49223));
    Span4Mux_s3_h I__10076 (
            .O(N__49223),
            .I(N__49220));
    Span4Mux_h I__10075 (
            .O(N__49220),
            .I(N__49216));
    IoInMux I__10074 (
            .O(N__49219),
            .I(N__49213));
    Span4Mux_h I__10073 (
            .O(N__49216),
            .I(N__49210));
    LocalMux I__10072 (
            .O(N__49213),
            .I(N__49207));
    Sp12to4 I__10071 (
            .O(N__49210),
            .I(N__49204));
    Span4Mux_s2_h I__10070 (
            .O(N__49207),
            .I(N__49201));
    Span12Mux_h I__10069 (
            .O(N__49204),
            .I(N__49198));
    Span4Mux_v I__10068 (
            .O(N__49201),
            .I(N__49195));
    Span12Mux_v I__10067 (
            .O(N__49198),
            .I(N__49189));
    Sp12to4 I__10066 (
            .O(N__49195),
            .I(N__49189));
    InMux I__10065 (
            .O(N__49194),
            .I(N__49186));
    Odrv12 I__10064 (
            .O(N__49189),
            .I(bus_15));
    LocalMux I__10063 (
            .O(N__49186),
            .I(bus_15));
    CascadeMux I__10062 (
            .O(N__49181),
            .I(N__49178));
    InMux I__10061 (
            .O(N__49178),
            .I(N__49174));
    CascadeMux I__10060 (
            .O(N__49177),
            .I(N__49171));
    LocalMux I__10059 (
            .O(N__49174),
            .I(N__49168));
    InMux I__10058 (
            .O(N__49171),
            .I(N__49165));
    Span4Mux_v I__10057 (
            .O(N__49168),
            .I(N__49159));
    LocalMux I__10056 (
            .O(N__49165),
            .I(N__49159));
    InMux I__10055 (
            .O(N__49164),
            .I(N__49156));
    Span4Mux_h I__10054 (
            .O(N__49159),
            .I(N__49153));
    LocalMux I__10053 (
            .O(N__49156),
            .I(N__49150));
    Span4Mux_h I__10052 (
            .O(N__49153),
            .I(N__49147));
    Span4Mux_h I__10051 (
            .O(N__49150),
            .I(N__49144));
    Span4Mux_v I__10050 (
            .O(N__49147),
            .I(N__49139));
    Span4Mux_h I__10049 (
            .O(N__49144),
            .I(N__49139));
    Odrv4 I__10048 (
            .O(N__49139),
            .I(f_1));
    CascadeMux I__10047 (
            .O(N__49136),
            .I(N__49133));
    InMux I__10046 (
            .O(N__49133),
            .I(N__49128));
    CascadeMux I__10045 (
            .O(N__49132),
            .I(N__49125));
    InMux I__10044 (
            .O(N__49131),
            .I(N__49122));
    LocalMux I__10043 (
            .O(N__49128),
            .I(N__49119));
    InMux I__10042 (
            .O(N__49125),
            .I(N__49116));
    LocalMux I__10041 (
            .O(N__49122),
            .I(N__49113));
    Span4Mux_v I__10040 (
            .O(N__49119),
            .I(N__49108));
    LocalMux I__10039 (
            .O(N__49116),
            .I(N__49108));
    Span4Mux_v I__10038 (
            .O(N__49113),
            .I(N__49105));
    Span4Mux_v I__10037 (
            .O(N__49108),
            .I(N__49102));
    Span4Mux_v I__10036 (
            .O(N__49105),
            .I(N__49097));
    Span4Mux_h I__10035 (
            .O(N__49102),
            .I(N__49097));
    Span4Mux_h I__10034 (
            .O(N__49097),
            .I(N__49094));
    Odrv4 I__10033 (
            .O(N__49094),
            .I(f_0));
    CascadeMux I__10032 (
            .O(N__49091),
            .I(N__49088));
    InMux I__10031 (
            .O(N__49088),
            .I(N__49085));
    LocalMux I__10030 (
            .O(N__49085),
            .I(N__49082));
    Span4Mux_v I__10029 (
            .O(N__49082),
            .I(N__49077));
    CascadeMux I__10028 (
            .O(N__49081),
            .I(N__49074));
    CascadeMux I__10027 (
            .O(N__49080),
            .I(N__49071));
    Span4Mux_h I__10026 (
            .O(N__49077),
            .I(N__49068));
    InMux I__10025 (
            .O(N__49074),
            .I(N__49063));
    InMux I__10024 (
            .O(N__49071),
            .I(N__49063));
    Span4Mux_h I__10023 (
            .O(N__49068),
            .I(N__49058));
    LocalMux I__10022 (
            .O(N__49063),
            .I(N__49058));
    Span4Mux_v I__10021 (
            .O(N__49058),
            .I(N__49055));
    Odrv4 I__10020 (
            .O(N__49055),
            .I(f_7));
    InMux I__10019 (
            .O(N__49052),
            .I(N__49049));
    LocalMux I__10018 (
            .O(N__49049),
            .I(N__49046));
    Span4Mux_h I__10017 (
            .O(N__49046),
            .I(N__49041));
    InMux I__10016 (
            .O(N__49045),
            .I(N__49038));
    CascadeMux I__10015 (
            .O(N__49044),
            .I(N__49035));
    Span4Mux_v I__10014 (
            .O(N__49041),
            .I(N__49030));
    LocalMux I__10013 (
            .O(N__49038),
            .I(N__49030));
    InMux I__10012 (
            .O(N__49035),
            .I(N__49027));
    Span4Mux_v I__10011 (
            .O(N__49030),
            .I(N__49024));
    LocalMux I__10010 (
            .O(N__49027),
            .I(N__49021));
    Span4Mux_h I__10009 (
            .O(N__49024),
            .I(N__49018));
    Span4Mux_v I__10008 (
            .O(N__49021),
            .I(N__49015));
    Sp12to4 I__10007 (
            .O(N__49018),
            .I(N__49012));
    Span4Mux_h I__10006 (
            .O(N__49015),
            .I(N__49009));
    Span12Mux_h I__10005 (
            .O(N__49012),
            .I(N__49006));
    Span4Mux_h I__10004 (
            .O(N__49009),
            .I(N__49003));
    Odrv12 I__10003 (
            .O(N__49006),
            .I(f_8));
    Odrv4 I__10002 (
            .O(N__49003),
            .I(f_8));
    InMux I__10001 (
            .O(N__48998),
            .I(N__48995));
    LocalMux I__10000 (
            .O(N__48995),
            .I(N__48992));
    Span4Mux_v I__9999 (
            .O(N__48992),
            .I(N__48988));
    CascadeMux I__9998 (
            .O(N__48991),
            .I(N__48985));
    Span4Mux_h I__9997 (
            .O(N__48988),
            .I(N__48982));
    InMux I__9996 (
            .O(N__48985),
            .I(N__48978));
    Span4Mux_h I__9995 (
            .O(N__48982),
            .I(N__48975));
    InMux I__9994 (
            .O(N__48981),
            .I(N__48972));
    LocalMux I__9993 (
            .O(N__48978),
            .I(N__48969));
    Span4Mux_v I__9992 (
            .O(N__48975),
            .I(N__48966));
    LocalMux I__9991 (
            .O(N__48972),
            .I(N__48963));
    Span12Mux_h I__9990 (
            .O(N__48969),
            .I(N__48960));
    Span4Mux_v I__9989 (
            .O(N__48966),
            .I(N__48955));
    Span4Mux_h I__9988 (
            .O(N__48963),
            .I(N__48955));
    Odrv12 I__9987 (
            .O(N__48960),
            .I(f_9));
    Odrv4 I__9986 (
            .O(N__48955),
            .I(f_9));
    InMux I__9985 (
            .O(N__48950),
            .I(N__48947));
    LocalMux I__9984 (
            .O(N__48947),
            .I(N__48944));
    Span4Mux_v I__9983 (
            .O(N__48944),
            .I(N__48939));
    InMux I__9982 (
            .O(N__48943),
            .I(N__48936));
    InMux I__9981 (
            .O(N__48942),
            .I(N__48933));
    Span4Mux_h I__9980 (
            .O(N__48939),
            .I(N__48928));
    LocalMux I__9979 (
            .O(N__48936),
            .I(N__48928));
    LocalMux I__9978 (
            .O(N__48933),
            .I(N__48925));
    Span4Mux_v I__9977 (
            .O(N__48928),
            .I(N__48920));
    Span4Mux_h I__9976 (
            .O(N__48925),
            .I(N__48920));
    Span4Mux_h I__9975 (
            .O(N__48920),
            .I(N__48917));
    Odrv4 I__9974 (
            .O(N__48917),
            .I(g_1));
    CascadeMux I__9973 (
            .O(N__48914),
            .I(N__48911));
    InMux I__9972 (
            .O(N__48911),
            .I(N__48908));
    LocalMux I__9971 (
            .O(N__48908),
            .I(N__48905));
    Span4Mux_v I__9970 (
            .O(N__48905),
            .I(N__48902));
    Span4Mux_h I__9969 (
            .O(N__48902),
            .I(N__48897));
    InMux I__9968 (
            .O(N__48901),
            .I(N__48894));
    InMux I__9967 (
            .O(N__48900),
            .I(N__48891));
    Span4Mux_h I__9966 (
            .O(N__48897),
            .I(N__48886));
    LocalMux I__9965 (
            .O(N__48894),
            .I(N__48886));
    LocalMux I__9964 (
            .O(N__48891),
            .I(N__48883));
    Span4Mux_v I__9963 (
            .O(N__48886),
            .I(N__48878));
    Span4Mux_h I__9962 (
            .O(N__48883),
            .I(N__48878));
    Span4Mux_h I__9961 (
            .O(N__48878),
            .I(N__48875));
    Odrv4 I__9960 (
            .O(N__48875),
            .I(g_0));
    InMux I__9959 (
            .O(N__48872),
            .I(N__48868));
    InMux I__9958 (
            .O(N__48871),
            .I(N__48864));
    LocalMux I__9957 (
            .O(N__48868),
            .I(N__48861));
    CascadeMux I__9956 (
            .O(N__48867),
            .I(N__48858));
    LocalMux I__9955 (
            .O(N__48864),
            .I(N__48855));
    Span12Mux_v I__9954 (
            .O(N__48861),
            .I(N__48852));
    InMux I__9953 (
            .O(N__48858),
            .I(N__48849));
    Span4Mux_v I__9952 (
            .O(N__48855),
            .I(N__48846));
    Span12Mux_h I__9951 (
            .O(N__48852),
            .I(N__48843));
    LocalMux I__9950 (
            .O(N__48849),
            .I(N__48838));
    Sp12to4 I__9949 (
            .O(N__48846),
            .I(N__48838));
    Odrv12 I__9948 (
            .O(N__48843),
            .I(g_7));
    Odrv12 I__9947 (
            .O(N__48838),
            .I(g_7));
    InMux I__9946 (
            .O(N__48833),
            .I(N__48829));
    InMux I__9945 (
            .O(N__48832),
            .I(N__48826));
    LocalMux I__9944 (
            .O(N__48829),
            .I(N__48823));
    LocalMux I__9943 (
            .O(N__48826),
            .I(N__48820));
    Span4Mux_v I__9942 (
            .O(N__48823),
            .I(N__48817));
    Span12Mux_h I__9941 (
            .O(N__48820),
            .I(N__48814));
    Sp12to4 I__9940 (
            .O(N__48817),
            .I(N__48811));
    Odrv12 I__9939 (
            .O(N__48814),
            .I(\ALU.bZ0Z_9 ));
    Odrv12 I__9938 (
            .O(N__48811),
            .I(\ALU.bZ0Z_9 ));
    CascadeMux I__9937 (
            .O(N__48806),
            .I(N__48803));
    InMux I__9936 (
            .O(N__48803),
            .I(N__48800));
    LocalMux I__9935 (
            .O(N__48800),
            .I(N__48797));
    Span4Mux_v I__9934 (
            .O(N__48797),
            .I(N__48794));
    Span4Mux_h I__9933 (
            .O(N__48794),
            .I(N__48791));
    Span4Mux_h I__9932 (
            .O(N__48791),
            .I(N__48787));
    InMux I__9931 (
            .O(N__48790),
            .I(N__48784));
    Odrv4 I__9930 (
            .O(N__48787),
            .I(\ALU.mult_9_8 ));
    LocalMux I__9929 (
            .O(N__48784),
            .I(\ALU.mult_9_8 ));
    InMux I__9928 (
            .O(N__48779),
            .I(N__48776));
    LocalMux I__9927 (
            .O(N__48776),
            .I(N__48773));
    Span4Mux_v I__9926 (
            .O(N__48773),
            .I(N__48769));
    CascadeMux I__9925 (
            .O(N__48772),
            .I(N__48766));
    Span4Mux_h I__9924 (
            .O(N__48769),
            .I(N__48763));
    InMux I__9923 (
            .O(N__48766),
            .I(N__48760));
    Odrv4 I__9922 (
            .O(N__48763),
            .I(\ALU.mult_25_8 ));
    LocalMux I__9921 (
            .O(N__48760),
            .I(\ALU.mult_25_8 ));
    CascadeMux I__9920 (
            .O(N__48755),
            .I(\ALU.mult_495_c_RNIKOB51JZ0_cascade_ ));
    InMux I__9919 (
            .O(N__48752),
            .I(N__48749));
    LocalMux I__9918 (
            .O(N__48749),
            .I(N__48746));
    Span4Mux_v I__9917 (
            .O(N__48746),
            .I(N__48742));
    InMux I__9916 (
            .O(N__48745),
            .I(N__48739));
    Span4Mux_h I__9915 (
            .O(N__48742),
            .I(N__48736));
    LocalMux I__9914 (
            .O(N__48739),
            .I(N__48733));
    Span4Mux_h I__9913 (
            .O(N__48736),
            .I(N__48730));
    Span12Mux_h I__9912 (
            .O(N__48733),
            .I(N__48727));
    Span4Mux_v I__9911 (
            .O(N__48730),
            .I(N__48724));
    Odrv12 I__9910 (
            .O(N__48727),
            .I(\ALU.aZ0Z_8 ));
    Odrv4 I__9909 (
            .O(N__48724),
            .I(\ALU.aZ0Z_8 ));
    CascadeMux I__9908 (
            .O(N__48719),
            .I(N__48716));
    InMux I__9907 (
            .O(N__48716),
            .I(N__48713));
    LocalMux I__9906 (
            .O(N__48713),
            .I(\ALU.lshift_15_ns_1_8 ));
    InMux I__9905 (
            .O(N__48710),
            .I(N__48706));
    InMux I__9904 (
            .O(N__48709),
            .I(N__48703));
    LocalMux I__9903 (
            .O(N__48706),
            .I(N__48700));
    LocalMux I__9902 (
            .O(N__48703),
            .I(N__48697));
    Span4Mux_h I__9901 (
            .O(N__48700),
            .I(N__48694));
    Span4Mux_v I__9900 (
            .O(N__48697),
            .I(N__48691));
    Span4Mux_h I__9899 (
            .O(N__48694),
            .I(N__48688));
    Span4Mux_h I__9898 (
            .O(N__48691),
            .I(N__48685));
    Span4Mux_v I__9897 (
            .O(N__48688),
            .I(N__48680));
    Span4Mux_h I__9896 (
            .O(N__48685),
            .I(N__48680));
    Odrv4 I__9895 (
            .O(N__48680),
            .I(\ALU.N_610 ));
    InMux I__9894 (
            .O(N__48677),
            .I(N__48674));
    LocalMux I__9893 (
            .O(N__48674),
            .I(N__48669));
    InMux I__9892 (
            .O(N__48673),
            .I(N__48666));
    InMux I__9891 (
            .O(N__48672),
            .I(N__48663));
    Span4Mux_v I__9890 (
            .O(N__48669),
            .I(N__48660));
    LocalMux I__9889 (
            .O(N__48666),
            .I(N__48657));
    LocalMux I__9888 (
            .O(N__48663),
            .I(N__48654));
    Span4Mux_h I__9887 (
            .O(N__48660),
            .I(N__48651));
    Span4Mux_h I__9886 (
            .O(N__48657),
            .I(N__48648));
    Span4Mux_v I__9885 (
            .O(N__48654),
            .I(N__48645));
    Span4Mux_h I__9884 (
            .O(N__48651),
            .I(N__48640));
    Span4Mux_v I__9883 (
            .O(N__48648),
            .I(N__48640));
    Span4Mux_h I__9882 (
            .O(N__48645),
            .I(N__48637));
    Sp12to4 I__9881 (
            .O(N__48640),
            .I(N__48634));
    Span4Mux_h I__9880 (
            .O(N__48637),
            .I(N__48631));
    Odrv12 I__9879 (
            .O(N__48634),
            .I(\ALU.N_608 ));
    Odrv4 I__9878 (
            .O(N__48631),
            .I(\ALU.N_608 ));
    InMux I__9877 (
            .O(N__48626),
            .I(N__48623));
    LocalMux I__9876 (
            .O(N__48623),
            .I(\ALU.N_640 ));
    CascadeMux I__9875 (
            .O(N__48620),
            .I(\ALU.addsub_cry_7_c_RNIDLTNZ0Z71_cascade_ ));
    InMux I__9874 (
            .O(N__48617),
            .I(N__48614));
    LocalMux I__9873 (
            .O(N__48614),
            .I(\ALU.lshift_8 ));
    InMux I__9872 (
            .O(N__48611),
            .I(N__48607));
    InMux I__9871 (
            .O(N__48610),
            .I(N__48604));
    LocalMux I__9870 (
            .O(N__48607),
            .I(N__48599));
    LocalMux I__9869 (
            .O(N__48604),
            .I(N__48599));
    Odrv4 I__9868 (
            .O(N__48599),
            .I(\ALU.N_636 ));
    CascadeMux I__9867 (
            .O(N__48596),
            .I(N__48592));
    CascadeMux I__9866 (
            .O(N__48595),
            .I(N__48589));
    InMux I__9865 (
            .O(N__48592),
            .I(N__48584));
    InMux I__9864 (
            .O(N__48589),
            .I(N__48584));
    LocalMux I__9863 (
            .O(N__48584),
            .I(N__48580));
    InMux I__9862 (
            .O(N__48583),
            .I(N__48577));
    Span4Mux_v I__9861 (
            .O(N__48580),
            .I(N__48574));
    LocalMux I__9860 (
            .O(N__48577),
            .I(N__48571));
    Span4Mux_v I__9859 (
            .O(N__48574),
            .I(N__48568));
    Span4Mux_v I__9858 (
            .O(N__48571),
            .I(N__48565));
    Span4Mux_h I__9857 (
            .O(N__48568),
            .I(N__48562));
    Span4Mux_v I__9856 (
            .O(N__48565),
            .I(N__48559));
    Odrv4 I__9855 (
            .O(N__48562),
            .I(\ALU.N_794_1 ));
    Odrv4 I__9854 (
            .O(N__48559),
            .I(\ALU.N_794_1 ));
    InMux I__9853 (
            .O(N__48554),
            .I(N__48551));
    LocalMux I__9852 (
            .O(N__48551),
            .I(N__48548));
    Span4Mux_v I__9851 (
            .O(N__48548),
            .I(N__48545));
    Span4Mux_h I__9850 (
            .O(N__48545),
            .I(N__48542));
    Span4Mux_h I__9849 (
            .O(N__48542),
            .I(N__48539));
    Span4Mux_h I__9848 (
            .O(N__48539),
            .I(N__48536));
    Span4Mux_h I__9847 (
            .O(N__48536),
            .I(N__48532));
    InMux I__9846 (
            .O(N__48535),
            .I(N__48529));
    Span4Mux_h I__9845 (
            .O(N__48532),
            .I(N__48526));
    LocalMux I__9844 (
            .O(N__48529),
            .I(N__48523));
    Odrv4 I__9843 (
            .O(N__48526),
            .I(\ALU.N_809 ));
    Odrv12 I__9842 (
            .O(N__48523),
            .I(\ALU.N_809 ));
    InMux I__9841 (
            .O(N__48518),
            .I(N__48515));
    LocalMux I__9840 (
            .O(N__48515),
            .I(N__48512));
    Span4Mux_h I__9839 (
            .O(N__48512),
            .I(N__48509));
    Odrv4 I__9838 (
            .O(N__48509),
            .I(\ALU.mult_12 ));
    InMux I__9837 (
            .O(N__48506),
            .I(N__48503));
    LocalMux I__9836 (
            .O(N__48503),
            .I(\ALU.mult_555_c_RNI5VJUOIZ0 ));
    InMux I__9835 (
            .O(N__48500),
            .I(N__48497));
    LocalMux I__9834 (
            .O(N__48497),
            .I(N__48494));
    Span4Mux_h I__9833 (
            .O(N__48494),
            .I(N__48491));
    Odrv4 I__9832 (
            .O(N__48491),
            .I(\ALU.mult_546_c_RNIG1E6IZ0Z8 ));
    CascadeMux I__9831 (
            .O(N__48488),
            .I(N__48484));
    InMux I__9830 (
            .O(N__48487),
            .I(N__48481));
    InMux I__9829 (
            .O(N__48484),
            .I(N__48478));
    LocalMux I__9828 (
            .O(N__48481),
            .I(N__48475));
    LocalMux I__9827 (
            .O(N__48478),
            .I(N__48472));
    Span4Mux_v I__9826 (
            .O(N__48475),
            .I(N__48469));
    Span4Mux_v I__9825 (
            .O(N__48472),
            .I(N__48465));
    Span4Mux_v I__9824 (
            .O(N__48469),
            .I(N__48460));
    InMux I__9823 (
            .O(N__48468),
            .I(N__48457));
    Span4Mux_h I__9822 (
            .O(N__48465),
            .I(N__48454));
    CascadeMux I__9821 (
            .O(N__48464),
            .I(N__48450));
    InMux I__9820 (
            .O(N__48463),
            .I(N__48447));
    Span4Mux_h I__9819 (
            .O(N__48460),
            .I(N__48440));
    LocalMux I__9818 (
            .O(N__48457),
            .I(N__48440));
    Span4Mux_h I__9817 (
            .O(N__48454),
            .I(N__48440));
    InMux I__9816 (
            .O(N__48453),
            .I(N__48435));
    InMux I__9815 (
            .O(N__48450),
            .I(N__48435));
    LocalMux I__9814 (
            .O(N__48447),
            .I(aluStatus_0));
    Odrv4 I__9813 (
            .O(N__48440),
            .I(aluStatus_0));
    LocalMux I__9812 (
            .O(N__48435),
            .I(aluStatus_0));
    CascadeMux I__9811 (
            .O(N__48428),
            .I(\ALU.status_14_12_0_cascade_ ));
    InMux I__9810 (
            .O(N__48425),
            .I(N__48422));
    LocalMux I__9809 (
            .O(N__48422),
            .I(N__48419));
    Span4Mux_h I__9808 (
            .O(N__48419),
            .I(N__48416));
    Span4Mux_v I__9807 (
            .O(N__48416),
            .I(N__48413));
    Odrv4 I__9806 (
            .O(N__48413),
            .I(\ALU.status_RNO_1Z0Z_0 ));
    InMux I__9805 (
            .O(N__48410),
            .I(N__48406));
    InMux I__9804 (
            .O(N__48409),
            .I(N__48403));
    LocalMux I__9803 (
            .O(N__48406),
            .I(N__48400));
    LocalMux I__9802 (
            .O(N__48403),
            .I(N__48397));
    Span4Mux_v I__9801 (
            .O(N__48400),
            .I(N__48392));
    Span4Mux_v I__9800 (
            .O(N__48397),
            .I(N__48392));
    Span4Mux_h I__9799 (
            .O(N__48392),
            .I(N__48389));
    Span4Mux_h I__9798 (
            .O(N__48389),
            .I(N__48386));
    Span4Mux_v I__9797 (
            .O(N__48386),
            .I(N__48383));
    Odrv4 I__9796 (
            .O(N__48383),
            .I(\ALU.bZ0Z_1 ));
    InMux I__9795 (
            .O(N__48380),
            .I(N__48377));
    LocalMux I__9794 (
            .O(N__48377),
            .I(N__48373));
    InMux I__9793 (
            .O(N__48376),
            .I(N__48370));
    Span4Mux_v I__9792 (
            .O(N__48373),
            .I(N__48367));
    LocalMux I__9791 (
            .O(N__48370),
            .I(N__48364));
    Span4Mux_h I__9790 (
            .O(N__48367),
            .I(N__48361));
    Span4Mux_h I__9789 (
            .O(N__48364),
            .I(N__48358));
    Span4Mux_h I__9788 (
            .O(N__48361),
            .I(N__48353));
    Span4Mux_h I__9787 (
            .O(N__48358),
            .I(N__48353));
    Span4Mux_v I__9786 (
            .O(N__48353),
            .I(N__48350));
    Odrv4 I__9785 (
            .O(N__48350),
            .I(\ALU.bZ0Z_0 ));
    InMux I__9784 (
            .O(N__48347),
            .I(N__48343));
    InMux I__9783 (
            .O(N__48346),
            .I(N__48340));
    LocalMux I__9782 (
            .O(N__48343),
            .I(N__48335));
    LocalMux I__9781 (
            .O(N__48340),
            .I(N__48335));
    Span4Mux_h I__9780 (
            .O(N__48335),
            .I(N__48332));
    Span4Mux_v I__9779 (
            .O(N__48332),
            .I(N__48329));
    Odrv4 I__9778 (
            .O(N__48329),
            .I(\ALU.bZ0Z_7 ));
    InMux I__9777 (
            .O(N__48326),
            .I(N__48322));
    InMux I__9776 (
            .O(N__48325),
            .I(N__48319));
    LocalMux I__9775 (
            .O(N__48322),
            .I(N__48316));
    LocalMux I__9774 (
            .O(N__48319),
            .I(N__48313));
    Span4Mux_h I__9773 (
            .O(N__48316),
            .I(N__48310));
    Span4Mux_v I__9772 (
            .O(N__48313),
            .I(N__48307));
    Span4Mux_h I__9771 (
            .O(N__48310),
            .I(N__48304));
    Span4Mux_h I__9770 (
            .O(N__48307),
            .I(N__48301));
    Span4Mux_h I__9769 (
            .O(N__48304),
            .I(N__48298));
    Span4Mux_h I__9768 (
            .O(N__48301),
            .I(N__48295));
    Odrv4 I__9767 (
            .O(N__48298),
            .I(\ALU.bZ0Z_8 ));
    Odrv4 I__9766 (
            .O(N__48295),
            .I(\ALU.bZ0Z_8 ));
    InMux I__9765 (
            .O(N__48290),
            .I(N__48287));
    LocalMux I__9764 (
            .O(N__48287),
            .I(N__48284));
    Span4Mux_v I__9763 (
            .O(N__48284),
            .I(N__48281));
    Span4Mux_h I__9762 (
            .O(N__48281),
            .I(N__48278));
    Span4Mux_h I__9761 (
            .O(N__48278),
            .I(N__48275));
    Odrv4 I__9760 (
            .O(N__48275),
            .I(\ALU.d_RNILTVJG3Z0Z_3 ));
    CascadeMux I__9759 (
            .O(N__48272),
            .I(\ALU.mult_555_c_RNIJF56AMZ0_cascade_ ));
    InMux I__9758 (
            .O(N__48269),
            .I(N__48266));
    LocalMux I__9757 (
            .O(N__48266),
            .I(N__48262));
    InMux I__9756 (
            .O(N__48265),
            .I(N__48259));
    Span4Mux_h I__9755 (
            .O(N__48262),
            .I(N__48256));
    LocalMux I__9754 (
            .O(N__48259),
            .I(N__48253));
    Span4Mux_h I__9753 (
            .O(N__48256),
            .I(N__48250));
    Span4Mux_v I__9752 (
            .O(N__48253),
            .I(N__48247));
    Span4Mux_v I__9751 (
            .O(N__48250),
            .I(N__48242));
    Span4Mux_h I__9750 (
            .O(N__48247),
            .I(N__48242));
    Span4Mux_h I__9749 (
            .O(N__48242),
            .I(N__48239));
    Odrv4 I__9748 (
            .O(N__48239),
            .I(\ALU.aZ0Z_12 ));
    InMux I__9747 (
            .O(N__48236),
            .I(N__48233));
    LocalMux I__9746 (
            .O(N__48233),
            .I(N__48229));
    InMux I__9745 (
            .O(N__48232),
            .I(N__48226));
    Span4Mux_v I__9744 (
            .O(N__48229),
            .I(N__48223));
    LocalMux I__9743 (
            .O(N__48226),
            .I(N__48220));
    Span4Mux_h I__9742 (
            .O(N__48223),
            .I(N__48217));
    Odrv4 I__9741 (
            .O(N__48220),
            .I(\ALU.N_612 ));
    Odrv4 I__9740 (
            .O(N__48217),
            .I(\ALU.N_612 ));
    CascadeMux I__9739 (
            .O(N__48212),
            .I(N__48209));
    InMux I__9738 (
            .O(N__48209),
            .I(N__48206));
    LocalMux I__9737 (
            .O(N__48206),
            .I(N__48203));
    Span4Mux_v I__9736 (
            .O(N__48203),
            .I(N__48200));
    Span4Mux_h I__9735 (
            .O(N__48200),
            .I(N__48197));
    Odrv4 I__9734 (
            .O(N__48197),
            .I(\ALU.N_614 ));
    CascadeMux I__9733 (
            .O(N__48194),
            .I(\ALU.lshift_7_ns_1_12_cascade_ ));
    CascadeMux I__9732 (
            .O(N__48191),
            .I(\ALU.N_704_cascade_ ));
    CascadeMux I__9731 (
            .O(N__48188),
            .I(N__48185));
    InMux I__9730 (
            .O(N__48185),
            .I(N__48182));
    LocalMux I__9729 (
            .O(N__48182),
            .I(\ALU.d_RNIGNBT49Z0Z_8 ));
    CascadeMux I__9728 (
            .O(N__48179),
            .I(\ALU.d_RNIGNBT49Z0Z_8_cascade_ ));
    InMux I__9727 (
            .O(N__48176),
            .I(N__48171));
    InMux I__9726 (
            .O(N__48175),
            .I(N__48166));
    InMux I__9725 (
            .O(N__48174),
            .I(N__48166));
    LocalMux I__9724 (
            .O(N__48171),
            .I(N__48163));
    LocalMux I__9723 (
            .O(N__48166),
            .I(N__48158));
    Span4Mux_h I__9722 (
            .O(N__48163),
            .I(N__48158));
    Span4Mux_v I__9721 (
            .O(N__48158),
            .I(N__48155));
    Span4Mux_h I__9720 (
            .O(N__48155),
            .I(N__48152));
    Span4Mux_v I__9719 (
            .O(N__48152),
            .I(N__48149));
    Odrv4 I__9718 (
            .O(N__48149),
            .I(\ALU.N_18_0 ));
    CascadeMux I__9717 (
            .O(N__48146),
            .I(N__48143));
    InMux I__9716 (
            .O(N__48143),
            .I(N__48138));
    InMux I__9715 (
            .O(N__48142),
            .I(N__48135));
    InMux I__9714 (
            .O(N__48141),
            .I(N__48132));
    LocalMux I__9713 (
            .O(N__48138),
            .I(N__48129));
    LocalMux I__9712 (
            .O(N__48135),
            .I(N__48126));
    LocalMux I__9711 (
            .O(N__48132),
            .I(N__48123));
    Span4Mux_v I__9710 (
            .O(N__48129),
            .I(N__48118));
    Span4Mux_h I__9709 (
            .O(N__48126),
            .I(N__48118));
    Span4Mux_h I__9708 (
            .O(N__48123),
            .I(N__48115));
    Span4Mux_h I__9707 (
            .O(N__48118),
            .I(N__48112));
    Span4Mux_v I__9706 (
            .O(N__48115),
            .I(N__48109));
    Span4Mux_h I__9705 (
            .O(N__48112),
            .I(N__48106));
    Span4Mux_h I__9704 (
            .O(N__48109),
            .I(N__48103));
    Span4Mux_v I__9703 (
            .O(N__48106),
            .I(N__48100));
    Sp12to4 I__9702 (
            .O(N__48103),
            .I(N__48097));
    Odrv4 I__9701 (
            .O(N__48100),
            .I(h_8));
    Odrv12 I__9700 (
            .O(N__48097),
            .I(h_8));
    CascadeMux I__9699 (
            .O(N__48092),
            .I(\ALU.lshift_3_ns_1_13_cascade_ ));
    CascadeMux I__9698 (
            .O(N__48089),
            .I(\ALU.N_645_cascade_ ));
    InMux I__9697 (
            .O(N__48086),
            .I(N__48083));
    LocalMux I__9696 (
            .O(N__48083),
            .I(N__48079));
    InMux I__9695 (
            .O(N__48082),
            .I(N__48076));
    Span4Mux_v I__9694 (
            .O(N__48079),
            .I(N__48073));
    LocalMux I__9693 (
            .O(N__48076),
            .I(N__48068));
    Span4Mux_h I__9692 (
            .O(N__48073),
            .I(N__48068));
    Odrv4 I__9691 (
            .O(N__48068),
            .I(\ALU.N_806_1 ));
    CascadeMux I__9690 (
            .O(N__48065),
            .I(\ALU.a_15_m1_am_1_13_cascade_ ));
    CascadeMux I__9689 (
            .O(N__48062),
            .I(\ALU.N_611_cascade_ ));
    InMux I__9688 (
            .O(N__48059),
            .I(N__48055));
    InMux I__9687 (
            .O(N__48058),
            .I(N__48052));
    LocalMux I__9686 (
            .O(N__48055),
            .I(N__48049));
    LocalMux I__9685 (
            .O(N__48052),
            .I(N__48046));
    Span4Mux_h I__9684 (
            .O(N__48049),
            .I(N__48043));
    Span12Mux_h I__9683 (
            .O(N__48046),
            .I(N__48040));
    Span4Mux_h I__9682 (
            .O(N__48043),
            .I(N__48037));
    Odrv12 I__9681 (
            .O(N__48040),
            .I(\ALU.N_609 ));
    Odrv4 I__9680 (
            .O(N__48037),
            .I(\ALU.N_609 ));
    InMux I__9679 (
            .O(N__48032),
            .I(N__48029));
    LocalMux I__9678 (
            .O(N__48029),
            .I(\ALU.N_641 ));
    CascadeMux I__9677 (
            .O(N__48026),
            .I(\ALU.N_641_cascade_ ));
    InMux I__9676 (
            .O(N__48023),
            .I(N__48020));
    LocalMux I__9675 (
            .O(N__48020),
            .I(N__48017));
    Span4Mux_v I__9674 (
            .O(N__48017),
            .I(N__48012));
    InMux I__9673 (
            .O(N__48016),
            .I(N__48007));
    InMux I__9672 (
            .O(N__48015),
            .I(N__48007));
    Odrv4 I__9671 (
            .O(N__48012),
            .I(\ALU.N_637 ));
    LocalMux I__9670 (
            .O(N__48007),
            .I(\ALU.N_637 ));
    InMux I__9669 (
            .O(N__48002),
            .I(N__47999));
    LocalMux I__9668 (
            .O(N__47999),
            .I(N__47996));
    Span12Mux_v I__9667 (
            .O(N__47996),
            .I(N__47993));
    Odrv12 I__9666 (
            .O(N__47993),
            .I(\ALU.d_RNITG2137Z0Z_0 ));
    CascadeMux I__9665 (
            .O(N__47990),
            .I(N__47987));
    InMux I__9664 (
            .O(N__47987),
            .I(N__47982));
    InMux I__9663 (
            .O(N__47986),
            .I(N__47979));
    InMux I__9662 (
            .O(N__47985),
            .I(N__47975));
    LocalMux I__9661 (
            .O(N__47982),
            .I(N__47972));
    LocalMux I__9660 (
            .O(N__47979),
            .I(N__47969));
    InMux I__9659 (
            .O(N__47978),
            .I(N__47966));
    LocalMux I__9658 (
            .O(N__47975),
            .I(N__47963));
    Span4Mux_h I__9657 (
            .O(N__47972),
            .I(N__47960));
    Span4Mux_v I__9656 (
            .O(N__47969),
            .I(N__47957));
    LocalMux I__9655 (
            .O(N__47966),
            .I(N__47954));
    Span4Mux_h I__9654 (
            .O(N__47963),
            .I(N__47949));
    Span4Mux_h I__9653 (
            .O(N__47960),
            .I(N__47949));
    Odrv4 I__9652 (
            .O(N__47957),
            .I(\ALU.N_765 ));
    Odrv12 I__9651 (
            .O(N__47954),
            .I(\ALU.N_765 ));
    Odrv4 I__9650 (
            .O(N__47949),
            .I(\ALU.N_765 ));
    InMux I__9649 (
            .O(N__47942),
            .I(N__47939));
    LocalMux I__9648 (
            .O(N__47939),
            .I(\ALU.a_15_m1_am_1_9 ));
    InMux I__9647 (
            .O(N__47936),
            .I(N__47933));
    LocalMux I__9646 (
            .O(N__47933),
            .I(N__47930));
    Span4Mux_h I__9645 (
            .O(N__47930),
            .I(N__47927));
    Span4Mux_h I__9644 (
            .O(N__47927),
            .I(N__47924));
    Span4Mux_h I__9643 (
            .O(N__47924),
            .I(N__47921));
    Odrv4 I__9642 (
            .O(N__47921),
            .I(\ALU.a_15_m3_d_d_0_ns_1_3 ));
    CascadeMux I__9641 (
            .O(N__47918),
            .I(\PROM.ROMDATA.m451_bm_cascade_ ));
    InMux I__9640 (
            .O(N__47915),
            .I(N__47912));
    LocalMux I__9639 (
            .O(N__47912),
            .I(N__47909));
    Odrv12 I__9638 (
            .O(N__47909),
            .I(\PROM.ROMDATA.m451_am ));
    CascadeMux I__9637 (
            .O(N__47906),
            .I(N__47903));
    InMux I__9636 (
            .O(N__47903),
            .I(N__47900));
    LocalMux I__9635 (
            .O(N__47900),
            .I(\PROM.ROMDATA.m451_ns ));
    CascadeMux I__9634 (
            .O(N__47897),
            .I(N__47894));
    InMux I__9633 (
            .O(N__47894),
            .I(N__47891));
    LocalMux I__9632 (
            .O(N__47891),
            .I(N__47888));
    Odrv12 I__9631 (
            .O(N__47888),
            .I(\PROM.ROMDATA.m375_bm ));
    CascadeMux I__9630 (
            .O(N__47885),
            .I(N__47882));
    InMux I__9629 (
            .O(N__47882),
            .I(N__47879));
    LocalMux I__9628 (
            .O(N__47879),
            .I(N__47876));
    Odrv4 I__9627 (
            .O(N__47876),
            .I(\PROM.ROMDATA.m376 ));
    InMux I__9626 (
            .O(N__47873),
            .I(N__47870));
    LocalMux I__9625 (
            .O(N__47870),
            .I(\PROM.ROMDATA.N_256_i ));
    InMux I__9624 (
            .O(N__47867),
            .I(N__47864));
    LocalMux I__9623 (
            .O(N__47864),
            .I(N__47861));
    Odrv4 I__9622 (
            .O(N__47861),
            .I(\PROM.ROMDATA.m389_bm ));
    CascadeMux I__9621 (
            .O(N__47858),
            .I(\PROM.ROMDATA.m389_am_cascade_ ));
    InMux I__9620 (
            .O(N__47855),
            .I(N__47852));
    LocalMux I__9619 (
            .O(N__47852),
            .I(N__47849));
    Odrv4 I__9618 (
            .O(N__47849),
            .I(\PROM.ROMDATA.m389_ns ));
    InMux I__9617 (
            .O(N__47846),
            .I(N__47843));
    LocalMux I__9616 (
            .O(N__47843),
            .I(N__47840));
    Span4Mux_v I__9615 (
            .O(N__47840),
            .I(N__47836));
    InMux I__9614 (
            .O(N__47839),
            .I(N__47833));
    Span4Mux_h I__9613 (
            .O(N__47836),
            .I(N__47830));
    LocalMux I__9612 (
            .O(N__47833),
            .I(N__47827));
    Span4Mux_h I__9611 (
            .O(N__47830),
            .I(N__47824));
    Span4Mux_h I__9610 (
            .O(N__47827),
            .I(N__47821));
    Odrv4 I__9609 (
            .O(N__47824),
            .I(\CONTROL.programCounter_1_6 ));
    Odrv4 I__9608 (
            .O(N__47821),
            .I(\CONTROL.programCounter_1_6 ));
    CascadeMux I__9607 (
            .O(N__47816),
            .I(N__47813));
    InMux I__9606 (
            .O(N__47813),
            .I(N__47810));
    LocalMux I__9605 (
            .O(N__47810),
            .I(N__47807));
    Odrv4 I__9604 (
            .O(N__47807),
            .I(\CONTROL.programCounter_1_reto_6 ));
    InMux I__9603 (
            .O(N__47804),
            .I(N__47801));
    LocalMux I__9602 (
            .O(N__47801),
            .I(\PROM.ROMDATA.m51 ));
    InMux I__9601 (
            .O(N__47798),
            .I(N__47795));
    LocalMux I__9600 (
            .O(N__47795),
            .I(N__47792));
    Span4Mux_h I__9599 (
            .O(N__47792),
            .I(N__47789));
    Odrv4 I__9598 (
            .O(N__47789),
            .I(\PROM.ROMDATA.m433_am ));
    CascadeMux I__9597 (
            .O(N__47786),
            .I(\PROM.ROMDATA.m399_am_cascade_ ));
    InMux I__9596 (
            .O(N__47783),
            .I(N__47780));
    LocalMux I__9595 (
            .O(N__47780),
            .I(N__47777));
    Span12Mux_v I__9594 (
            .O(N__47777),
            .I(N__47774));
    Odrv12 I__9593 (
            .O(N__47774),
            .I(\PROM.ROMDATA.m399_bm ));
    InMux I__9592 (
            .O(N__47771),
            .I(N__47768));
    LocalMux I__9591 (
            .O(N__47768),
            .I(N__47765));
    Odrv4 I__9590 (
            .O(N__47765),
            .I(\PROM.ROMDATA.m399_ns ));
    InMux I__9589 (
            .O(N__47762),
            .I(N__47759));
    LocalMux I__9588 (
            .O(N__47759),
            .I(N__47756));
    Span4Mux_h I__9587 (
            .O(N__47756),
            .I(N__47753));
    Span4Mux_h I__9586 (
            .O(N__47753),
            .I(N__47750));
    Span4Mux_h I__9585 (
            .O(N__47750),
            .I(N__47747));
    Odrv4 I__9584 (
            .O(N__47747),
            .I(\PROM.ROMDATA.m461_ns_1 ));
    InMux I__9583 (
            .O(N__47744),
            .I(N__47741));
    LocalMux I__9582 (
            .O(N__47741),
            .I(N__47738));
    Span4Mux_v I__9581 (
            .O(N__47738),
            .I(N__47735));
    Span4Mux_h I__9580 (
            .O(N__47735),
            .I(N__47732));
    Span4Mux_h I__9579 (
            .O(N__47732),
            .I(N__47729));
    Odrv4 I__9578 (
            .O(N__47729),
            .I(\CONTROL.addrstack_4 ));
    InMux I__9577 (
            .O(N__47726),
            .I(N__47723));
    LocalMux I__9576 (
            .O(N__47723),
            .I(N__47720));
    Odrv12 I__9575 (
            .O(N__47720),
            .I(\PROM.ROMDATA.m22 ));
    CascadeMux I__9574 (
            .O(N__47717),
            .I(\PROM.ROMDATA.m215_ns_1_1_1_cascade_ ));
    InMux I__9573 (
            .O(N__47714),
            .I(N__47711));
    LocalMux I__9572 (
            .O(N__47711),
            .I(\PROM.ROMDATA.m215_ns_1_1 ));
    InMux I__9571 (
            .O(N__47708),
            .I(N__47705));
    LocalMux I__9570 (
            .O(N__47705),
            .I(\PROM.ROMDATA.m256 ));
    InMux I__9569 (
            .O(N__47702),
            .I(N__47699));
    LocalMux I__9568 (
            .O(N__47699),
            .I(N__47696));
    Odrv12 I__9567 (
            .O(N__47696),
            .I(\PROM.ROMDATA.m38 ));
    InMux I__9566 (
            .O(N__47693),
            .I(N__47690));
    LocalMux I__9565 (
            .O(N__47690),
            .I(\PROM.ROMDATA.m251 ));
    InMux I__9564 (
            .O(N__47687),
            .I(N__47684));
    LocalMux I__9563 (
            .O(N__47684),
            .I(\PROM.ROMDATA.m253 ));
    CascadeMux I__9562 (
            .O(N__47681),
            .I(N__47677));
    CascadeMux I__9561 (
            .O(N__47680),
            .I(N__47674));
    InMux I__9560 (
            .O(N__47677),
            .I(N__47669));
    InMux I__9559 (
            .O(N__47674),
            .I(N__47669));
    LocalMux I__9558 (
            .O(N__47669),
            .I(N__47666));
    Span4Mux_v I__9557 (
            .O(N__47666),
            .I(N__47663));
    Odrv4 I__9556 (
            .O(N__47663),
            .I(N_419));
    InMux I__9555 (
            .O(N__47660),
            .I(N__47657));
    LocalMux I__9554 (
            .O(N__47657),
            .I(N__47654));
    Span4Mux_v I__9553 (
            .O(N__47654),
            .I(N__47651));
    Span4Mux_h I__9552 (
            .O(N__47651),
            .I(N__47648));
    Span4Mux_h I__9551 (
            .O(N__47648),
            .I(N__47645));
    Span4Mux_h I__9550 (
            .O(N__47645),
            .I(N__47642));
    Odrv4 I__9549 (
            .O(N__47642),
            .I(\CONTROL.addrstackZ0Z_1 ));
    InMux I__9548 (
            .O(N__47639),
            .I(N__47636));
    LocalMux I__9547 (
            .O(N__47636),
            .I(N__47632));
    InMux I__9546 (
            .O(N__47635),
            .I(N__47629));
    Odrv4 I__9545 (
            .O(N__47632),
            .I(\CONTROL.dout_reto_3 ));
    LocalMux I__9544 (
            .O(N__47629),
            .I(\CONTROL.dout_reto_3 ));
    CascadeMux I__9543 (
            .O(N__47624),
            .I(\CONTROL.programCounter_ret_1_RNILA8IZ0Z_3_cascade_ ));
    InMux I__9542 (
            .O(N__47621),
            .I(N__47618));
    LocalMux I__9541 (
            .O(N__47618),
            .I(\CONTROL.programCounter_ret_19_RNIEO8JZ0Z_3 ));
    InMux I__9540 (
            .O(N__47615),
            .I(N__47612));
    LocalMux I__9539 (
            .O(N__47612),
            .I(N__47608));
    InMux I__9538 (
            .O(N__47611),
            .I(N__47605));
    Odrv4 I__9537 (
            .O(N__47608),
            .I(\CONTROL.programCounter_1_reto_0 ));
    LocalMux I__9536 (
            .O(N__47605),
            .I(\CONTROL.programCounter_1_reto_0 ));
    InMux I__9535 (
            .O(N__47600),
            .I(N__47597));
    LocalMux I__9534 (
            .O(N__47597),
            .I(N__47594));
    Span12Mux_v I__9533 (
            .O(N__47594),
            .I(N__47591));
    Odrv12 I__9532 (
            .O(N__47591),
            .I(\CONTROL.addrstack_3 ));
    InMux I__9531 (
            .O(N__47588),
            .I(N__47585));
    LocalMux I__9530 (
            .O(N__47585),
            .I(\PROM.ROMDATA.m30 ));
    InMux I__9529 (
            .O(N__47582),
            .I(N__47579));
    LocalMux I__9528 (
            .O(N__47579),
            .I(N__47576));
    Span4Mux_h I__9527 (
            .O(N__47576),
            .I(N__47573));
    Odrv4 I__9526 (
            .O(N__47573),
            .I(\PROM.ROMDATA.m35_1 ));
    InMux I__9525 (
            .O(N__47570),
            .I(N__47567));
    LocalMux I__9524 (
            .O(N__47567),
            .I(\PROM.ROMDATA.m35 ));
    InMux I__9523 (
            .O(N__47564),
            .I(N__47560));
    InMux I__9522 (
            .O(N__47563),
            .I(N__47557));
    LocalMux I__9521 (
            .O(N__47560),
            .I(\CONTROL.programCounter_1_reto_2 ));
    LocalMux I__9520 (
            .O(N__47557),
            .I(\CONTROL.programCounter_1_reto_2 ));
    InMux I__9519 (
            .O(N__47552),
            .I(N__47549));
    LocalMux I__9518 (
            .O(N__47549),
            .I(N__47546));
    Span4Mux_v I__9517 (
            .O(N__47546),
            .I(N__47543));
    Odrv4 I__9516 (
            .O(N__47543),
            .I(\PROM.ROMDATA.m392_am ));
    CascadeMux I__9515 (
            .O(N__47540),
            .I(\PROM.ROMDATA.m163_cascade_ ));
    InMux I__9514 (
            .O(N__47537),
            .I(N__47534));
    LocalMux I__9513 (
            .O(N__47534),
            .I(N__47531));
    Odrv4 I__9512 (
            .O(N__47531),
            .I(\PROM.ROMDATA.m176_x ));
    CascadeMux I__9511 (
            .O(N__47528),
            .I(N__47525));
    InMux I__9510 (
            .O(N__47525),
            .I(N__47518));
    InMux I__9509 (
            .O(N__47524),
            .I(N__47518));
    CascadeMux I__9508 (
            .O(N__47523),
            .I(N__47515));
    LocalMux I__9507 (
            .O(N__47518),
            .I(N__47511));
    InMux I__9506 (
            .O(N__47515),
            .I(N__47508));
    InMux I__9505 (
            .O(N__47514),
            .I(N__47505));
    Span4Mux_v I__9504 (
            .O(N__47511),
            .I(N__47502));
    LocalMux I__9503 (
            .O(N__47508),
            .I(\PROM.ROMDATA.N_543_mux_2 ));
    LocalMux I__9502 (
            .O(N__47505),
            .I(\PROM.ROMDATA.N_543_mux_2 ));
    Odrv4 I__9501 (
            .O(N__47502),
            .I(\PROM.ROMDATA.N_543_mux_2 ));
    CascadeMux I__9500 (
            .O(N__47495),
            .I(N__47491));
    InMux I__9499 (
            .O(N__47494),
            .I(N__47485));
    InMux I__9498 (
            .O(N__47491),
            .I(N__47478));
    InMux I__9497 (
            .O(N__47490),
            .I(N__47478));
    InMux I__9496 (
            .O(N__47489),
            .I(N__47478));
    CascadeMux I__9495 (
            .O(N__47488),
            .I(N__47472));
    LocalMux I__9494 (
            .O(N__47485),
            .I(N__47469));
    LocalMux I__9493 (
            .O(N__47478),
            .I(N__47466));
    InMux I__9492 (
            .O(N__47477),
            .I(N__47463));
    InMux I__9491 (
            .O(N__47476),
            .I(N__47456));
    InMux I__9490 (
            .O(N__47475),
            .I(N__47456));
    InMux I__9489 (
            .O(N__47472),
            .I(N__47456));
    Span4Mux_v I__9488 (
            .O(N__47469),
            .I(N__47453));
    Sp12to4 I__9487 (
            .O(N__47466),
            .I(N__47450));
    LocalMux I__9486 (
            .O(N__47463),
            .I(N__47447));
    LocalMux I__9485 (
            .O(N__47456),
            .I(N__47442));
    Sp12to4 I__9484 (
            .O(N__47453),
            .I(N__47442));
    Span12Mux_v I__9483 (
            .O(N__47450),
            .I(N__47437));
    Span12Mux_h I__9482 (
            .O(N__47447),
            .I(N__47437));
    Span12Mux_h I__9481 (
            .O(N__47442),
            .I(N__47434));
    Odrv12 I__9480 (
            .O(N__47437),
            .I(\PROM.ROMDATA.N_569_mux ));
    Odrv12 I__9479 (
            .O(N__47434),
            .I(\PROM.ROMDATA.N_569_mux ));
    CascadeMux I__9478 (
            .O(N__47429),
            .I(\PROM.ROMDATA.m109_am_1_cascade_ ));
    InMux I__9477 (
            .O(N__47426),
            .I(N__47423));
    LocalMux I__9476 (
            .O(N__47423),
            .I(N__47420));
    Sp12to4 I__9475 (
            .O(N__47420),
            .I(N__47417));
    Span12Mux_v I__9474 (
            .O(N__47417),
            .I(N__47414));
    Span12Mux_h I__9473 (
            .O(N__47414),
            .I(N__47411));
    Odrv12 I__9472 (
            .O(N__47411),
            .I(\CONTROL.addrstack_0 ));
    InMux I__9471 (
            .O(N__47408),
            .I(N__47404));
    InMux I__9470 (
            .O(N__47407),
            .I(N__47400));
    LocalMux I__9469 (
            .O(N__47404),
            .I(N__47397));
    InMux I__9468 (
            .O(N__47403),
            .I(N__47394));
    LocalMux I__9467 (
            .O(N__47400),
            .I(N__47391));
    Sp12to4 I__9466 (
            .O(N__47397),
            .I(N__47388));
    LocalMux I__9465 (
            .O(N__47394),
            .I(N__47383));
    Span4Mux_h I__9464 (
            .O(N__47391),
            .I(N__47383));
    Span12Mux_v I__9463 (
            .O(N__47388),
            .I(N__47380));
    Span4Mux_v I__9462 (
            .O(N__47383),
            .I(N__47377));
    Odrv12 I__9461 (
            .O(N__47380),
            .I(N_415));
    Odrv4 I__9460 (
            .O(N__47377),
            .I(N_415));
    InMux I__9459 (
            .O(N__47372),
            .I(N__47369));
    LocalMux I__9458 (
            .O(N__47369),
            .I(\PROM.ROMDATA.m422_am ));
    CascadeMux I__9457 (
            .O(N__47366),
            .I(\PROM.ROMDATA.m422_bm_cascade_ ));
    CascadeMux I__9456 (
            .O(N__47363),
            .I(N__47360));
    InMux I__9455 (
            .O(N__47360),
            .I(N__47357));
    LocalMux I__9454 (
            .O(N__47357),
            .I(N__47354));
    Span4Mux_h I__9453 (
            .O(N__47354),
            .I(N__47351));
    Span4Mux_v I__9452 (
            .O(N__47351),
            .I(N__47348));
    Odrv4 I__9451 (
            .O(N__47348),
            .I(\PROM.ROMDATA.m381_bm ));
    InMux I__9450 (
            .O(N__47345),
            .I(N__47342));
    LocalMux I__9449 (
            .O(N__47342),
            .I(N__47339));
    Span4Mux_v I__9448 (
            .O(N__47339),
            .I(N__47336));
    Span4Mux_h I__9447 (
            .O(N__47336),
            .I(N__47333));
    Odrv4 I__9446 (
            .O(N__47333),
            .I(\PROM.ROMDATA.m298_am ));
    InMux I__9445 (
            .O(N__47330),
            .I(N__47327));
    LocalMux I__9444 (
            .O(N__47327),
            .I(N__47324));
    Span4Mux_v I__9443 (
            .O(N__47324),
            .I(N__47321));
    Span4Mux_h I__9442 (
            .O(N__47321),
            .I(N__47318));
    Span4Mux_h I__9441 (
            .O(N__47318),
            .I(N__47315));
    Odrv4 I__9440 (
            .O(N__47315),
            .I(\CONTROL.programCounter_1_axb_4 ));
    CascadeMux I__9439 (
            .O(N__47312),
            .I(\PROM.ROMDATA.N_543_mux_2_cascade_ ));
    InMux I__9438 (
            .O(N__47309),
            .I(N__47306));
    LocalMux I__9437 (
            .O(N__47306),
            .I(N__47302));
    InMux I__9436 (
            .O(N__47305),
            .I(N__47299));
    Span4Mux_v I__9435 (
            .O(N__47302),
            .I(N__47296));
    LocalMux I__9434 (
            .O(N__47299),
            .I(N__47293));
    Span4Mux_h I__9433 (
            .O(N__47296),
            .I(N__47288));
    Span4Mux_h I__9432 (
            .O(N__47293),
            .I(N__47288));
    Odrv4 I__9431 (
            .O(N__47288),
            .I(\PROM.ROMDATA.N_559_mux ));
    InMux I__9430 (
            .O(N__47285),
            .I(N__47281));
    InMux I__9429 (
            .O(N__47284),
            .I(N__47278));
    LocalMux I__9428 (
            .O(N__47281),
            .I(N__47268));
    LocalMux I__9427 (
            .O(N__47278),
            .I(N__47265));
    InMux I__9426 (
            .O(N__47277),
            .I(N__47260));
    InMux I__9425 (
            .O(N__47276),
            .I(N__47260));
    InMux I__9424 (
            .O(N__47275),
            .I(N__47255));
    InMux I__9423 (
            .O(N__47274),
            .I(N__47255));
    InMux I__9422 (
            .O(N__47273),
            .I(N__47250));
    InMux I__9421 (
            .O(N__47272),
            .I(N__47250));
    CascadeMux I__9420 (
            .O(N__47271),
            .I(N__47247));
    Span4Mux_h I__9419 (
            .O(N__47268),
            .I(N__47243));
    Span4Mux_h I__9418 (
            .O(N__47265),
            .I(N__47240));
    LocalMux I__9417 (
            .O(N__47260),
            .I(N__47237));
    LocalMux I__9416 (
            .O(N__47255),
            .I(N__47232));
    LocalMux I__9415 (
            .O(N__47250),
            .I(N__47232));
    InMux I__9414 (
            .O(N__47247),
            .I(N__47227));
    InMux I__9413 (
            .O(N__47246),
            .I(N__47227));
    Odrv4 I__9412 (
            .O(N__47243),
            .I(aluOperand1_2));
    Odrv4 I__9411 (
            .O(N__47240),
            .I(aluOperand1_2));
    Odrv4 I__9410 (
            .O(N__47237),
            .I(aluOperand1_2));
    Odrv12 I__9409 (
            .O(N__47232),
            .I(aluOperand1_2));
    LocalMux I__9408 (
            .O(N__47227),
            .I(aluOperand1_2));
    CascadeMux I__9407 (
            .O(N__47216),
            .I(\ALU.dout_6_ns_1_14_cascade_ ));
    InMux I__9406 (
            .O(N__47213),
            .I(N__47205));
    InMux I__9405 (
            .O(N__47212),
            .I(N__47205));
    InMux I__9404 (
            .O(N__47211),
            .I(N__47196));
    InMux I__9403 (
            .O(N__47210),
            .I(N__47196));
    LocalMux I__9402 (
            .O(N__47205),
            .I(N__47185));
    InMux I__9401 (
            .O(N__47204),
            .I(N__47180));
    InMux I__9400 (
            .O(N__47203),
            .I(N__47180));
    InMux I__9399 (
            .O(N__47202),
            .I(N__47175));
    InMux I__9398 (
            .O(N__47201),
            .I(N__47175));
    LocalMux I__9397 (
            .O(N__47196),
            .I(N__47172));
    InMux I__9396 (
            .O(N__47195),
            .I(N__47167));
    InMux I__9395 (
            .O(N__47194),
            .I(N__47167));
    InMux I__9394 (
            .O(N__47193),
            .I(N__47162));
    InMux I__9393 (
            .O(N__47192),
            .I(N__47162));
    InMux I__9392 (
            .O(N__47191),
            .I(N__47157));
    InMux I__9391 (
            .O(N__47190),
            .I(N__47157));
    InMux I__9390 (
            .O(N__47189),
            .I(N__47152));
    InMux I__9389 (
            .O(N__47188),
            .I(N__47152));
    Span4Mux_h I__9388 (
            .O(N__47185),
            .I(N__47149));
    LocalMux I__9387 (
            .O(N__47180),
            .I(N__47146));
    LocalMux I__9386 (
            .O(N__47175),
            .I(N__47139));
    Span4Mux_h I__9385 (
            .O(N__47172),
            .I(N__47136));
    LocalMux I__9384 (
            .O(N__47167),
            .I(N__47133));
    LocalMux I__9383 (
            .O(N__47162),
            .I(N__47128));
    LocalMux I__9382 (
            .O(N__47157),
            .I(N__47128));
    LocalMux I__9381 (
            .O(N__47152),
            .I(N__47121));
    Span4Mux_v I__9380 (
            .O(N__47149),
            .I(N__47121));
    Span4Mux_h I__9379 (
            .O(N__47146),
            .I(N__47121));
    InMux I__9378 (
            .O(N__47145),
            .I(N__47112));
    InMux I__9377 (
            .O(N__47144),
            .I(N__47112));
    InMux I__9376 (
            .O(N__47143),
            .I(N__47112));
    InMux I__9375 (
            .O(N__47142),
            .I(N__47112));
    Odrv4 I__9374 (
            .O(N__47139),
            .I(aluOperand1_1));
    Odrv4 I__9373 (
            .O(N__47136),
            .I(aluOperand1_1));
    Odrv4 I__9372 (
            .O(N__47133),
            .I(aluOperand1_1));
    Odrv12 I__9371 (
            .O(N__47128),
            .I(aluOperand1_1));
    Odrv4 I__9370 (
            .O(N__47121),
            .I(aluOperand1_1));
    LocalMux I__9369 (
            .O(N__47112),
            .I(aluOperand1_1));
    InMux I__9368 (
            .O(N__47099),
            .I(N__47096));
    LocalMux I__9367 (
            .O(N__47096),
            .I(\ALU.N_1099 ));
    CascadeMux I__9366 (
            .O(N__47093),
            .I(\ALU.N_1147_cascade_ ));
    InMux I__9365 (
            .O(N__47090),
            .I(N__47087));
    LocalMux I__9364 (
            .O(N__47087),
            .I(N__47084));
    Span4Mux_v I__9363 (
            .O(N__47084),
            .I(N__47081));
    Sp12to4 I__9362 (
            .O(N__47081),
            .I(N__47078));
    Odrv12 I__9361 (
            .O(N__47078),
            .I(DROM_ROMDATA_dintern_14ro));
    CascadeMux I__9360 (
            .O(N__47075),
            .I(aluOut_14_cascade_));
    InMux I__9359 (
            .O(N__47072),
            .I(N__47069));
    LocalMux I__9358 (
            .O(N__47069),
            .I(N__47066));
    Span4Mux_h I__9357 (
            .O(N__47066),
            .I(N__47063));
    Span4Mux_h I__9356 (
            .O(N__47063),
            .I(N__47059));
    InMux I__9355 (
            .O(N__47062),
            .I(N__47056));
    Odrv4 I__9354 (
            .O(N__47059),
            .I(N_207));
    LocalMux I__9353 (
            .O(N__47056),
            .I(N_207));
    InMux I__9352 (
            .O(N__47051),
            .I(N__47047));
    InMux I__9351 (
            .O(N__47050),
            .I(N__47044));
    LocalMux I__9350 (
            .O(N__47047),
            .I(N__47040));
    LocalMux I__9349 (
            .O(N__47044),
            .I(N__47037));
    InMux I__9348 (
            .O(N__47043),
            .I(N__47034));
    Span4Mux_h I__9347 (
            .O(N__47040),
            .I(N__47030));
    Span4Mux_h I__9346 (
            .O(N__47037),
            .I(N__47025));
    LocalMux I__9345 (
            .O(N__47034),
            .I(N__47025));
    InMux I__9344 (
            .O(N__47033),
            .I(N__47022));
    Odrv4 I__9343 (
            .O(N__47030),
            .I(\CONTROL.un1_busState114_2_0_o2_0_0 ));
    Odrv4 I__9342 (
            .O(N__47025),
            .I(\CONTROL.un1_busState114_2_0_o2_0_0 ));
    LocalMux I__9341 (
            .O(N__47022),
            .I(\CONTROL.un1_busState114_2_0_o2_0_0 ));
    InMux I__9340 (
            .O(N__47015),
            .I(N__47012));
    LocalMux I__9339 (
            .O(N__47012),
            .I(N__47006));
    InMux I__9338 (
            .O(N__47011),
            .I(N__47003));
    InMux I__9337 (
            .O(N__47010),
            .I(N__46997));
    InMux I__9336 (
            .O(N__47009),
            .I(N__46997));
    Span4Mux_v I__9335 (
            .O(N__47006),
            .I(N__46994));
    LocalMux I__9334 (
            .O(N__47003),
            .I(N__46991));
    InMux I__9333 (
            .O(N__47002),
            .I(N__46988));
    LocalMux I__9332 (
            .O(N__46997),
            .I(N__46985));
    Span4Mux_v I__9331 (
            .O(N__46994),
            .I(N__46981));
    Span4Mux_h I__9330 (
            .O(N__46991),
            .I(N__46974));
    LocalMux I__9329 (
            .O(N__46988),
            .I(N__46974));
    Span4Mux_v I__9328 (
            .O(N__46985),
            .I(N__46974));
    InMux I__9327 (
            .O(N__46984),
            .I(N__46971));
    Odrv4 I__9326 (
            .O(N__46981),
            .I(\CONTROL.N_361_1 ));
    Odrv4 I__9325 (
            .O(N__46974),
            .I(\CONTROL.N_361_1 ));
    LocalMux I__9324 (
            .O(N__46971),
            .I(\CONTROL.N_361_1 ));
    CascadeMux I__9323 (
            .O(N__46964),
            .I(N__46961));
    InMux I__9322 (
            .O(N__46961),
            .I(N__46958));
    LocalMux I__9321 (
            .O(N__46958),
            .I(N__46955));
    Span4Mux_h I__9320 (
            .O(N__46955),
            .I(N__46952));
    Span4Mux_h I__9319 (
            .O(N__46952),
            .I(N__46949));
    Odrv4 I__9318 (
            .O(N__46949),
            .I(\CONTROL.un1_busState114_2_0_0_0 ));
    InMux I__9317 (
            .O(N__46946),
            .I(N__46939));
    CascadeMux I__9316 (
            .O(N__46945),
            .I(N__46936));
    InMux I__9315 (
            .O(N__46944),
            .I(N__46932));
    InMux I__9314 (
            .O(N__46943),
            .I(N__46927));
    InMux I__9313 (
            .O(N__46942),
            .I(N__46927));
    LocalMux I__9312 (
            .O(N__46939),
            .I(N__46919));
    InMux I__9311 (
            .O(N__46936),
            .I(N__46914));
    InMux I__9310 (
            .O(N__46935),
            .I(N__46914));
    LocalMux I__9309 (
            .O(N__46932),
            .I(N__46909));
    LocalMux I__9308 (
            .O(N__46927),
            .I(N__46909));
    InMux I__9307 (
            .O(N__46926),
            .I(N__46904));
    InMux I__9306 (
            .O(N__46925),
            .I(N__46904));
    InMux I__9305 (
            .O(N__46924),
            .I(N__46899));
    InMux I__9304 (
            .O(N__46923),
            .I(N__46899));
    CascadeMux I__9303 (
            .O(N__46922),
            .I(N__46893));
    Span4Mux_v I__9302 (
            .O(N__46919),
            .I(N__46889));
    LocalMux I__9301 (
            .O(N__46914),
            .I(N__46884));
    Span4Mux_h I__9300 (
            .O(N__46909),
            .I(N__46884));
    LocalMux I__9299 (
            .O(N__46904),
            .I(N__46881));
    LocalMux I__9298 (
            .O(N__46899),
            .I(N__46878));
    InMux I__9297 (
            .O(N__46898),
            .I(N__46871));
    InMux I__9296 (
            .O(N__46897),
            .I(N__46871));
    InMux I__9295 (
            .O(N__46896),
            .I(N__46871));
    InMux I__9294 (
            .O(N__46893),
            .I(N__46866));
    InMux I__9293 (
            .O(N__46892),
            .I(N__46866));
    Span4Mux_h I__9292 (
            .O(N__46889),
            .I(N__46859));
    Span4Mux_h I__9291 (
            .O(N__46884),
            .I(N__46859));
    Span4Mux_v I__9290 (
            .O(N__46881),
            .I(N__46859));
    Odrv4 I__9289 (
            .O(N__46878),
            .I(aluOperand2_2_rep2));
    LocalMux I__9288 (
            .O(N__46871),
            .I(aluOperand2_2_rep2));
    LocalMux I__9287 (
            .O(N__46866),
            .I(aluOperand2_2_rep2));
    Odrv4 I__9286 (
            .O(N__46859),
            .I(aluOperand2_2_rep2));
    InMux I__9285 (
            .O(N__46850),
            .I(N__46847));
    LocalMux I__9284 (
            .O(N__46847),
            .I(\ALU.c_RNI9SHFZ0Z_14 ));
    CascadeMux I__9283 (
            .O(N__46844),
            .I(\ALU.a_RNI5CPUZ0Z_14_cascade_ ));
    InMux I__9282 (
            .O(N__46841),
            .I(N__46837));
    InMux I__9281 (
            .O(N__46840),
            .I(N__46833));
    LocalMux I__9280 (
            .O(N__46837),
            .I(N__46828));
    InMux I__9279 (
            .O(N__46836),
            .I(N__46824));
    LocalMux I__9278 (
            .O(N__46833),
            .I(N__46821));
    InMux I__9277 (
            .O(N__46832),
            .I(N__46816));
    InMux I__9276 (
            .O(N__46831),
            .I(N__46816));
    Span4Mux_h I__9275 (
            .O(N__46828),
            .I(N__46808));
    InMux I__9274 (
            .O(N__46827),
            .I(N__46805));
    LocalMux I__9273 (
            .O(N__46824),
            .I(N__46798));
    Span4Mux_h I__9272 (
            .O(N__46821),
            .I(N__46798));
    LocalMux I__9271 (
            .O(N__46816),
            .I(N__46798));
    InMux I__9270 (
            .O(N__46815),
            .I(N__46789));
    InMux I__9269 (
            .O(N__46814),
            .I(N__46789));
    InMux I__9268 (
            .O(N__46813),
            .I(N__46789));
    InMux I__9267 (
            .O(N__46812),
            .I(N__46789));
    InMux I__9266 (
            .O(N__46811),
            .I(N__46786));
    Span4Mux_h I__9265 (
            .O(N__46808),
            .I(N__46783));
    LocalMux I__9264 (
            .O(N__46805),
            .I(N__46776));
    Span4Mux_h I__9263 (
            .O(N__46798),
            .I(N__46773));
    LocalMux I__9262 (
            .O(N__46789),
            .I(N__46770));
    LocalMux I__9261 (
            .O(N__46786),
            .I(N__46767));
    Span4Mux_h I__9260 (
            .O(N__46783),
            .I(N__46764));
    InMux I__9259 (
            .O(N__46782),
            .I(N__46761));
    InMux I__9258 (
            .O(N__46781),
            .I(N__46756));
    InMux I__9257 (
            .O(N__46780),
            .I(N__46756));
    InMux I__9256 (
            .O(N__46779),
            .I(N__46753));
    Span4Mux_h I__9255 (
            .O(N__46776),
            .I(N__46746));
    Span4Mux_h I__9254 (
            .O(N__46773),
            .I(N__46746));
    Span4Mux_h I__9253 (
            .O(N__46770),
            .I(N__46746));
    Odrv12 I__9252 (
            .O(N__46767),
            .I(aluOperand2_1));
    Odrv4 I__9251 (
            .O(N__46764),
            .I(aluOperand2_1));
    LocalMux I__9250 (
            .O(N__46761),
            .I(aluOperand2_1));
    LocalMux I__9249 (
            .O(N__46756),
            .I(aluOperand2_1));
    LocalMux I__9248 (
            .O(N__46753),
            .I(aluOperand2_1));
    Odrv4 I__9247 (
            .O(N__46746),
            .I(aluOperand2_1));
    InMux I__9246 (
            .O(N__46733),
            .I(N__46730));
    LocalMux I__9245 (
            .O(N__46730),
            .I(N__46727));
    Odrv12 I__9244 (
            .O(N__46727),
            .I(\ALU.d_RNICJCTZ0Z_14 ));
    CascadeMux I__9243 (
            .O(N__46724),
            .I(\ALU.operand2_7_ns_1_14_cascade_ ));
    InMux I__9242 (
            .O(N__46721),
            .I(N__46718));
    LocalMux I__9241 (
            .O(N__46718),
            .I(N__46715));
    Odrv4 I__9240 (
            .O(N__46715),
            .I(\ALU.b_RNI83KC1Z0Z_14 ));
    InMux I__9239 (
            .O(N__46712),
            .I(N__46709));
    LocalMux I__9238 (
            .O(N__46709),
            .I(N__46706));
    Span4Mux_h I__9237 (
            .O(N__46706),
            .I(N__46703));
    Odrv4 I__9236 (
            .O(N__46703),
            .I(N_191));
    CascadeMux I__9235 (
            .O(N__46700),
            .I(\ALU.operand2_14_cascade_ ));
    CascadeMux I__9234 (
            .O(N__46697),
            .I(N__46694));
    InMux I__9233 (
            .O(N__46694),
            .I(N__46691));
    LocalMux I__9232 (
            .O(N__46691),
            .I(\ALU.d_RNINISC7Z0Z_14 ));
    CascadeMux I__9231 (
            .O(N__46688),
            .I(\ALU.dout_3_ns_1_14_cascade_ ));
    InMux I__9230 (
            .O(N__46685),
            .I(N__46679));
    InMux I__9229 (
            .O(N__46684),
            .I(N__46679));
    LocalMux I__9228 (
            .O(N__46679),
            .I(N__46676));
    Span4Mux_h I__9227 (
            .O(N__46676),
            .I(N__46673));
    Span4Mux_h I__9226 (
            .O(N__46673),
            .I(N__46670));
    Odrv4 I__9225 (
            .O(N__46670),
            .I(\ALU.cZ0Z_15 ));
    InMux I__9224 (
            .O(N__46667),
            .I(N__46664));
    LocalMux I__9223 (
            .O(N__46664),
            .I(N__46661));
    Span4Mux_v I__9222 (
            .O(N__46661),
            .I(N__46658));
    Span4Mux_h I__9221 (
            .O(N__46658),
            .I(N__46655));
    Span4Mux_h I__9220 (
            .O(N__46655),
            .I(N__46651));
    InMux I__9219 (
            .O(N__46654),
            .I(N__46648));
    Odrv4 I__9218 (
            .O(N__46651),
            .I(\ALU.cZ0Z_9 ));
    LocalMux I__9217 (
            .O(N__46648),
            .I(\ALU.cZ0Z_9 ));
    CascadeMux I__9216 (
            .O(N__46643),
            .I(\ALU.log_1_7_cascade_ ));
    InMux I__9215 (
            .O(N__46640),
            .I(N__46637));
    LocalMux I__9214 (
            .O(N__46637),
            .I(N__46634));
    Span4Mux_v I__9213 (
            .O(N__46634),
            .I(N__46631));
    Span4Mux_h I__9212 (
            .O(N__46631),
            .I(N__46628));
    Odrv4 I__9211 (
            .O(N__46628),
            .I(\ALU.mult_7 ));
    CascadeMux I__9210 (
            .O(N__46625),
            .I(\ALU.mult_492_c_RNIQ5BZ0Z457_cascade_ ));
    InMux I__9209 (
            .O(N__46622),
            .I(N__46619));
    LocalMux I__9208 (
            .O(N__46619),
            .I(N__46616));
    Odrv12 I__9207 (
            .O(N__46616),
            .I(\ALU.lshift_7 ));
    CascadeMux I__9206 (
            .O(N__46613),
            .I(\ALU.mult_492_c_RNIGN2JECZ0_cascade_ ));
    InMux I__9205 (
            .O(N__46610),
            .I(N__46606));
    CascadeMux I__9204 (
            .O(N__46609),
            .I(N__46603));
    LocalMux I__9203 (
            .O(N__46606),
            .I(N__46600));
    InMux I__9202 (
            .O(N__46603),
            .I(N__46597));
    Span4Mux_h I__9201 (
            .O(N__46600),
            .I(N__46594));
    LocalMux I__9200 (
            .O(N__46597),
            .I(N__46591));
    Odrv4 I__9199 (
            .O(N__46594),
            .I(\ALU.aZ0Z_7 ));
    Odrv4 I__9198 (
            .O(N__46591),
            .I(\ALU.aZ0Z_7 ));
    CascadeMux I__9197 (
            .O(N__46586),
            .I(N__46583));
    InMux I__9196 (
            .O(N__46583),
            .I(N__46580));
    LocalMux I__9195 (
            .O(N__46580),
            .I(N__46577));
    Span4Mux_h I__9194 (
            .O(N__46577),
            .I(N__46574));
    Span4Mux_v I__9193 (
            .O(N__46574),
            .I(N__46571));
    Span4Mux_h I__9192 (
            .O(N__46571),
            .I(N__46568));
    Odrv4 I__9191 (
            .O(N__46568),
            .I(\ALU.d_RNIO75BGZ0Z_7 ));
    InMux I__9190 (
            .O(N__46565),
            .I(N__46562));
    LocalMux I__9189 (
            .O(N__46562),
            .I(N__46559));
    Span4Mux_h I__9188 (
            .O(N__46559),
            .I(N__46556));
    Odrv4 I__9187 (
            .O(N__46556),
            .I(\ALU.c_RNIE4B6N4Z0Z_15 ));
    CascadeMux I__9186 (
            .O(N__46553),
            .I(\ALU.a_15_1_15_cascade_ ));
    InMux I__9185 (
            .O(N__46550),
            .I(N__46546));
    InMux I__9184 (
            .O(N__46549),
            .I(N__46543));
    LocalMux I__9183 (
            .O(N__46546),
            .I(N__46538));
    LocalMux I__9182 (
            .O(N__46543),
            .I(N__46538));
    Span4Mux_v I__9181 (
            .O(N__46538),
            .I(N__46535));
    Span4Mux_h I__9180 (
            .O(N__46535),
            .I(N__46532));
    Sp12to4 I__9179 (
            .O(N__46532),
            .I(N__46529));
    Span12Mux_v I__9178 (
            .O(N__46529),
            .I(N__46526));
    Odrv12 I__9177 (
            .O(N__46526),
            .I(\ALU.aZ0Z_15 ));
    InMux I__9176 (
            .O(N__46523),
            .I(N__46520));
    LocalMux I__9175 (
            .O(N__46520),
            .I(\ALU.N_812 ));
    CascadeMux I__9174 (
            .O(N__46517),
            .I(\ALU.N_812_cascade_ ));
    InMux I__9173 (
            .O(N__46514),
            .I(N__46511));
    LocalMux I__9172 (
            .O(N__46511),
            .I(\ALU.addsub_cry_14_c_RNI134CVZ0Z5 ));
    CascadeMux I__9171 (
            .O(N__46508),
            .I(N__46505));
    InMux I__9170 (
            .O(N__46505),
            .I(N__46502));
    LocalMux I__9169 (
            .O(N__46502),
            .I(N__46497));
    InMux I__9168 (
            .O(N__46501),
            .I(N__46494));
    InMux I__9167 (
            .O(N__46500),
            .I(N__46491));
    Span4Mux_h I__9166 (
            .O(N__46497),
            .I(N__46488));
    LocalMux I__9165 (
            .O(N__46494),
            .I(\ALU.N_635 ));
    LocalMux I__9164 (
            .O(N__46491),
            .I(\ALU.N_635 ));
    Odrv4 I__9163 (
            .O(N__46488),
            .I(\ALU.N_635 ));
    CascadeMux I__9162 (
            .O(N__46481),
            .I(N__46478));
    InMux I__9161 (
            .O(N__46478),
            .I(N__46472));
    InMux I__9160 (
            .O(N__46477),
            .I(N__46472));
    LocalMux I__9159 (
            .O(N__46472),
            .I(N__46469));
    Span4Mux_v I__9158 (
            .O(N__46469),
            .I(N__46466));
    Odrv4 I__9157 (
            .O(N__46466),
            .I(\ALU.N_639 ));
    InMux I__9156 (
            .O(N__46463),
            .I(N__46459));
    InMux I__9155 (
            .O(N__46462),
            .I(N__46456));
    LocalMux I__9154 (
            .O(N__46459),
            .I(N__46453));
    LocalMux I__9153 (
            .O(N__46456),
            .I(N__46450));
    Span4Mux_v I__9152 (
            .O(N__46453),
            .I(N__46447));
    Span4Mux_h I__9151 (
            .O(N__46450),
            .I(N__46444));
    Span4Mux_h I__9150 (
            .O(N__46447),
            .I(N__46441));
    Span4Mux_h I__9149 (
            .O(N__46444),
            .I(N__46438));
    Odrv4 I__9148 (
            .O(N__46441),
            .I(\ALU.cZ0Z_1 ));
    Odrv4 I__9147 (
            .O(N__46438),
            .I(\ALU.cZ0Z_1 ));
    InMux I__9146 (
            .O(N__46433),
            .I(N__46430));
    LocalMux I__9145 (
            .O(N__46430),
            .I(N__46426));
    InMux I__9144 (
            .O(N__46429),
            .I(N__46423));
    Span4Mux_h I__9143 (
            .O(N__46426),
            .I(N__46420));
    LocalMux I__9142 (
            .O(N__46423),
            .I(N__46417));
    Span4Mux_h I__9141 (
            .O(N__46420),
            .I(N__46414));
    Span4Mux_h I__9140 (
            .O(N__46417),
            .I(N__46411));
    Span4Mux_v I__9139 (
            .O(N__46414),
            .I(N__46408));
    Odrv4 I__9138 (
            .O(N__46411),
            .I(\ALU.cZ0Z_0 ));
    Odrv4 I__9137 (
            .O(N__46408),
            .I(\ALU.cZ0Z_0 ));
    InMux I__9136 (
            .O(N__46403),
            .I(N__46399));
    InMux I__9135 (
            .O(N__46402),
            .I(N__46396));
    LocalMux I__9134 (
            .O(N__46399),
            .I(N__46393));
    LocalMux I__9133 (
            .O(N__46396),
            .I(N__46390));
    Span4Mux_v I__9132 (
            .O(N__46393),
            .I(N__46387));
    Span4Mux_v I__9131 (
            .O(N__46390),
            .I(N__46382));
    Span4Mux_h I__9130 (
            .O(N__46387),
            .I(N__46382));
    Odrv4 I__9129 (
            .O(N__46382),
            .I(\ALU.cZ0Z_7 ));
    InMux I__9128 (
            .O(N__46379),
            .I(N__46373));
    InMux I__9127 (
            .O(N__46378),
            .I(N__46373));
    LocalMux I__9126 (
            .O(N__46373),
            .I(N__46370));
    Span4Mux_h I__9125 (
            .O(N__46370),
            .I(N__46367));
    Span4Mux_h I__9124 (
            .O(N__46367),
            .I(N__46364));
    Span4Mux_h I__9123 (
            .O(N__46364),
            .I(N__46361));
    Odrv4 I__9122 (
            .O(N__46361),
            .I(\ALU.cZ0Z_8 ));
    CascadeMux I__9121 (
            .O(N__46358),
            .I(N__46355));
    InMux I__9120 (
            .O(N__46355),
            .I(N__46352));
    LocalMux I__9119 (
            .O(N__46352),
            .I(N__46348));
    CascadeMux I__9118 (
            .O(N__46351),
            .I(N__46345));
    Span4Mux_h I__9117 (
            .O(N__46348),
            .I(N__46342));
    InMux I__9116 (
            .O(N__46345),
            .I(N__46339));
    Span4Mux_v I__9115 (
            .O(N__46342),
            .I(N__46334));
    LocalMux I__9114 (
            .O(N__46339),
            .I(N__46334));
    Span4Mux_v I__9113 (
            .O(N__46334),
            .I(N__46331));
    Span4Mux_h I__9112 (
            .O(N__46331),
            .I(N__46328));
    Odrv4 I__9111 (
            .O(N__46328),
            .I(\ALU.eZ0Z_1 ));
    InMux I__9110 (
            .O(N__46325),
            .I(N__46321));
    InMux I__9109 (
            .O(N__46324),
            .I(N__46318));
    LocalMux I__9108 (
            .O(N__46321),
            .I(N__46315));
    LocalMux I__9107 (
            .O(N__46318),
            .I(N__46312));
    Span4Mux_v I__9106 (
            .O(N__46315),
            .I(N__46307));
    Span4Mux_h I__9105 (
            .O(N__46312),
            .I(N__46307));
    Span4Mux_h I__9104 (
            .O(N__46307),
            .I(N__46304));
    Span4Mux_v I__9103 (
            .O(N__46304),
            .I(N__46301));
    Odrv4 I__9102 (
            .O(N__46301),
            .I(\ALU.eZ0Z_0 ));
    CascadeMux I__9101 (
            .O(N__46298),
            .I(N__46295));
    InMux I__9100 (
            .O(N__46295),
            .I(N__46289));
    InMux I__9099 (
            .O(N__46294),
            .I(N__46289));
    LocalMux I__9098 (
            .O(N__46289),
            .I(N__46286));
    Sp12to4 I__9097 (
            .O(N__46286),
            .I(N__46283));
    Odrv12 I__9096 (
            .O(N__46283),
            .I(\ALU.eZ0Z_7 ));
    InMux I__9095 (
            .O(N__46280),
            .I(N__46276));
    CascadeMux I__9094 (
            .O(N__46279),
            .I(N__46273));
    LocalMux I__9093 (
            .O(N__46276),
            .I(N__46270));
    InMux I__9092 (
            .O(N__46273),
            .I(N__46267));
    Span4Mux_h I__9091 (
            .O(N__46270),
            .I(N__46264));
    LocalMux I__9090 (
            .O(N__46267),
            .I(N__46261));
    Span4Mux_v I__9089 (
            .O(N__46264),
            .I(N__46258));
    Span4Mux_v I__9088 (
            .O(N__46261),
            .I(N__46255));
    Span4Mux_h I__9087 (
            .O(N__46258),
            .I(N__46252));
    Span4Mux_h I__9086 (
            .O(N__46255),
            .I(N__46249));
    Sp12to4 I__9085 (
            .O(N__46252),
            .I(N__46246));
    Span4Mux_h I__9084 (
            .O(N__46249),
            .I(N__46243));
    Odrv12 I__9083 (
            .O(N__46246),
            .I(\ALU.eZ0Z_8 ));
    Odrv4 I__9082 (
            .O(N__46243),
            .I(\ALU.eZ0Z_8 ));
    CascadeMux I__9081 (
            .O(N__46238),
            .I(N__46234));
    CascadeMux I__9080 (
            .O(N__46237),
            .I(N__46231));
    InMux I__9079 (
            .O(N__46234),
            .I(N__46228));
    InMux I__9078 (
            .O(N__46231),
            .I(N__46225));
    LocalMux I__9077 (
            .O(N__46228),
            .I(N__46220));
    LocalMux I__9076 (
            .O(N__46225),
            .I(N__46220));
    Span4Mux_v I__9075 (
            .O(N__46220),
            .I(N__46217));
    Span4Mux_h I__9074 (
            .O(N__46217),
            .I(N__46214));
    Odrv4 I__9073 (
            .O(N__46214),
            .I(\ALU.eZ0Z_15 ));
    CascadeMux I__9072 (
            .O(N__46211),
            .I(N__46208));
    InMux I__9071 (
            .O(N__46208),
            .I(N__46204));
    InMux I__9070 (
            .O(N__46207),
            .I(N__46201));
    LocalMux I__9069 (
            .O(N__46204),
            .I(N__46198));
    LocalMux I__9068 (
            .O(N__46201),
            .I(N__46195));
    Span4Mux_v I__9067 (
            .O(N__46198),
            .I(N__46192));
    Span4Mux_v I__9066 (
            .O(N__46195),
            .I(N__46189));
    Span4Mux_h I__9065 (
            .O(N__46192),
            .I(N__46186));
    Span4Mux_h I__9064 (
            .O(N__46189),
            .I(N__46183));
    Odrv4 I__9063 (
            .O(N__46186),
            .I(\ALU.eZ0Z_9 ));
    Odrv4 I__9062 (
            .O(N__46183),
            .I(\ALU.eZ0Z_9 ));
    InMux I__9061 (
            .O(N__46178),
            .I(N__46175));
    LocalMux I__9060 (
            .O(N__46175),
            .I(N__46172));
    Span4Mux_h I__9059 (
            .O(N__46172),
            .I(N__46169));
    Span4Mux_v I__9058 (
            .O(N__46169),
            .I(N__46166));
    Odrv4 I__9057 (
            .O(N__46166),
            .I(\ALU.N_647 ));
    InMux I__9056 (
            .O(N__46163),
            .I(N__46160));
    LocalMux I__9055 (
            .O(N__46160),
            .I(N__46156));
    InMux I__9054 (
            .O(N__46159),
            .I(N__46153));
    Span4Mux_h I__9053 (
            .O(N__46156),
            .I(N__46150));
    LocalMux I__9052 (
            .O(N__46153),
            .I(N__46147));
    Span4Mux_h I__9051 (
            .O(N__46150),
            .I(N__46144));
    Odrv12 I__9050 (
            .O(N__46147),
            .I(\ALU.N_643 ));
    Odrv4 I__9049 (
            .O(N__46144),
            .I(\ALU.N_643 ));
    InMux I__9048 (
            .O(N__46139),
            .I(N__46136));
    LocalMux I__9047 (
            .O(N__46136),
            .I(\ALU.N_707 ));
    CascadeMux I__9046 (
            .O(N__46133),
            .I(\ALU.addsub_cry_14_c_RNI134CV5Z0Z_0_cascade_ ));
    CascadeMux I__9045 (
            .O(N__46130),
            .I(\ALU.addsub_cry_14_c_RNIKS9S5HZ0_cascade_ ));
    InMux I__9044 (
            .O(N__46127),
            .I(N__46124));
    LocalMux I__9043 (
            .O(N__46124),
            .I(\ALU.mult_335_c_RNOZ0Z_0 ));
    CascadeMux I__9042 (
            .O(N__46121),
            .I(\ALU.N_835_cascade_ ));
    InMux I__9041 (
            .O(N__46118),
            .I(N__46114));
    CascadeMux I__9040 (
            .O(N__46117),
            .I(N__46111));
    LocalMux I__9039 (
            .O(N__46114),
            .I(N__46108));
    InMux I__9038 (
            .O(N__46111),
            .I(N__46105));
    Odrv4 I__9037 (
            .O(N__46108),
            .I(\ALU.N_852 ));
    LocalMux I__9036 (
            .O(N__46105),
            .I(\ALU.N_852 ));
    CascadeMux I__9035 (
            .O(N__46100),
            .I(\ALU.rshift_7_ns_1_7_cascade_ ));
    CascadeMux I__9034 (
            .O(N__46097),
            .I(\ALU.N_925_cascade_ ));
    CascadeMux I__9033 (
            .O(N__46094),
            .I(N__46091));
    InMux I__9032 (
            .O(N__46091),
            .I(N__46088));
    LocalMux I__9031 (
            .O(N__46088),
            .I(N__46085));
    Span4Mux_v I__9030 (
            .O(N__46085),
            .I(N__46082));
    Sp12to4 I__9029 (
            .O(N__46082),
            .I(N__46079));
    Odrv12 I__9028 (
            .O(N__46079),
            .I(\ALU.N_833 ));
    InMux I__9027 (
            .O(N__46076),
            .I(N__46070));
    InMux I__9026 (
            .O(N__46075),
            .I(N__46070));
    LocalMux I__9025 (
            .O(N__46070),
            .I(N__46067));
    Span4Mux_h I__9024 (
            .O(N__46067),
            .I(N__46063));
    InMux I__9023 (
            .O(N__46066),
            .I(N__46060));
    Odrv4 I__9022 (
            .O(N__46063),
            .I(\ALU.N_837 ));
    LocalMux I__9021 (
            .O(N__46060),
            .I(\ALU.N_837 ));
    CascadeMux I__9020 (
            .O(N__46055),
            .I(\ALU.rshift_7_ns_1_3_cascade_ ));
    InMux I__9019 (
            .O(N__46052),
            .I(N__46049));
    LocalMux I__9018 (
            .O(N__46049),
            .I(N__46046));
    Odrv4 I__9017 (
            .O(N__46046),
            .I(\ALU.N_921 ));
    IoInMux I__9016 (
            .O(N__46043),
            .I(N__46040));
    LocalMux I__9015 (
            .O(N__46040),
            .I(N__46036));
    IoInMux I__9014 (
            .O(N__46039),
            .I(N__46033));
    Span4Mux_s0_h I__9013 (
            .O(N__46036),
            .I(N__46029));
    LocalMux I__9012 (
            .O(N__46033),
            .I(N__46026));
    InMux I__9011 (
            .O(N__46032),
            .I(N__46023));
    Span4Mux_h I__9010 (
            .O(N__46029),
            .I(N__46020));
    IoSpan4Mux I__9009 (
            .O(N__46026),
            .I(N__46017));
    LocalMux I__9008 (
            .O(N__46023),
            .I(N__46014));
    Sp12to4 I__9007 (
            .O(N__46020),
            .I(N__46011));
    Span4Mux_s3_h I__9006 (
            .O(N__46017),
            .I(N__46008));
    Span4Mux_v I__9005 (
            .O(N__46014),
            .I(N__46005));
    Span12Mux_v I__9004 (
            .O(N__46011),
            .I(N__46002));
    Sp12to4 I__9003 (
            .O(N__46008),
            .I(N__45999));
    Span4Mux_v I__9002 (
            .O(N__46005),
            .I(N__45996));
    Span12Mux_h I__9001 (
            .O(N__46002),
            .I(N__45991));
    Span12Mux_v I__9000 (
            .O(N__45999),
            .I(N__45991));
    Span4Mux_h I__8999 (
            .O(N__45996),
            .I(N__45988));
    Odrv12 I__8998 (
            .O(N__45991),
            .I(bus_7));
    Odrv4 I__8997 (
            .O(N__45988),
            .I(bus_7));
    InMux I__8996 (
            .O(N__45983),
            .I(N__45980));
    LocalMux I__8995 (
            .O(N__45980),
            .I(N__45977));
    Span4Mux_v I__8994 (
            .O(N__45977),
            .I(N__45974));
    Span4Mux_h I__8993 (
            .O(N__45974),
            .I(N__45971));
    Odrv4 I__8992 (
            .O(N__45971),
            .I(\ALU.N_1030 ));
    InMux I__8991 (
            .O(N__45968),
            .I(N__45965));
    LocalMux I__8990 (
            .O(N__45965),
            .I(\ALU.c_RNI08R632Z0Z_15 ));
    InMux I__8989 (
            .O(N__45962),
            .I(N__45959));
    LocalMux I__8988 (
            .O(N__45959),
            .I(N__45956));
    Span4Mux_v I__8987 (
            .O(N__45956),
            .I(N__45953));
    Span4Mux_h I__8986 (
            .O(N__45953),
            .I(N__45950));
    Odrv4 I__8985 (
            .O(N__45950),
            .I(\ALU.lshift_3_ns_1_11 ));
    InMux I__8984 (
            .O(N__45947),
            .I(N__45944));
    LocalMux I__8983 (
            .O(N__45944),
            .I(N__45941));
    Odrv4 I__8982 (
            .O(N__45941),
            .I(\ALU.d_RNI4N3K21Z0Z_8 ));
    CascadeMux I__8981 (
            .O(N__45938),
            .I(N__45935));
    InMux I__8980 (
            .O(N__45935),
            .I(N__45932));
    LocalMux I__8979 (
            .O(N__45932),
            .I(\ALU.d_RNIH8D821Z0Z_8 ));
    CascadeMux I__8978 (
            .O(N__45929),
            .I(N__45926));
    InMux I__8977 (
            .O(N__45926),
            .I(N__45923));
    LocalMux I__8976 (
            .O(N__45923),
            .I(N__45920));
    Odrv4 I__8975 (
            .O(N__45920),
            .I(\ALU.mult_335_c_RNOZ0 ));
    InMux I__8974 (
            .O(N__45917),
            .I(N__45914));
    LocalMux I__8973 (
            .O(N__45914),
            .I(\ALU.c_RNIBQSTOZ0Z_11 ));
    CascadeMux I__8972 (
            .O(N__45911),
            .I(N__45908));
    InMux I__8971 (
            .O(N__45908),
            .I(N__45905));
    LocalMux I__8970 (
            .O(N__45905),
            .I(\ALU.c_RNIG5G6F1Z0Z_10 ));
    CascadeMux I__8969 (
            .O(N__45902),
            .I(N__45899));
    InMux I__8968 (
            .O(N__45899),
            .I(N__45896));
    LocalMux I__8967 (
            .O(N__45896),
            .I(\ALU.mult_11_12 ));
    InMux I__8966 (
            .O(N__45893),
            .I(\ALU.mult_11_c11 ));
    InMux I__8965 (
            .O(N__45890),
            .I(N__45887));
    LocalMux I__8964 (
            .O(N__45887),
            .I(N__45884));
    Span4Mux_h I__8963 (
            .O(N__45884),
            .I(N__45881));
    Odrv4 I__8962 (
            .O(N__45881),
            .I(\ALU.c_RNIN266MZ0Z_11 ));
    CascadeMux I__8961 (
            .O(N__45878),
            .I(N__45875));
    InMux I__8960 (
            .O(N__45875),
            .I(N__45872));
    LocalMux I__8959 (
            .O(N__45872),
            .I(\ALU.c_RNIT73F71Z0Z_10 ));
    CascadeMux I__8958 (
            .O(N__45869),
            .I(N__45866));
    InMux I__8957 (
            .O(N__45866),
            .I(N__45863));
    LocalMux I__8956 (
            .O(N__45863),
            .I(\ALU.mult_11_13 ));
    InMux I__8955 (
            .O(N__45860),
            .I(\ALU.mult_11_c12 ));
    CascadeMux I__8954 (
            .O(N__45857),
            .I(N__45854));
    InMux I__8953 (
            .O(N__45854),
            .I(N__45851));
    LocalMux I__8952 (
            .O(N__45851),
            .I(N__45848));
    Span4Mux_v I__8951 (
            .O(N__45848),
            .I(N__45845));
    Span4Mux_h I__8950 (
            .O(N__45845),
            .I(N__45842));
    Span4Mux_h I__8949 (
            .O(N__45842),
            .I(N__45839));
    Odrv4 I__8948 (
            .O(N__45839),
            .I(\ALU.c_RNIK31N31Z0Z_10 ));
    CascadeMux I__8947 (
            .O(N__45836),
            .I(N__45833));
    InMux I__8946 (
            .O(N__45833),
            .I(N__45830));
    LocalMux I__8945 (
            .O(N__45830),
            .I(\ALU.mult_11_14 ));
    InMux I__8944 (
            .O(N__45827),
            .I(\ALU.mult_11_c13 ));
    InMux I__8943 (
            .O(N__45824),
            .I(\ALU.mult_11_c14 ));
    InMux I__8942 (
            .O(N__45821),
            .I(N__45818));
    LocalMux I__8941 (
            .O(N__45818),
            .I(\ALU.mult_11_c14_THRU_CO ));
    InMux I__8940 (
            .O(N__45815),
            .I(N__45812));
    LocalMux I__8939 (
            .O(N__45812),
            .I(\ALU.c_RNIOSF6HZ0Z_11 ));
    InMux I__8938 (
            .O(N__45809),
            .I(N__45806));
    LocalMux I__8937 (
            .O(N__45806),
            .I(N__45802));
    CascadeMux I__8936 (
            .O(N__45805),
            .I(N__45799));
    Span4Mux_v I__8935 (
            .O(N__45802),
            .I(N__45796));
    InMux I__8934 (
            .O(N__45799),
            .I(N__45793));
    Span4Mux_v I__8933 (
            .O(N__45796),
            .I(N__45790));
    LocalMux I__8932 (
            .O(N__45793),
            .I(\PROM.ROMDATA.m134 ));
    Odrv4 I__8931 (
            .O(N__45790),
            .I(\PROM.ROMDATA.m134 ));
    InMux I__8930 (
            .O(N__45785),
            .I(N__45782));
    LocalMux I__8929 (
            .O(N__45782),
            .I(\PROM.ROMDATA.m396_bm ));
    CascadeMux I__8928 (
            .O(N__45779),
            .I(\PROM.ROMDATA.m396_am_cascade_ ));
    CascadeMux I__8927 (
            .O(N__45776),
            .I(\PROM.ROMDATA.m396_ns_cascade_ ));
    InMux I__8926 (
            .O(N__45773),
            .I(N__45770));
    LocalMux I__8925 (
            .O(N__45770),
            .I(\PROM.ROMDATA.m401_ns_1 ));
    InMux I__8924 (
            .O(N__45767),
            .I(N__45763));
    InMux I__8923 (
            .O(N__45766),
            .I(N__45760));
    LocalMux I__8922 (
            .O(N__45763),
            .I(N__45757));
    LocalMux I__8921 (
            .O(N__45760),
            .I(N__45754));
    Span4Mux_h I__8920 (
            .O(N__45757),
            .I(N__45751));
    Span4Mux_h I__8919 (
            .O(N__45754),
            .I(N__45748));
    Span4Mux_v I__8918 (
            .O(N__45751),
            .I(N__45745));
    Odrv4 I__8917 (
            .O(N__45748),
            .I(\PROM.ROMDATA.m401_ns ));
    Odrv4 I__8916 (
            .O(N__45745),
            .I(\PROM.ROMDATA.m401_ns ));
    CascadeMux I__8915 (
            .O(N__45740),
            .I(N__45737));
    InMux I__8914 (
            .O(N__45737),
            .I(N__45734));
    LocalMux I__8913 (
            .O(N__45734),
            .I(N__45731));
    Odrv4 I__8912 (
            .O(N__45731),
            .I(\ALU.N_607 ));
    InMux I__8911 (
            .O(N__45728),
            .I(N__45725));
    LocalMux I__8910 (
            .O(N__45725),
            .I(N__45720));
    InMux I__8909 (
            .O(N__45724),
            .I(N__45717));
    CascadeMux I__8908 (
            .O(N__45723),
            .I(N__45714));
    Span4Mux_h I__8907 (
            .O(N__45720),
            .I(N__45711));
    LocalMux I__8906 (
            .O(N__45717),
            .I(N__45708));
    InMux I__8905 (
            .O(N__45714),
            .I(N__45705));
    Span4Mux_v I__8904 (
            .O(N__45711),
            .I(N__45702));
    Span4Mux_v I__8903 (
            .O(N__45708),
            .I(N__45699));
    LocalMux I__8902 (
            .O(N__45705),
            .I(N__45696));
    Span4Mux_h I__8901 (
            .O(N__45702),
            .I(N__45693));
    Span4Mux_h I__8900 (
            .O(N__45699),
            .I(N__45690));
    Odrv12 I__8899 (
            .O(N__45696),
            .I(\ALU.N_767 ));
    Odrv4 I__8898 (
            .O(N__45693),
            .I(\ALU.N_767 ));
    Odrv4 I__8897 (
            .O(N__45690),
            .I(\ALU.N_767 ));
    CascadeMux I__8896 (
            .O(N__45683),
            .I(\ALU.N_607_cascade_ ));
    InMux I__8895 (
            .O(N__45680),
            .I(N__45677));
    LocalMux I__8894 (
            .O(N__45677),
            .I(N__45674));
    Span12Mux_v I__8893 (
            .O(N__45674),
            .I(N__45670));
    InMux I__8892 (
            .O(N__45673),
            .I(N__45667));
    Odrv12 I__8891 (
            .O(N__45670),
            .I(\CONTROL.ctrlOut_5 ));
    LocalMux I__8890 (
            .O(N__45667),
            .I(\CONTROL.ctrlOut_5 ));
    InMux I__8889 (
            .O(N__45662),
            .I(N__45659));
    LocalMux I__8888 (
            .O(N__45659),
            .I(N__45655));
    InMux I__8887 (
            .O(N__45658),
            .I(N__45652));
    Span4Mux_v I__8886 (
            .O(N__45655),
            .I(N__45649));
    LocalMux I__8885 (
            .O(N__45652),
            .I(N__45646));
    Odrv4 I__8884 (
            .O(N__45649),
            .I(\CONTROL.dout_reto_5 ));
    Odrv4 I__8883 (
            .O(N__45646),
            .I(\CONTROL.dout_reto_5 ));
    InMux I__8882 (
            .O(N__45641),
            .I(N__45638));
    LocalMux I__8881 (
            .O(N__45638),
            .I(N__45635));
    Odrv12 I__8880 (
            .O(N__45635),
            .I(\CONTROL.programCounter_ret_19_RNIV5IGZ0Z_6 ));
    InMux I__8879 (
            .O(N__45632),
            .I(N__45629));
    LocalMux I__8878 (
            .O(N__45629),
            .I(N__45626));
    Span4Mux_h I__8877 (
            .O(N__45626),
            .I(N__45623));
    Span4Mux_h I__8876 (
            .O(N__45623),
            .I(N__45620));
    Span4Mux_h I__8875 (
            .O(N__45620),
            .I(N__45617));
    Odrv4 I__8874 (
            .O(N__45617),
            .I(\CONTROL.addrstack_6 ));
    InMux I__8873 (
            .O(N__45614),
            .I(N__45610));
    InMux I__8872 (
            .O(N__45613),
            .I(N__45607));
    LocalMux I__8871 (
            .O(N__45610),
            .I(N__45604));
    LocalMux I__8870 (
            .O(N__45607),
            .I(\CONTROL.addrstack_reto_6 ));
    Odrv12 I__8869 (
            .O(N__45604),
            .I(\CONTROL.addrstack_reto_6 ));
    InMux I__8868 (
            .O(N__45599),
            .I(N__45596));
    LocalMux I__8867 (
            .O(N__45596),
            .I(\PROM.ROMDATA.m48 ));
    InMux I__8866 (
            .O(N__45593),
            .I(N__45590));
    LocalMux I__8865 (
            .O(N__45590),
            .I(N__45587));
    Span4Mux_v I__8864 (
            .O(N__45587),
            .I(N__45584));
    Sp12to4 I__8863 (
            .O(N__45584),
            .I(N__45580));
    InMux I__8862 (
            .O(N__45583),
            .I(N__45577));
    Odrv12 I__8861 (
            .O(N__45580),
            .I(\CONTROL.ctrlOut_6 ));
    LocalMux I__8860 (
            .O(N__45577),
            .I(\CONTROL.ctrlOut_6 ));
    InMux I__8859 (
            .O(N__45572),
            .I(N__45569));
    LocalMux I__8858 (
            .O(N__45569),
            .I(\CONTROL.dout_reto_6 ));
    InMux I__8857 (
            .O(N__45566),
            .I(N__45563));
    LocalMux I__8856 (
            .O(N__45563),
            .I(\PROM.ROMDATA.m7 ));
    CascadeMux I__8855 (
            .O(N__45560),
            .I(\PROM.ROMDATA.m392_bm_cascade_ ));
    CascadeMux I__8854 (
            .O(N__45557),
            .I(\PROM.ROMDATA.m392_ns_cascade_ ));
    CascadeMux I__8853 (
            .O(N__45554),
            .I(N__45551));
    InMux I__8852 (
            .O(N__45551),
            .I(N__45548));
    LocalMux I__8851 (
            .O(N__45548),
            .I(N__45545));
    Odrv12 I__8850 (
            .O(N__45545),
            .I(\PROM.ROMDATA.m36 ));
    CascadeMux I__8849 (
            .O(N__45542),
            .I(\PROM.ROMDATA.N_526_mux_cascade_ ));
    InMux I__8848 (
            .O(N__45539),
            .I(N__45536));
    LocalMux I__8847 (
            .O(N__45536),
            .I(N__45533));
    Span4Mux_h I__8846 (
            .O(N__45533),
            .I(N__45530));
    Span4Mux_v I__8845 (
            .O(N__45530),
            .I(N__45527));
    Odrv4 I__8844 (
            .O(N__45527),
            .I(\PROM.ROMDATA.m238_bm ));
    CascadeMux I__8843 (
            .O(N__45524),
            .I(N__45520));
    CascadeMux I__8842 (
            .O(N__45523),
            .I(N__45517));
    InMux I__8841 (
            .O(N__45520),
            .I(N__45510));
    InMux I__8840 (
            .O(N__45517),
            .I(N__45510));
    CascadeMux I__8839 (
            .O(N__45516),
            .I(N__45506));
    CascadeMux I__8838 (
            .O(N__45515),
            .I(N__45502));
    LocalMux I__8837 (
            .O(N__45510),
            .I(N__45499));
    InMux I__8836 (
            .O(N__45509),
            .I(N__45492));
    InMux I__8835 (
            .O(N__45506),
            .I(N__45492));
    InMux I__8834 (
            .O(N__45505),
            .I(N__45492));
    InMux I__8833 (
            .O(N__45502),
            .I(N__45489));
    Span4Mux_h I__8832 (
            .O(N__45499),
            .I(N__45486));
    LocalMux I__8831 (
            .O(N__45492),
            .I(N__45483));
    LocalMux I__8830 (
            .O(N__45489),
            .I(N__45480));
    Span4Mux_h I__8829 (
            .O(N__45486),
            .I(N__45476));
    Span4Mux_h I__8828 (
            .O(N__45483),
            .I(N__45473));
    Span4Mux_v I__8827 (
            .O(N__45480),
            .I(N__45470));
    CascadeMux I__8826 (
            .O(N__45479),
            .I(N__45467));
    Span4Mux_h I__8825 (
            .O(N__45476),
            .I(N__45464));
    Span4Mux_v I__8824 (
            .O(N__45473),
            .I(N__45461));
    Span4Mux_v I__8823 (
            .O(N__45470),
            .I(N__45458));
    InMux I__8822 (
            .O(N__45467),
            .I(N__45455));
    Span4Mux_v I__8821 (
            .O(N__45464),
            .I(N__45452));
    Span4Mux_h I__8820 (
            .O(N__45461),
            .I(N__45449));
    Span4Mux_h I__8819 (
            .O(N__45458),
            .I(N__45445));
    LocalMux I__8818 (
            .O(N__45455),
            .I(N__45442));
    Span4Mux_v I__8817 (
            .O(N__45452),
            .I(N__45439));
    Span4Mux_h I__8816 (
            .O(N__45449),
            .I(N__45436));
    InMux I__8815 (
            .O(N__45448),
            .I(N__45433));
    Span4Mux_v I__8814 (
            .O(N__45445),
            .I(N__45430));
    Span12Mux_v I__8813 (
            .O(N__45442),
            .I(N__45427));
    Span4Mux_v I__8812 (
            .O(N__45439),
            .I(N__45424));
    Span4Mux_v I__8811 (
            .O(N__45436),
            .I(N__45421));
    LocalMux I__8810 (
            .O(N__45433),
            .I(aluStatus_i_3));
    Odrv4 I__8809 (
            .O(N__45430),
            .I(aluStatus_i_3));
    Odrv12 I__8808 (
            .O(N__45427),
            .I(aluStatus_i_3));
    Odrv4 I__8807 (
            .O(N__45424),
            .I(aluStatus_i_3));
    Odrv4 I__8806 (
            .O(N__45421),
            .I(aluStatus_i_3));
    InMux I__8805 (
            .O(N__45410),
            .I(N__45407));
    LocalMux I__8804 (
            .O(N__45407),
            .I(N__45404));
    Span4Mux_v I__8803 (
            .O(N__45404),
            .I(N__45398));
    InMux I__8802 (
            .O(N__45403),
            .I(N__45393));
    InMux I__8801 (
            .O(N__45402),
            .I(N__45393));
    InMux I__8800 (
            .O(N__45401),
            .I(N__45387));
    Span4Mux_h I__8799 (
            .O(N__45398),
            .I(N__45382));
    LocalMux I__8798 (
            .O(N__45393),
            .I(N__45382));
    InMux I__8797 (
            .O(N__45392),
            .I(N__45375));
    InMux I__8796 (
            .O(N__45391),
            .I(N__45375));
    InMux I__8795 (
            .O(N__45390),
            .I(N__45375));
    LocalMux I__8794 (
            .O(N__45387),
            .I(PROM_ROMDATA_dintern_10ro));
    Odrv4 I__8793 (
            .O(N__45382),
            .I(PROM_ROMDATA_dintern_10ro));
    LocalMux I__8792 (
            .O(N__45375),
            .I(PROM_ROMDATA_dintern_10ro));
    CascadeMux I__8791 (
            .O(N__45368),
            .I(N__45365));
    InMux I__8790 (
            .O(N__45365),
            .I(N__45362));
    LocalMux I__8789 (
            .O(N__45362),
            .I(N__45359));
    Odrv12 I__8788 (
            .O(N__45359),
            .I(\CONTROL.g0_5Z0Z_0 ));
    InMux I__8787 (
            .O(N__45356),
            .I(N__45353));
    LocalMux I__8786 (
            .O(N__45353),
            .I(N__45350));
    Span4Mux_h I__8785 (
            .O(N__45350),
            .I(N__45347));
    Odrv4 I__8784 (
            .O(N__45347),
            .I(\PROM.ROMDATA.m258_am ));
    CascadeMux I__8783 (
            .O(N__45344),
            .I(N__45340));
    InMux I__8782 (
            .O(N__45343),
            .I(N__45335));
    InMux I__8781 (
            .O(N__45340),
            .I(N__45335));
    LocalMux I__8780 (
            .O(N__45335),
            .I(N__45332));
    Span4Mux_h I__8779 (
            .O(N__45332),
            .I(N__45329));
    Odrv4 I__8778 (
            .O(N__45329),
            .I(PROM_ROMDATA_dintern_31_0__N_555_mux));
    CascadeMux I__8777 (
            .O(N__45326),
            .I(N_417_cascade_));
    InMux I__8776 (
            .O(N__45323),
            .I(N__45320));
    LocalMux I__8775 (
            .O(N__45320),
            .I(N__45317));
    Span4Mux_v I__8774 (
            .O(N__45317),
            .I(N__45313));
    InMux I__8773 (
            .O(N__45316),
            .I(N__45310));
    Span4Mux_h I__8772 (
            .O(N__45313),
            .I(N__45305));
    LocalMux I__8771 (
            .O(N__45310),
            .I(N__45305));
    Span4Mux_h I__8770 (
            .O(N__45305),
            .I(N__45302));
    Span4Mux_v I__8769 (
            .O(N__45302),
            .I(N__45299));
    Odrv4 I__8768 (
            .O(N__45299),
            .I(\CONTROL.programCounter_1_2 ));
    InMux I__8767 (
            .O(N__45296),
            .I(N__45293));
    LocalMux I__8766 (
            .O(N__45293),
            .I(\CONTROL.programCounter_ret_1_RNI6OHFZ0Z_6 ));
    InMux I__8765 (
            .O(N__45290),
            .I(N__45287));
    LocalMux I__8764 (
            .O(N__45287),
            .I(N__45284));
    Span4Mux_v I__8763 (
            .O(N__45284),
            .I(N__45281));
    Span4Mux_h I__8762 (
            .O(N__45281),
            .I(N__45277));
    InMux I__8761 (
            .O(N__45280),
            .I(N__45274));
    Sp12to4 I__8760 (
            .O(N__45277),
            .I(N__45269));
    LocalMux I__8759 (
            .O(N__45274),
            .I(N__45269));
    Odrv12 I__8758 (
            .O(N__45269),
            .I(\CONTROL.ctrlOut_3 ));
    InMux I__8757 (
            .O(N__45266),
            .I(N__45263));
    LocalMux I__8756 (
            .O(N__45263),
            .I(N__45259));
    InMux I__8755 (
            .O(N__45262),
            .I(N__45256));
    Span4Mux_v I__8754 (
            .O(N__45259),
            .I(N__45253));
    LocalMux I__8753 (
            .O(N__45256),
            .I(N__45250));
    Span4Mux_h I__8752 (
            .O(N__45253),
            .I(N__45245));
    Span4Mux_v I__8751 (
            .O(N__45250),
            .I(N__45245));
    Odrv4 I__8750 (
            .O(N__45245),
            .I(\CONTROL.programCounter_1_4 ));
    CascadeMux I__8749 (
            .O(N__45242),
            .I(\PROM.ROMDATA.m215_ns_1_N_2L1_cascade_ ));
    InMux I__8748 (
            .O(N__45239),
            .I(N__45233));
    InMux I__8747 (
            .O(N__45238),
            .I(N__45233));
    LocalMux I__8746 (
            .O(N__45233),
            .I(N__45230));
    Span4Mux_h I__8745 (
            .O(N__45230),
            .I(N__45227));
    Span4Mux_v I__8744 (
            .O(N__45227),
            .I(N__45224));
    Odrv4 I__8743 (
            .O(N__45224),
            .I(\PROM.ROMDATA.m215_ns_1 ));
    InMux I__8742 (
            .O(N__45221),
            .I(N__45218));
    LocalMux I__8741 (
            .O(N__45218),
            .I(N__45215));
    Span4Mux_v I__8740 (
            .O(N__45215),
            .I(N__45212));
    Span4Mux_h I__8739 (
            .O(N__45212),
            .I(N__45209));
    Odrv4 I__8738 (
            .O(N__45209),
            .I(\CONTROL.g0_3_i_a7_0_0 ));
    InMux I__8737 (
            .O(N__45206),
            .I(N__45203));
    LocalMux I__8736 (
            .O(N__45203),
            .I(N__45200));
    Span12Mux_v I__8735 (
            .O(N__45200),
            .I(N__45197));
    Odrv12 I__8734 (
            .O(N__45197),
            .I(\CONTROL.addrstack_2 ));
    InMux I__8733 (
            .O(N__45194),
            .I(N__45191));
    LocalMux I__8732 (
            .O(N__45191),
            .I(\PROM.ROMDATA.m258_bm ));
    InMux I__8731 (
            .O(N__45188),
            .I(N__45184));
    InMux I__8730 (
            .O(N__45187),
            .I(N__45181));
    LocalMux I__8729 (
            .O(N__45184),
            .I(N__45178));
    LocalMux I__8728 (
            .O(N__45181),
            .I(N__45175));
    Span4Mux_h I__8727 (
            .O(N__45178),
            .I(N__45172));
    Span12Mux_h I__8726 (
            .O(N__45175),
            .I(N__45169));
    Span4Mux_v I__8725 (
            .O(N__45172),
            .I(N__45166));
    Odrv12 I__8724 (
            .O(N__45169),
            .I(\CONTROL.programCounter_1_1 ));
    Odrv4 I__8723 (
            .O(N__45166),
            .I(\CONTROL.programCounter_1_1 ));
    InMux I__8722 (
            .O(N__45161),
            .I(N__45158));
    LocalMux I__8721 (
            .O(N__45158),
            .I(\CONTROL.programCounter_ret_19_RNIT3IGZ0Z_5 ));
    InMux I__8720 (
            .O(N__45155),
            .I(N__45152));
    LocalMux I__8719 (
            .O(N__45152),
            .I(N__45149));
    Odrv4 I__8718 (
            .O(N__45149),
            .I(\CONTROL.programCounter_ret_1_RNI4MHFZ0Z_5 ));
    InMux I__8717 (
            .O(N__45146),
            .I(N__45138));
    InMux I__8716 (
            .O(N__45145),
            .I(N__45138));
    InMux I__8715 (
            .O(N__45144),
            .I(N__45133));
    InMux I__8714 (
            .O(N__45143),
            .I(N__45133));
    LocalMux I__8713 (
            .O(N__45138),
            .I(N__45130));
    LocalMux I__8712 (
            .O(N__45133),
            .I(N__45127));
    Span4Mux_v I__8711 (
            .O(N__45130),
            .I(N__45122));
    Span4Mux_h I__8710 (
            .O(N__45127),
            .I(N__45122));
    Span4Mux_h I__8709 (
            .O(N__45122),
            .I(N__45116));
    InMux I__8708 (
            .O(N__45121),
            .I(N__45113));
    InMux I__8707 (
            .O(N__45120),
            .I(N__45110));
    InMux I__8706 (
            .O(N__45119),
            .I(N__45107));
    Odrv4 I__8705 (
            .O(N__45116),
            .I(\CONTROL.un1_programCounter9_reto ));
    LocalMux I__8704 (
            .O(N__45113),
            .I(\CONTROL.un1_programCounter9_reto ));
    LocalMux I__8703 (
            .O(N__45110),
            .I(\CONTROL.un1_programCounter9_reto ));
    LocalMux I__8702 (
            .O(N__45107),
            .I(\CONTROL.un1_programCounter9_reto ));
    CascadeMux I__8701 (
            .O(N__45098),
            .I(progRomAddress_5_cascade_));
    CascadeMux I__8700 (
            .O(N__45095),
            .I(\PROM.ROMDATA.m243_1_cascade_ ));
    InMux I__8699 (
            .O(N__45092),
            .I(N__45089));
    LocalMux I__8698 (
            .O(N__45089),
            .I(N__45086));
    Span4Mux_h I__8697 (
            .O(N__45086),
            .I(N__45083));
    Odrv4 I__8696 (
            .O(N__45083),
            .I(\PROM.ROMDATA.m244_ns_1_1 ));
    InMux I__8695 (
            .O(N__45080),
            .I(N__45077));
    LocalMux I__8694 (
            .O(N__45077),
            .I(N__45073));
    InMux I__8693 (
            .O(N__45076),
            .I(N__45070));
    Odrv12 I__8692 (
            .O(N__45073),
            .I(\CONTROL.ctrlOut_0 ));
    LocalMux I__8691 (
            .O(N__45070),
            .I(\CONTROL.ctrlOut_0 ));
    InMux I__8690 (
            .O(N__45065),
            .I(N__45062));
    LocalMux I__8689 (
            .O(N__45062),
            .I(\PROM.ROMDATA.m243_1 ));
    CascadeMux I__8688 (
            .O(N__45059),
            .I(N__45055));
    CascadeMux I__8687 (
            .O(N__45058),
            .I(N__45052));
    InMux I__8686 (
            .O(N__45055),
            .I(N__45045));
    InMux I__8685 (
            .O(N__45052),
            .I(N__45045));
    InMux I__8684 (
            .O(N__45051),
            .I(N__45040));
    InMux I__8683 (
            .O(N__45050),
            .I(N__45040));
    LocalMux I__8682 (
            .O(N__45045),
            .I(N__45035));
    LocalMux I__8681 (
            .O(N__45040),
            .I(N__45035));
    Span4Mux_h I__8680 (
            .O(N__45035),
            .I(N__45032));
    Span4Mux_v I__8679 (
            .O(N__45032),
            .I(N__45028));
    InMux I__8678 (
            .O(N__45031),
            .I(N__45025));
    Odrv4 I__8677 (
            .O(N__45028),
            .I(\PROM.ROMDATA.m260_1 ));
    LocalMux I__8676 (
            .O(N__45025),
            .I(\PROM.ROMDATA.m260_1 ));
    InMux I__8675 (
            .O(N__45020),
            .I(N__45017));
    LocalMux I__8674 (
            .O(N__45017),
            .I(N__45014));
    Span4Mux_h I__8673 (
            .O(N__45014),
            .I(N__45011));
    Span4Mux_h I__8672 (
            .O(N__45011),
            .I(N__45006));
    InMux I__8671 (
            .O(N__45010),
            .I(N__45003));
    InMux I__8670 (
            .O(N__45009),
            .I(N__45000));
    Span4Mux_h I__8669 (
            .O(N__45006),
            .I(N__44995));
    LocalMux I__8668 (
            .O(N__45003),
            .I(N__44995));
    LocalMux I__8667 (
            .O(N__45000),
            .I(N__44992));
    Span4Mux_v I__8666 (
            .O(N__44995),
            .I(N__44989));
    Span4Mux_h I__8665 (
            .O(N__44992),
            .I(N__44986));
    Span4Mux_h I__8664 (
            .O(N__44989),
            .I(N__44983));
    Odrv4 I__8663 (
            .O(N__44986),
            .I(controlWord_31));
    Odrv4 I__8662 (
            .O(N__44983),
            .I(controlWord_31));
    IoInMux I__8661 (
            .O(N__44978),
            .I(N__44975));
    LocalMux I__8660 (
            .O(N__44975),
            .I(N__44972));
    IoSpan4Mux I__8659 (
            .O(N__44972),
            .I(N__44969));
    Span4Mux_s1_v I__8658 (
            .O(N__44969),
            .I(N__44966));
    Sp12to4 I__8657 (
            .O(N__44966),
            .I(N__44963));
    Span12Mux_h I__8656 (
            .O(N__44963),
            .I(N__44959));
    CascadeMux I__8655 (
            .O(N__44962),
            .I(N__44956));
    Span12Mux_v I__8654 (
            .O(N__44959),
            .I(N__44953));
    InMux I__8653 (
            .O(N__44956),
            .I(N__44950));
    Odrv12 I__8652 (
            .O(N__44953),
            .I(A15_c));
    LocalMux I__8651 (
            .O(N__44950),
            .I(A15_c));
    InMux I__8650 (
            .O(N__44945),
            .I(N__44942));
    LocalMux I__8649 (
            .O(N__44942),
            .I(\PROM.ROMDATA.m266 ));
    CascadeMux I__8648 (
            .O(N__44939),
            .I(\PROM.ROMDATA.m157_cascade_ ));
    CascadeMux I__8647 (
            .O(N__44936),
            .I(\PROM.ROMDATA.m265_cascade_ ));
    InMux I__8646 (
            .O(N__44933),
            .I(N__44930));
    LocalMux I__8645 (
            .O(N__44930),
            .I(\PROM.ROMDATA.m268 ));
    InMux I__8644 (
            .O(N__44927),
            .I(N__44924));
    LocalMux I__8643 (
            .O(N__44924),
            .I(N__44921));
    Span4Mux_h I__8642 (
            .O(N__44921),
            .I(N__44917));
    InMux I__8641 (
            .O(N__44920),
            .I(N__44914));
    Odrv4 I__8640 (
            .O(N__44917),
            .I(\PROM.ROMDATA.m270_bm ));
    LocalMux I__8639 (
            .O(N__44914),
            .I(\PROM.ROMDATA.m270_bm ));
    InMux I__8638 (
            .O(N__44909),
            .I(N__44906));
    LocalMux I__8637 (
            .O(N__44906),
            .I(\CONTROL.aluOperation_12_i_0_6 ));
    InMux I__8636 (
            .O(N__44903),
            .I(N__44891));
    InMux I__8635 (
            .O(N__44902),
            .I(N__44891));
    InMux I__8634 (
            .O(N__44901),
            .I(N__44888));
    InMux I__8633 (
            .O(N__44900),
            .I(N__44885));
    InMux I__8632 (
            .O(N__44899),
            .I(N__44879));
    InMux I__8631 (
            .O(N__44898),
            .I(N__44872));
    InMux I__8630 (
            .O(N__44897),
            .I(N__44872));
    InMux I__8629 (
            .O(N__44896),
            .I(N__44872));
    LocalMux I__8628 (
            .O(N__44891),
            .I(N__44859));
    LocalMux I__8627 (
            .O(N__44888),
            .I(N__44854));
    LocalMux I__8626 (
            .O(N__44885),
            .I(N__44854));
    InMux I__8625 (
            .O(N__44884),
            .I(N__44849));
    InMux I__8624 (
            .O(N__44883),
            .I(N__44849));
    InMux I__8623 (
            .O(N__44882),
            .I(N__44846));
    LocalMux I__8622 (
            .O(N__44879),
            .I(N__44841));
    LocalMux I__8621 (
            .O(N__44872),
            .I(N__44841));
    InMux I__8620 (
            .O(N__44871),
            .I(N__44836));
    InMux I__8619 (
            .O(N__44870),
            .I(N__44827));
    InMux I__8618 (
            .O(N__44869),
            .I(N__44827));
    InMux I__8617 (
            .O(N__44868),
            .I(N__44827));
    InMux I__8616 (
            .O(N__44867),
            .I(N__44827));
    InMux I__8615 (
            .O(N__44866),
            .I(N__44824));
    InMux I__8614 (
            .O(N__44865),
            .I(N__44819));
    InMux I__8613 (
            .O(N__44864),
            .I(N__44819));
    InMux I__8612 (
            .O(N__44863),
            .I(N__44816));
    InMux I__8611 (
            .O(N__44862),
            .I(N__44813));
    Span4Mux_h I__8610 (
            .O(N__44859),
            .I(N__44810));
    Span4Mux_h I__8609 (
            .O(N__44854),
            .I(N__44801));
    LocalMux I__8608 (
            .O(N__44849),
            .I(N__44801));
    LocalMux I__8607 (
            .O(N__44846),
            .I(N__44801));
    Span4Mux_h I__8606 (
            .O(N__44841),
            .I(N__44801));
    InMux I__8605 (
            .O(N__44840),
            .I(N__44796));
    InMux I__8604 (
            .O(N__44839),
            .I(N__44796));
    LocalMux I__8603 (
            .O(N__44836),
            .I(N__44791));
    LocalMux I__8602 (
            .O(N__44827),
            .I(N__44791));
    LocalMux I__8601 (
            .O(N__44824),
            .I(controlWord_3));
    LocalMux I__8600 (
            .O(N__44819),
            .I(controlWord_3));
    LocalMux I__8599 (
            .O(N__44816),
            .I(controlWord_3));
    LocalMux I__8598 (
            .O(N__44813),
            .I(controlWord_3));
    Odrv4 I__8597 (
            .O(N__44810),
            .I(controlWord_3));
    Odrv4 I__8596 (
            .O(N__44801),
            .I(controlWord_3));
    LocalMux I__8595 (
            .O(N__44796),
            .I(controlWord_3));
    Odrv4 I__8594 (
            .O(N__44791),
            .I(controlWord_3));
    CascadeMux I__8593 (
            .O(N__44774),
            .I(N__44770));
    CascadeMux I__8592 (
            .O(N__44773),
            .I(N__44766));
    InMux I__8591 (
            .O(N__44770),
            .I(N__44763));
    InMux I__8590 (
            .O(N__44769),
            .I(N__44760));
    InMux I__8589 (
            .O(N__44766),
            .I(N__44756));
    LocalMux I__8588 (
            .O(N__44763),
            .I(N__44753));
    LocalMux I__8587 (
            .O(N__44760),
            .I(N__44750));
    CascadeMux I__8586 (
            .O(N__44759),
            .I(N__44745));
    LocalMux I__8585 (
            .O(N__44756),
            .I(N__44742));
    Span4Mux_h I__8584 (
            .O(N__44753),
            .I(N__44739));
    Span4Mux_h I__8583 (
            .O(N__44750),
            .I(N__44736));
    InMux I__8582 (
            .O(N__44749),
            .I(N__44731));
    InMux I__8581 (
            .O(N__44748),
            .I(N__44731));
    InMux I__8580 (
            .O(N__44745),
            .I(N__44728));
    Span4Mux_h I__8579 (
            .O(N__44742),
            .I(N__44725));
    Odrv4 I__8578 (
            .O(N__44739),
            .I(\CONTROL.N_219 ));
    Odrv4 I__8577 (
            .O(N__44736),
            .I(\CONTROL.N_219 ));
    LocalMux I__8576 (
            .O(N__44731),
            .I(\CONTROL.N_219 ));
    LocalMux I__8575 (
            .O(N__44728),
            .I(\CONTROL.N_219 ));
    Odrv4 I__8574 (
            .O(N__44725),
            .I(\CONTROL.N_219 ));
    InMux I__8573 (
            .O(N__44714),
            .I(N__44709));
    CascadeMux I__8572 (
            .O(N__44713),
            .I(N__44697));
    InMux I__8571 (
            .O(N__44712),
            .I(N__44693));
    LocalMux I__8570 (
            .O(N__44709),
            .I(N__44690));
    InMux I__8569 (
            .O(N__44708),
            .I(N__44687));
    InMux I__8568 (
            .O(N__44707),
            .I(N__44680));
    InMux I__8567 (
            .O(N__44706),
            .I(N__44680));
    InMux I__8566 (
            .O(N__44705),
            .I(N__44680));
    InMux I__8565 (
            .O(N__44704),
            .I(N__44676));
    InMux I__8564 (
            .O(N__44703),
            .I(N__44673));
    InMux I__8563 (
            .O(N__44702),
            .I(N__44670));
    InMux I__8562 (
            .O(N__44701),
            .I(N__44667));
    InMux I__8561 (
            .O(N__44700),
            .I(N__44664));
    InMux I__8560 (
            .O(N__44697),
            .I(N__44651));
    InMux I__8559 (
            .O(N__44696),
            .I(N__44646));
    LocalMux I__8558 (
            .O(N__44693),
            .I(N__44641));
    Span4Mux_v I__8557 (
            .O(N__44690),
            .I(N__44641));
    LocalMux I__8556 (
            .O(N__44687),
            .I(N__44626));
    LocalMux I__8555 (
            .O(N__44680),
            .I(N__44626));
    InMux I__8554 (
            .O(N__44679),
            .I(N__44623));
    LocalMux I__8553 (
            .O(N__44676),
            .I(N__44620));
    LocalMux I__8552 (
            .O(N__44673),
            .I(N__44615));
    LocalMux I__8551 (
            .O(N__44670),
            .I(N__44615));
    LocalMux I__8550 (
            .O(N__44667),
            .I(N__44612));
    LocalMux I__8549 (
            .O(N__44664),
            .I(N__44609));
    InMux I__8548 (
            .O(N__44663),
            .I(N__44604));
    InMux I__8547 (
            .O(N__44662),
            .I(N__44604));
    InMux I__8546 (
            .O(N__44661),
            .I(N__44601));
    InMux I__8545 (
            .O(N__44660),
            .I(N__44594));
    InMux I__8544 (
            .O(N__44659),
            .I(N__44594));
    InMux I__8543 (
            .O(N__44658),
            .I(N__44594));
    InMux I__8542 (
            .O(N__44657),
            .I(N__44585));
    InMux I__8541 (
            .O(N__44656),
            .I(N__44585));
    InMux I__8540 (
            .O(N__44655),
            .I(N__44585));
    InMux I__8539 (
            .O(N__44654),
            .I(N__44585));
    LocalMux I__8538 (
            .O(N__44651),
            .I(N__44582));
    InMux I__8537 (
            .O(N__44650),
            .I(N__44579));
    InMux I__8536 (
            .O(N__44649),
            .I(N__44576));
    LocalMux I__8535 (
            .O(N__44646),
            .I(N__44573));
    Span4Mux_h I__8534 (
            .O(N__44641),
            .I(N__44570));
    InMux I__8533 (
            .O(N__44640),
            .I(N__44565));
    InMux I__8532 (
            .O(N__44639),
            .I(N__44565));
    InMux I__8531 (
            .O(N__44638),
            .I(N__44560));
    InMux I__8530 (
            .O(N__44637),
            .I(N__44560));
    InMux I__8529 (
            .O(N__44636),
            .I(N__44549));
    InMux I__8528 (
            .O(N__44635),
            .I(N__44549));
    InMux I__8527 (
            .O(N__44634),
            .I(N__44549));
    InMux I__8526 (
            .O(N__44633),
            .I(N__44549));
    InMux I__8525 (
            .O(N__44632),
            .I(N__44549));
    InMux I__8524 (
            .O(N__44631),
            .I(N__44546));
    Span4Mux_v I__8523 (
            .O(N__44626),
            .I(N__44541));
    LocalMux I__8522 (
            .O(N__44623),
            .I(N__44541));
    Span4Mux_v I__8521 (
            .O(N__44620),
            .I(N__44530));
    Span4Mux_v I__8520 (
            .O(N__44615),
            .I(N__44530));
    Span4Mux_h I__8519 (
            .O(N__44612),
            .I(N__44530));
    Span4Mux_v I__8518 (
            .O(N__44609),
            .I(N__44530));
    LocalMux I__8517 (
            .O(N__44604),
            .I(N__44530));
    LocalMux I__8516 (
            .O(N__44601),
            .I(N__44523));
    LocalMux I__8515 (
            .O(N__44594),
            .I(N__44523));
    LocalMux I__8514 (
            .O(N__44585),
            .I(N__44523));
    Odrv4 I__8513 (
            .O(N__44582),
            .I(controlWord_2));
    LocalMux I__8512 (
            .O(N__44579),
            .I(controlWord_2));
    LocalMux I__8511 (
            .O(N__44576),
            .I(controlWord_2));
    Odrv12 I__8510 (
            .O(N__44573),
            .I(controlWord_2));
    Odrv4 I__8509 (
            .O(N__44570),
            .I(controlWord_2));
    LocalMux I__8508 (
            .O(N__44565),
            .I(controlWord_2));
    LocalMux I__8507 (
            .O(N__44560),
            .I(controlWord_2));
    LocalMux I__8506 (
            .O(N__44549),
            .I(controlWord_2));
    LocalMux I__8505 (
            .O(N__44546),
            .I(controlWord_2));
    Odrv4 I__8504 (
            .O(N__44541),
            .I(controlWord_2));
    Odrv4 I__8503 (
            .O(N__44530),
            .I(controlWord_2));
    Odrv4 I__8502 (
            .O(N__44523),
            .I(controlWord_2));
    InMux I__8501 (
            .O(N__44498),
            .I(N__44490));
    InMux I__8500 (
            .O(N__44497),
            .I(N__44490));
    InMux I__8499 (
            .O(N__44496),
            .I(N__44485));
    InMux I__8498 (
            .O(N__44495),
            .I(N__44485));
    LocalMux I__8497 (
            .O(N__44490),
            .I(N__44482));
    LocalMux I__8496 (
            .O(N__44485),
            .I(N__44479));
    Span12Mux_v I__8495 (
            .O(N__44482),
            .I(N__44475));
    Span4Mux_v I__8494 (
            .O(N__44479),
            .I(N__44472));
    InMux I__8493 (
            .O(N__44478),
            .I(N__44469));
    Odrv12 I__8492 (
            .O(N__44475),
            .I(\PROM.ROMDATA.N_544_mux ));
    Odrv4 I__8491 (
            .O(N__44472),
            .I(\PROM.ROMDATA.N_544_mux ));
    LocalMux I__8490 (
            .O(N__44469),
            .I(\PROM.ROMDATA.N_544_mux ));
    CEMux I__8489 (
            .O(N__44462),
            .I(N__44458));
    CEMux I__8488 (
            .O(N__44461),
            .I(N__44454));
    LocalMux I__8487 (
            .O(N__44458),
            .I(N__44449));
    CEMux I__8486 (
            .O(N__44457),
            .I(N__44446));
    LocalMux I__8485 (
            .O(N__44454),
            .I(N__44442));
    CEMux I__8484 (
            .O(N__44453),
            .I(N__44439));
    CEMux I__8483 (
            .O(N__44452),
            .I(N__44436));
    Span4Mux_h I__8482 (
            .O(N__44449),
            .I(N__44429));
    LocalMux I__8481 (
            .O(N__44446),
            .I(N__44429));
    CEMux I__8480 (
            .O(N__44445),
            .I(N__44426));
    Span4Mux_h I__8479 (
            .O(N__44442),
            .I(N__44419));
    LocalMux I__8478 (
            .O(N__44439),
            .I(N__44419));
    LocalMux I__8477 (
            .O(N__44436),
            .I(N__44419));
    CEMux I__8476 (
            .O(N__44435),
            .I(N__44416));
    CEMux I__8475 (
            .O(N__44434),
            .I(N__44412));
    Span4Mux_h I__8474 (
            .O(N__44429),
            .I(N__44407));
    LocalMux I__8473 (
            .O(N__44426),
            .I(N__44407));
    Span4Mux_v I__8472 (
            .O(N__44419),
            .I(N__44402));
    LocalMux I__8471 (
            .O(N__44416),
            .I(N__44402));
    CEMux I__8470 (
            .O(N__44415),
            .I(N__44399));
    LocalMux I__8469 (
            .O(N__44412),
            .I(N__44393));
    Span4Mux_v I__8468 (
            .O(N__44407),
            .I(N__44390));
    Span4Mux_v I__8467 (
            .O(N__44402),
            .I(N__44385));
    LocalMux I__8466 (
            .O(N__44399),
            .I(N__44385));
    CEMux I__8465 (
            .O(N__44398),
            .I(N__44382));
    CEMux I__8464 (
            .O(N__44397),
            .I(N__44379));
    CEMux I__8463 (
            .O(N__44396),
            .I(N__44376));
    Span4Mux_h I__8462 (
            .O(N__44393),
            .I(N__44373));
    Span4Mux_h I__8461 (
            .O(N__44390),
            .I(N__44370));
    Span4Mux_h I__8460 (
            .O(N__44385),
            .I(N__44365));
    LocalMux I__8459 (
            .O(N__44382),
            .I(N__44365));
    LocalMux I__8458 (
            .O(N__44379),
            .I(N__44362));
    LocalMux I__8457 (
            .O(N__44376),
            .I(N__44359));
    Span4Mux_h I__8456 (
            .O(N__44373),
            .I(N__44356));
    Span4Mux_h I__8455 (
            .O(N__44370),
            .I(N__44353));
    Span4Mux_h I__8454 (
            .O(N__44365),
            .I(N__44350));
    Span4Mux_v I__8453 (
            .O(N__44362),
            .I(N__44345));
    Span4Mux_v I__8452 (
            .O(N__44359),
            .I(N__44345));
    Odrv4 I__8451 (
            .O(N__44356),
            .I(\CONTROL.N_35 ));
    Odrv4 I__8450 (
            .O(N__44353),
            .I(\CONTROL.N_35 ));
    Odrv4 I__8449 (
            .O(N__44350),
            .I(\CONTROL.N_35 ));
    Odrv4 I__8448 (
            .O(N__44345),
            .I(\CONTROL.N_35 ));
    InMux I__8447 (
            .O(N__44336),
            .I(N__44333));
    LocalMux I__8446 (
            .O(N__44333),
            .I(N__44330));
    Odrv4 I__8445 (
            .O(N__44330),
            .I(\PROM.ROMDATA.m444_am ));
    CascadeMux I__8444 (
            .O(N__44327),
            .I(\PROM.ROMDATA.m444_bm_cascade_ ));
    CascadeMux I__8443 (
            .O(N__44324),
            .I(N__44321));
    InMux I__8442 (
            .O(N__44321),
            .I(N__44315));
    InMux I__8441 (
            .O(N__44320),
            .I(N__44315));
    LocalMux I__8440 (
            .O(N__44315),
            .I(N__44312));
    Span4Mux_h I__8439 (
            .O(N__44312),
            .I(N__44309));
    Span4Mux_h I__8438 (
            .O(N__44309),
            .I(N__44304));
    InMux I__8437 (
            .O(N__44308),
            .I(N__44299));
    InMux I__8436 (
            .O(N__44307),
            .I(N__44299));
    Odrv4 I__8435 (
            .O(N__44304),
            .I(\PROM.ROMDATA.m289 ));
    LocalMux I__8434 (
            .O(N__44299),
            .I(\PROM.ROMDATA.m289 ));
    CascadeMux I__8433 (
            .O(N__44294),
            .I(N__44291));
    InMux I__8432 (
            .O(N__44291),
            .I(N__44288));
    LocalMux I__8431 (
            .O(N__44288),
            .I(N__44285));
    Span4Mux_v I__8430 (
            .O(N__44285),
            .I(N__44282));
    Odrv4 I__8429 (
            .O(N__44282),
            .I(\PROM.ROMDATA.m418_ns_1 ));
    InMux I__8428 (
            .O(N__44279),
            .I(N__44273));
    InMux I__8427 (
            .O(N__44278),
            .I(N__44273));
    LocalMux I__8426 (
            .O(N__44273),
            .I(N__44270));
    Span4Mux_h I__8425 (
            .O(N__44270),
            .I(N__44267));
    Span4Mux_h I__8424 (
            .O(N__44267),
            .I(N__44264));
    Span4Mux_h I__8423 (
            .O(N__44264),
            .I(N__44261));
    Odrv4 I__8422 (
            .O(N__44261),
            .I(PROM_ROMDATA_dintern_19ro));
    CascadeMux I__8421 (
            .O(N__44258),
            .I(PROM_ROMDATA_dintern_19ro_cascade_));
    InMux I__8420 (
            .O(N__44255),
            .I(N__44252));
    LocalMux I__8419 (
            .O(N__44252),
            .I(N__44249));
    Span12Mux_h I__8418 (
            .O(N__44249),
            .I(N__44246));
    Odrv12 I__8417 (
            .O(N__44246),
            .I(controlWord_19));
    InMux I__8416 (
            .O(N__44243),
            .I(N__44239));
    CascadeMux I__8415 (
            .O(N__44242),
            .I(N__44236));
    LocalMux I__8414 (
            .O(N__44239),
            .I(N__44232));
    InMux I__8413 (
            .O(N__44236),
            .I(N__44229));
    CascadeMux I__8412 (
            .O(N__44235),
            .I(N__44226));
    Span4Mux_v I__8411 (
            .O(N__44232),
            .I(N__44223));
    LocalMux I__8410 (
            .O(N__44229),
            .I(N__44220));
    InMux I__8409 (
            .O(N__44226),
            .I(N__44217));
    Span4Mux_h I__8408 (
            .O(N__44223),
            .I(N__44212));
    Span4Mux_v I__8407 (
            .O(N__44220),
            .I(N__44212));
    LocalMux I__8406 (
            .O(N__44217),
            .I(N__44209));
    Span4Mux_v I__8405 (
            .O(N__44212),
            .I(N__44206));
    Span4Mux_v I__8404 (
            .O(N__44209),
            .I(N__44203));
    Sp12to4 I__8403 (
            .O(N__44206),
            .I(N__44200));
    Odrv4 I__8402 (
            .O(N__44203),
            .I(f_3));
    Odrv12 I__8401 (
            .O(N__44200),
            .I(f_3));
    CascadeMux I__8400 (
            .O(N__44195),
            .I(controlWord_19_cascade_));
    InMux I__8399 (
            .O(N__44192),
            .I(N__44189));
    LocalMux I__8398 (
            .O(N__44189),
            .I(N__44185));
    InMux I__8397 (
            .O(N__44188),
            .I(N__44182));
    Span4Mux_h I__8396 (
            .O(N__44185),
            .I(N__44179));
    LocalMux I__8395 (
            .O(N__44182),
            .I(N__44173));
    Span4Mux_h I__8394 (
            .O(N__44179),
            .I(N__44173));
    InMux I__8393 (
            .O(N__44178),
            .I(N__44170));
    Span4Mux_h I__8392 (
            .O(N__44173),
            .I(N__44167));
    LocalMux I__8391 (
            .O(N__44170),
            .I(controlWord_20));
    Odrv4 I__8390 (
            .O(N__44167),
            .I(controlWord_20));
    CascadeMux I__8389 (
            .O(N__44162),
            .I(N__44159));
    InMux I__8388 (
            .O(N__44159),
            .I(N__44156));
    LocalMux I__8387 (
            .O(N__44156),
            .I(N__44152));
    CascadeMux I__8386 (
            .O(N__44155),
            .I(N__44149));
    Span4Mux_h I__8385 (
            .O(N__44152),
            .I(N__44146));
    InMux I__8384 (
            .O(N__44149),
            .I(N__44143));
    Span4Mux_h I__8383 (
            .O(N__44146),
            .I(N__44140));
    LocalMux I__8382 (
            .O(N__44143),
            .I(N__44136));
    Span4Mux_v I__8381 (
            .O(N__44140),
            .I(N__44133));
    InMux I__8380 (
            .O(N__44139),
            .I(N__44130));
    Span4Mux_h I__8379 (
            .O(N__44136),
            .I(N__44127));
    Span4Mux_h I__8378 (
            .O(N__44133),
            .I(N__44122));
    LocalMux I__8377 (
            .O(N__44130),
            .I(N__44122));
    Span4Mux_h I__8376 (
            .O(N__44127),
            .I(N__44119));
    Span4Mux_h I__8375 (
            .O(N__44122),
            .I(N__44116));
    Odrv4 I__8374 (
            .O(N__44119),
            .I(f_4));
    Odrv4 I__8373 (
            .O(N__44116),
            .I(f_4));
    IoInMux I__8372 (
            .O(N__44111),
            .I(N__44108));
    LocalMux I__8371 (
            .O(N__44108),
            .I(N__44105));
    Span4Mux_s2_v I__8370 (
            .O(N__44105),
            .I(N__44102));
    Span4Mux_h I__8369 (
            .O(N__44102),
            .I(N__44098));
    InMux I__8368 (
            .O(N__44101),
            .I(N__44095));
    Span4Mux_h I__8367 (
            .O(N__44098),
            .I(N__44092));
    LocalMux I__8366 (
            .O(N__44095),
            .I(N__44089));
    Span4Mux_h I__8365 (
            .O(N__44092),
            .I(N__44086));
    Span4Mux_v I__8364 (
            .O(N__44089),
            .I(N__44083));
    Span4Mux_v I__8363 (
            .O(N__44086),
            .I(N__44078));
    Span4Mux_v I__8362 (
            .O(N__44083),
            .I(N__44078));
    Span4Mux_h I__8361 (
            .O(N__44078),
            .I(N__44075));
    Odrv4 I__8360 (
            .O(N__44075),
            .I(A14_c));
    IoInMux I__8359 (
            .O(N__44072),
            .I(N__44069));
    LocalMux I__8358 (
            .O(N__44069),
            .I(N__44066));
    Span4Mux_s2_h I__8357 (
            .O(N__44066),
            .I(N__44063));
    Span4Mux_v I__8356 (
            .O(N__44063),
            .I(N__44060));
    Sp12to4 I__8355 (
            .O(N__44060),
            .I(N__44056));
    InMux I__8354 (
            .O(N__44059),
            .I(N__44053));
    Odrv12 I__8353 (
            .O(N__44056),
            .I(A4_c));
    LocalMux I__8352 (
            .O(N__44053),
            .I(A4_c));
    IoInMux I__8351 (
            .O(N__44048),
            .I(N__44045));
    LocalMux I__8350 (
            .O(N__44045),
            .I(N__44042));
    Span4Mux_s1_h I__8349 (
            .O(N__44042),
            .I(N__44039));
    Sp12to4 I__8348 (
            .O(N__44039),
            .I(N__44036));
    Span12Mux_v I__8347 (
            .O(N__44036),
            .I(N__44033));
    Span12Mux_h I__8346 (
            .O(N__44033),
            .I(N__44029));
    InMux I__8345 (
            .O(N__44032),
            .I(N__44026));
    Odrv12 I__8344 (
            .O(N__44029),
            .I(A3_c));
    LocalMux I__8343 (
            .O(N__44026),
            .I(A3_c));
    InMux I__8342 (
            .O(N__44021),
            .I(N__44018));
    LocalMux I__8341 (
            .O(N__44018),
            .I(N__44015));
    Span4Mux_h I__8340 (
            .O(N__44015),
            .I(N__44012));
    Span4Mux_v I__8339 (
            .O(N__44012),
            .I(N__44009));
    Sp12to4 I__8338 (
            .O(N__44009),
            .I(N__44006));
    Span12Mux_h I__8337 (
            .O(N__44006),
            .I(N__44003));
    Odrv12 I__8336 (
            .O(N__44003),
            .I(\RAM.un1_WR_105_0Z0Z_7 ));
    InMux I__8335 (
            .O(N__44000),
            .I(N__43992));
    InMux I__8334 (
            .O(N__43999),
            .I(N__43992));
    InMux I__8333 (
            .O(N__43998),
            .I(N__43987));
    InMux I__8332 (
            .O(N__43997),
            .I(N__43987));
    LocalMux I__8331 (
            .O(N__43992),
            .I(N__43984));
    LocalMux I__8330 (
            .O(N__43987),
            .I(N__43976));
    Span4Mux_h I__8329 (
            .O(N__43984),
            .I(N__43971));
    InMux I__8328 (
            .O(N__43983),
            .I(N__43964));
    InMux I__8327 (
            .O(N__43982),
            .I(N__43964));
    InMux I__8326 (
            .O(N__43981),
            .I(N__43964));
    InMux I__8325 (
            .O(N__43980),
            .I(N__43959));
    InMux I__8324 (
            .O(N__43979),
            .I(N__43959));
    Span4Mux_h I__8323 (
            .O(N__43976),
            .I(N__43956));
    InMux I__8322 (
            .O(N__43975),
            .I(N__43951));
    InMux I__8321 (
            .O(N__43974),
            .I(N__43951));
    Span4Mux_h I__8320 (
            .O(N__43971),
            .I(N__43948));
    LocalMux I__8319 (
            .O(N__43964),
            .I(aluOperand2_2_rep1));
    LocalMux I__8318 (
            .O(N__43959),
            .I(aluOperand2_2_rep1));
    Odrv4 I__8317 (
            .O(N__43956),
            .I(aluOperand2_2_rep1));
    LocalMux I__8316 (
            .O(N__43951),
            .I(aluOperand2_2_rep1));
    Odrv4 I__8315 (
            .O(N__43948),
            .I(aluOperand2_2_rep1));
    InMux I__8314 (
            .O(N__43937),
            .I(N__43934));
    LocalMux I__8313 (
            .O(N__43934),
            .I(\ALU.operand2_3_ns_1_7 ));
    InMux I__8312 (
            .O(N__43931),
            .I(N__43925));
    InMux I__8311 (
            .O(N__43930),
            .I(N__43925));
    LocalMux I__8310 (
            .O(N__43925),
            .I(N__43922));
    Span4Mux_h I__8309 (
            .O(N__43922),
            .I(N__43909));
    InMux I__8308 (
            .O(N__43921),
            .I(N__43904));
    InMux I__8307 (
            .O(N__43920),
            .I(N__43904));
    InMux I__8306 (
            .O(N__43919),
            .I(N__43898));
    InMux I__8305 (
            .O(N__43918),
            .I(N__43898));
    InMux I__8304 (
            .O(N__43917),
            .I(N__43891));
    InMux I__8303 (
            .O(N__43916),
            .I(N__43891));
    InMux I__8302 (
            .O(N__43915),
            .I(N__43886));
    InMux I__8301 (
            .O(N__43914),
            .I(N__43886));
    InMux I__8300 (
            .O(N__43913),
            .I(N__43881));
    InMux I__8299 (
            .O(N__43912),
            .I(N__43881));
    Span4Mux_h I__8298 (
            .O(N__43909),
            .I(N__43878));
    LocalMux I__8297 (
            .O(N__43904),
            .I(N__43875));
    InMux I__8296 (
            .O(N__43903),
            .I(N__43872));
    LocalMux I__8295 (
            .O(N__43898),
            .I(N__43869));
    InMux I__8294 (
            .O(N__43897),
            .I(N__43866));
    InMux I__8293 (
            .O(N__43896),
            .I(N__43863));
    LocalMux I__8292 (
            .O(N__43891),
            .I(N__43858));
    LocalMux I__8291 (
            .O(N__43886),
            .I(N__43858));
    LocalMux I__8290 (
            .O(N__43881),
            .I(N__43853));
    Span4Mux_v I__8289 (
            .O(N__43878),
            .I(N__43853));
    Span4Mux_v I__8288 (
            .O(N__43875),
            .I(N__43850));
    LocalMux I__8287 (
            .O(N__43872),
            .I(aluOperand1_1_rep1));
    Odrv4 I__8286 (
            .O(N__43869),
            .I(aluOperand1_1_rep1));
    LocalMux I__8285 (
            .O(N__43866),
            .I(aluOperand1_1_rep1));
    LocalMux I__8284 (
            .O(N__43863),
            .I(aluOperand1_1_rep1));
    Odrv12 I__8283 (
            .O(N__43858),
            .I(aluOperand1_1_rep1));
    Odrv4 I__8282 (
            .O(N__43853),
            .I(aluOperand1_1_rep1));
    Odrv4 I__8281 (
            .O(N__43850),
            .I(aluOperand1_1_rep1));
    InMux I__8280 (
            .O(N__43835),
            .I(N__43832));
    LocalMux I__8279 (
            .O(N__43832),
            .I(N__43829));
    Span4Mux_v I__8278 (
            .O(N__43829),
            .I(N__43826));
    Span4Mux_v I__8277 (
            .O(N__43826),
            .I(N__43823));
    Sp12to4 I__8276 (
            .O(N__43823),
            .I(N__43819));
    CascadeMux I__8275 (
            .O(N__43822),
            .I(N__43816));
    Span12Mux_h I__8274 (
            .O(N__43819),
            .I(N__43812));
    InMux I__8273 (
            .O(N__43816),
            .I(N__43809));
    InMux I__8272 (
            .O(N__43815),
            .I(N__43806));
    Odrv12 I__8271 (
            .O(N__43812),
            .I(h_7));
    LocalMux I__8270 (
            .O(N__43809),
            .I(h_7));
    LocalMux I__8269 (
            .O(N__43806),
            .I(h_7));
    CascadeMux I__8268 (
            .O(N__43799),
            .I(\ALU.dout_6_ns_1_7_cascade_ ));
    CascadeMux I__8267 (
            .O(N__43796),
            .I(\ALU.N_1140_cascade_ ));
    InMux I__8266 (
            .O(N__43793),
            .I(N__43790));
    LocalMux I__8265 (
            .O(N__43790),
            .I(\ALU.N_1092 ));
    InMux I__8264 (
            .O(N__43787),
            .I(N__43784));
    LocalMux I__8263 (
            .O(N__43784),
            .I(N__43781));
    Span4Mux_h I__8262 (
            .O(N__43781),
            .I(N__43778));
    Span4Mux_h I__8261 (
            .O(N__43778),
            .I(N__43775));
    Odrv4 I__8260 (
            .O(N__43775),
            .I(DROM_ROMDATA_dintern_7ro));
    CascadeMux I__8259 (
            .O(N__43772),
            .I(aluOut_7_cascade_));
    InMux I__8258 (
            .O(N__43769),
            .I(N__43766));
    LocalMux I__8257 (
            .O(N__43766),
            .I(N__43763));
    Span4Mux_h I__8256 (
            .O(N__43763),
            .I(N__43760));
    Span4Mux_h I__8255 (
            .O(N__43760),
            .I(N__43756));
    InMux I__8254 (
            .O(N__43759),
            .I(N__43753));
    Odrv4 I__8253 (
            .O(N__43756),
            .I(N_200));
    LocalMux I__8252 (
            .O(N__43753),
            .I(N_200));
    CascadeMux I__8251 (
            .O(N__43748),
            .I(\PROM.ROMDATA.m267_cascade_ ));
    CascadeMux I__8250 (
            .O(N__43745),
            .I(N__43741));
    InMux I__8249 (
            .O(N__43744),
            .I(N__43736));
    InMux I__8248 (
            .O(N__43741),
            .I(N__43736));
    LocalMux I__8247 (
            .O(N__43736),
            .I(N__43733));
    Span4Mux_v I__8246 (
            .O(N__43733),
            .I(N__43730));
    Sp12to4 I__8245 (
            .O(N__43730),
            .I(N__43727));
    Span12Mux_h I__8244 (
            .O(N__43727),
            .I(N__43724));
    Odrv12 I__8243 (
            .O(N__43724),
            .I(\PROM.ROMDATA.m442 ));
    InMux I__8242 (
            .O(N__43721),
            .I(N__43718));
    LocalMux I__8241 (
            .O(N__43718),
            .I(N__43715));
    Span12Mux_h I__8240 (
            .O(N__43715),
            .I(N__43711));
    InMux I__8239 (
            .O(N__43714),
            .I(N__43708));
    Odrv12 I__8238 (
            .O(N__43711),
            .I(\PROM.ROMDATA.m282 ));
    LocalMux I__8237 (
            .O(N__43708),
            .I(\PROM.ROMDATA.m282 ));
    InMux I__8236 (
            .O(N__43703),
            .I(N__43700));
    LocalMux I__8235 (
            .O(N__43700),
            .I(N__43697));
    Span4Mux_h I__8234 (
            .O(N__43697),
            .I(N__43694));
    Span4Mux_h I__8233 (
            .O(N__43694),
            .I(N__43691));
    Span4Mux_h I__8232 (
            .O(N__43691),
            .I(N__43687));
    InMux I__8231 (
            .O(N__43690),
            .I(N__43684));
    Odrv4 I__8230 (
            .O(N__43687),
            .I(\PROM.ROMDATA.dintern_29dfltZ0Z_1 ));
    LocalMux I__8229 (
            .O(N__43684),
            .I(\PROM.ROMDATA.dintern_29dfltZ0Z_1 ));
    CascadeMux I__8228 (
            .O(N__43679),
            .I(\PROM.ROMDATA.m282_cascade_ ));
    InMux I__8227 (
            .O(N__43676),
            .I(N__43673));
    LocalMux I__8226 (
            .O(N__43673),
            .I(N__43670));
    Span4Mux_v I__8225 (
            .O(N__43670),
            .I(N__43666));
    InMux I__8224 (
            .O(N__43669),
            .I(N__43663));
    Span4Mux_h I__8223 (
            .O(N__43666),
            .I(N__43658));
    LocalMux I__8222 (
            .O(N__43663),
            .I(N__43658));
    Span4Mux_v I__8221 (
            .O(N__43658),
            .I(N__43655));
    Span4Mux_h I__8220 (
            .O(N__43655),
            .I(N__43652));
    Odrv4 I__8219 (
            .O(N__43652),
            .I(\CONTROL.ctrlOut_13 ));
    CascadeMux I__8218 (
            .O(N__43649),
            .I(\ALU.N_1252_cascade_ ));
    InMux I__8217 (
            .O(N__43646),
            .I(N__43643));
    LocalMux I__8216 (
            .O(N__43643),
            .I(\ALU.N_1204 ));
    CascadeMux I__8215 (
            .O(N__43640),
            .I(\ALU.d_RNIO5IF4Z0Z_7_cascade_ ));
    InMux I__8214 (
            .O(N__43637),
            .I(N__43634));
    LocalMux I__8213 (
            .O(N__43634),
            .I(N__43631));
    Span4Mux_h I__8212 (
            .O(N__43631),
            .I(N__43628));
    Span4Mux_h I__8211 (
            .O(N__43628),
            .I(N__43625));
    Odrv4 I__8210 (
            .O(N__43625),
            .I(\ALU.combOperand2_d_bmZ0Z_7 ));
    CascadeMux I__8209 (
            .O(N__43622),
            .I(\ALU.d_RNIM3JB6Z0Z_7_cascade_ ));
    CascadeMux I__8208 (
            .O(N__43619),
            .I(\ALU.dout_3_ns_1_7_cascade_ ));
    InMux I__8207 (
            .O(N__43616),
            .I(N__43613));
    LocalMux I__8206 (
            .O(N__43613),
            .I(\ALU.operand2_6_ns_1_7 ));
    InMux I__8205 (
            .O(N__43610),
            .I(N__43607));
    LocalMux I__8204 (
            .O(N__43607),
            .I(\ALU.N_606 ));
    CascadeMux I__8203 (
            .O(N__43604),
            .I(N__43600));
    InMux I__8202 (
            .O(N__43603),
            .I(N__43596));
    InMux I__8201 (
            .O(N__43600),
            .I(N__43591));
    InMux I__8200 (
            .O(N__43599),
            .I(N__43591));
    LocalMux I__8199 (
            .O(N__43596),
            .I(N__43585));
    LocalMux I__8198 (
            .O(N__43591),
            .I(N__43585));
    InMux I__8197 (
            .O(N__43590),
            .I(N__43582));
    Span4Mux_h I__8196 (
            .O(N__43585),
            .I(N__43579));
    LocalMux I__8195 (
            .O(N__43582),
            .I(\ALU.N_638 ));
    Odrv4 I__8194 (
            .O(N__43579),
            .I(\ALU.N_638 ));
    InMux I__8193 (
            .O(N__43574),
            .I(N__43568));
    InMux I__8192 (
            .O(N__43573),
            .I(N__43568));
    LocalMux I__8191 (
            .O(N__43568),
            .I(N__43565));
    Span4Mux_v I__8190 (
            .O(N__43565),
            .I(N__43562));
    Span4Mux_h I__8189 (
            .O(N__43562),
            .I(N__43559));
    Odrv4 I__8188 (
            .O(N__43559),
            .I(\ALU.a_15_m0_amZ0Z_2 ));
    CascadeMux I__8187 (
            .O(N__43556),
            .I(\ALU.a_15_m1_9_cascade_ ));
    InMux I__8186 (
            .O(N__43553),
            .I(N__43549));
    InMux I__8185 (
            .O(N__43552),
            .I(N__43546));
    LocalMux I__8184 (
            .O(N__43549),
            .I(N__43543));
    LocalMux I__8183 (
            .O(N__43546),
            .I(N__43540));
    Span4Mux_h I__8182 (
            .O(N__43543),
            .I(N__43535));
    Span4Mux_v I__8181 (
            .O(N__43540),
            .I(N__43535));
    Odrv4 I__8180 (
            .O(N__43535),
            .I(\ALU.aZ0Z_9 ));
    InMux I__8179 (
            .O(N__43532),
            .I(N__43526));
    InMux I__8178 (
            .O(N__43531),
            .I(N__43526));
    LocalMux I__8177 (
            .O(N__43526),
            .I(N__43523));
    Span4Mux_h I__8176 (
            .O(N__43523),
            .I(N__43520));
    Span4Mux_h I__8175 (
            .O(N__43520),
            .I(N__43517));
    Span4Mux_h I__8174 (
            .O(N__43517),
            .I(N__43514));
    Odrv4 I__8173 (
            .O(N__43514),
            .I(N_227_0));
    CascadeMux I__8172 (
            .O(N__43511),
            .I(N__43508));
    InMux I__8171 (
            .O(N__43508),
            .I(N__43502));
    InMux I__8170 (
            .O(N__43507),
            .I(N__43502));
    LocalMux I__8169 (
            .O(N__43502),
            .I(N__43499));
    Span4Mux_v I__8168 (
            .O(N__43499),
            .I(N__43496));
    Span4Mux_h I__8167 (
            .O(N__43496),
            .I(N__43491));
    InMux I__8166 (
            .O(N__43495),
            .I(N__43486));
    InMux I__8165 (
            .O(N__43494),
            .I(N__43486));
    Odrv4 I__8164 (
            .O(N__43491),
            .I(N_179));
    LocalMux I__8163 (
            .O(N__43486),
            .I(N_179));
    IoInMux I__8162 (
            .O(N__43481),
            .I(N__43478));
    LocalMux I__8161 (
            .O(N__43478),
            .I(N__43475));
    IoSpan4Mux I__8160 (
            .O(N__43475),
            .I(N__43471));
    IoInMux I__8159 (
            .O(N__43474),
            .I(N__43468));
    Span4Mux_s3_h I__8158 (
            .O(N__43471),
            .I(N__43465));
    LocalMux I__8157 (
            .O(N__43468),
            .I(N__43462));
    Sp12to4 I__8156 (
            .O(N__43465),
            .I(N__43459));
    Span12Mux_s6_h I__8155 (
            .O(N__43462),
            .I(N__43456));
    Span12Mux_h I__8154 (
            .O(N__43459),
            .I(N__43451));
    Span12Mux_h I__8153 (
            .O(N__43456),
            .I(N__43451));
    Odrv12 I__8152 (
            .O(N__43451),
            .I(bus_2));
    InMux I__8151 (
            .O(N__43448),
            .I(N__43445));
    LocalMux I__8150 (
            .O(N__43445),
            .I(N__43441));
    InMux I__8149 (
            .O(N__43444),
            .I(N__43438));
    Span12Mux_h I__8148 (
            .O(N__43441),
            .I(N__43435));
    LocalMux I__8147 (
            .O(N__43438),
            .I(\ALU.bZ0Z_4 ));
    Odrv12 I__8146 (
            .O(N__43435),
            .I(\ALU.bZ0Z_4 ));
    InMux I__8145 (
            .O(N__43430),
            .I(N__43427));
    LocalMux I__8144 (
            .O(N__43427),
            .I(N__43424));
    Span4Mux_h I__8143 (
            .O(N__43424),
            .I(N__43421));
    Span4Mux_h I__8142 (
            .O(N__43421),
            .I(N__43418));
    Odrv4 I__8141 (
            .O(N__43418),
            .I(\ALU.b_RNI5FSPZ0Z_4 ));
    InMux I__8140 (
            .O(N__43415),
            .I(N__43412));
    LocalMux I__8139 (
            .O(N__43412),
            .I(N__43409));
    Span4Mux_h I__8138 (
            .O(N__43409),
            .I(N__43406));
    Odrv4 I__8137 (
            .O(N__43406),
            .I(\ALU.c_RNIHV2SZ0Z_9 ));
    CascadeMux I__8136 (
            .O(N__43403),
            .I(N__43399));
    InMux I__8135 (
            .O(N__43402),
            .I(N__43396));
    InMux I__8134 (
            .O(N__43399),
            .I(N__43393));
    LocalMux I__8133 (
            .O(N__43396),
            .I(N__43390));
    LocalMux I__8132 (
            .O(N__43393),
            .I(N__43387));
    Span4Mux_v I__8131 (
            .O(N__43390),
            .I(N__43383));
    Span4Mux_v I__8130 (
            .O(N__43387),
            .I(N__43380));
    InMux I__8129 (
            .O(N__43386),
            .I(N__43377));
    Span4Mux_v I__8128 (
            .O(N__43383),
            .I(N__43374));
    Span4Mux_v I__8127 (
            .O(N__43380),
            .I(N__43371));
    LocalMux I__8126 (
            .O(N__43377),
            .I(N__43368));
    Span4Mux_h I__8125 (
            .O(N__43374),
            .I(N__43365));
    Span4Mux_h I__8124 (
            .O(N__43371),
            .I(N__43362));
    Span4Mux_v I__8123 (
            .O(N__43368),
            .I(N__43359));
    Sp12to4 I__8122 (
            .O(N__43365),
            .I(N__43356));
    Odrv4 I__8121 (
            .O(N__43362),
            .I(h_4));
    Odrv4 I__8120 (
            .O(N__43359),
            .I(h_4));
    Odrv12 I__8119 (
            .O(N__43356),
            .I(h_4));
    InMux I__8118 (
            .O(N__43349),
            .I(N__43345));
    InMux I__8117 (
            .O(N__43348),
            .I(N__43342));
    LocalMux I__8116 (
            .O(N__43345),
            .I(N__43339));
    LocalMux I__8115 (
            .O(N__43342),
            .I(N__43336));
    Span4Mux_h I__8114 (
            .O(N__43339),
            .I(N__43331));
    Span4Mux_v I__8113 (
            .O(N__43336),
            .I(N__43331));
    Span4Mux_h I__8112 (
            .O(N__43331),
            .I(N__43328));
    Odrv4 I__8111 (
            .O(N__43328),
            .I(\ALU.dZ0Z_4 ));
    InMux I__8110 (
            .O(N__43325),
            .I(N__43322));
    LocalMux I__8109 (
            .O(N__43322),
            .I(N__43319));
    Span4Mux_h I__8108 (
            .O(N__43319),
            .I(N__43316));
    Span4Mux_h I__8107 (
            .O(N__43316),
            .I(N__43313));
    Odrv4 I__8106 (
            .O(N__43313),
            .I(\ALU.d_RNI9R8EZ0Z_4 ));
    InMux I__8105 (
            .O(N__43310),
            .I(N__43300));
    InMux I__8104 (
            .O(N__43309),
            .I(N__43297));
    InMux I__8103 (
            .O(N__43308),
            .I(N__43288));
    InMux I__8102 (
            .O(N__43307),
            .I(N__43288));
    InMux I__8101 (
            .O(N__43306),
            .I(N__43280));
    InMux I__8100 (
            .O(N__43305),
            .I(N__43280));
    InMux I__8099 (
            .O(N__43304),
            .I(N__43280));
    InMux I__8098 (
            .O(N__43303),
            .I(N__43274));
    LocalMux I__8097 (
            .O(N__43300),
            .I(N__43269));
    LocalMux I__8096 (
            .O(N__43297),
            .I(N__43269));
    InMux I__8095 (
            .O(N__43296),
            .I(N__43260));
    InMux I__8094 (
            .O(N__43295),
            .I(N__43260));
    InMux I__8093 (
            .O(N__43294),
            .I(N__43260));
    InMux I__8092 (
            .O(N__43293),
            .I(N__43260));
    LocalMux I__8091 (
            .O(N__43288),
            .I(N__43257));
    InMux I__8090 (
            .O(N__43287),
            .I(N__43254));
    LocalMux I__8089 (
            .O(N__43280),
            .I(N__43251));
    InMux I__8088 (
            .O(N__43279),
            .I(N__43244));
    InMux I__8087 (
            .O(N__43278),
            .I(N__43244));
    InMux I__8086 (
            .O(N__43277),
            .I(N__43244));
    LocalMux I__8085 (
            .O(N__43274),
            .I(N__43239));
    Span4Mux_v I__8084 (
            .O(N__43269),
            .I(N__43234));
    LocalMux I__8083 (
            .O(N__43260),
            .I(N__43231));
    Span4Mux_v I__8082 (
            .O(N__43257),
            .I(N__43222));
    LocalMux I__8081 (
            .O(N__43254),
            .I(N__43222));
    Span4Mux_v I__8080 (
            .O(N__43251),
            .I(N__43222));
    LocalMux I__8079 (
            .O(N__43244),
            .I(N__43222));
    InMux I__8078 (
            .O(N__43243),
            .I(N__43217));
    InMux I__8077 (
            .O(N__43242),
            .I(N__43217));
    Span4Mux_v I__8076 (
            .O(N__43239),
            .I(N__43214));
    InMux I__8075 (
            .O(N__43238),
            .I(N__43209));
    InMux I__8074 (
            .O(N__43237),
            .I(N__43209));
    Span4Mux_h I__8073 (
            .O(N__43234),
            .I(N__43206));
    Span4Mux_v I__8072 (
            .O(N__43231),
            .I(N__43201));
    Span4Mux_h I__8071 (
            .O(N__43222),
            .I(N__43201));
    LocalMux I__8070 (
            .O(N__43217),
            .I(N__43198));
    Odrv4 I__8069 (
            .O(N__43214),
            .I(aluOperand2_2));
    LocalMux I__8068 (
            .O(N__43209),
            .I(aluOperand2_2));
    Odrv4 I__8067 (
            .O(N__43206),
            .I(aluOperand2_2));
    Odrv4 I__8066 (
            .O(N__43201),
            .I(aluOperand2_2));
    Odrv4 I__8065 (
            .O(N__43198),
            .I(aluOperand2_2));
    CascadeMux I__8064 (
            .O(N__43187),
            .I(\ALU.N_852_cascade_ ));
    InMux I__8063 (
            .O(N__43184),
            .I(N__43180));
    InMux I__8062 (
            .O(N__43183),
            .I(N__43177));
    LocalMux I__8061 (
            .O(N__43180),
            .I(N__43174));
    LocalMux I__8060 (
            .O(N__43177),
            .I(\ALU.N_966 ));
    Odrv4 I__8059 (
            .O(N__43174),
            .I(\ALU.N_966 ));
    CascadeMux I__8058 (
            .O(N__43169),
            .I(\ALU.N_766_cascade_ ));
    InMux I__8057 (
            .O(N__43166),
            .I(N__43161));
    CascadeMux I__8056 (
            .O(N__43165),
            .I(N__43157));
    CascadeMux I__8055 (
            .O(N__43164),
            .I(N__43154));
    LocalMux I__8054 (
            .O(N__43161),
            .I(N__43151));
    InMux I__8053 (
            .O(N__43160),
            .I(N__43146));
    InMux I__8052 (
            .O(N__43157),
            .I(N__43146));
    InMux I__8051 (
            .O(N__43154),
            .I(N__43143));
    Span12Mux_h I__8050 (
            .O(N__43151),
            .I(N__43140));
    LocalMux I__8049 (
            .O(N__43146),
            .I(N__43137));
    LocalMux I__8048 (
            .O(N__43143),
            .I(N__43134));
    Odrv12 I__8047 (
            .O(N__43140),
            .I(\ALU.N_634 ));
    Odrv4 I__8046 (
            .O(N__43137),
            .I(\ALU.N_634 ));
    Odrv12 I__8045 (
            .O(N__43134),
            .I(\ALU.N_634 ));
    CascadeMux I__8044 (
            .O(N__43127),
            .I(\ALU.N_634_cascade_ ));
    CascadeMux I__8043 (
            .O(N__43124),
            .I(\ALU.N_811_cascade_ ));
    InMux I__8042 (
            .O(N__43121),
            .I(N__43115));
    InMux I__8041 (
            .O(N__43120),
            .I(N__43112));
    InMux I__8040 (
            .O(N__43119),
            .I(N__43109));
    InMux I__8039 (
            .O(N__43118),
            .I(N__43106));
    LocalMux I__8038 (
            .O(N__43115),
            .I(N__43101));
    LocalMux I__8037 (
            .O(N__43112),
            .I(N__43096));
    LocalMux I__8036 (
            .O(N__43109),
            .I(N__43096));
    LocalMux I__8035 (
            .O(N__43106),
            .I(N__43093));
    InMux I__8034 (
            .O(N__43105),
            .I(N__43090));
    InMux I__8033 (
            .O(N__43104),
            .I(N__43087));
    Span4Mux_h I__8032 (
            .O(N__43101),
            .I(N__43075));
    Span4Mux_v I__8031 (
            .O(N__43096),
            .I(N__43075));
    Span4Mux_v I__8030 (
            .O(N__43093),
            .I(N__43075));
    LocalMux I__8029 (
            .O(N__43090),
            .I(N__43075));
    LocalMux I__8028 (
            .O(N__43087),
            .I(N__43075));
    InMux I__8027 (
            .O(N__43086),
            .I(N__43072));
    Odrv4 I__8026 (
            .O(N__43075),
            .I(\ALU.d_RNIK8M6K5Z0Z_6 ));
    LocalMux I__8025 (
            .O(N__43072),
            .I(\ALU.d_RNIK8M6K5Z0Z_6 ));
    InMux I__8024 (
            .O(N__43067),
            .I(N__43062));
    InMux I__8023 (
            .O(N__43066),
            .I(N__43059));
    InMux I__8022 (
            .O(N__43065),
            .I(N__43056));
    LocalMux I__8021 (
            .O(N__43062),
            .I(N__43052));
    LocalMux I__8020 (
            .O(N__43059),
            .I(N__43048));
    LocalMux I__8019 (
            .O(N__43056),
            .I(N__43045));
    InMux I__8018 (
            .O(N__43055),
            .I(N__43042));
    Span4Mux_h I__8017 (
            .O(N__43052),
            .I(N__43034));
    InMux I__8016 (
            .O(N__43051),
            .I(N__43031));
    Span4Mux_v I__8015 (
            .O(N__43048),
            .I(N__43024));
    Span4Mux_v I__8014 (
            .O(N__43045),
            .I(N__43024));
    LocalMux I__8013 (
            .O(N__43042),
            .I(N__43024));
    InMux I__8012 (
            .O(N__43041),
            .I(N__43021));
    InMux I__8011 (
            .O(N__43040),
            .I(N__43018));
    InMux I__8010 (
            .O(N__43039),
            .I(N__43015));
    InMux I__8009 (
            .O(N__43038),
            .I(N__43010));
    InMux I__8008 (
            .O(N__43037),
            .I(N__43010));
    Odrv4 I__8007 (
            .O(N__43034),
            .I(\ALU.a_15_sZ0Z_11 ));
    LocalMux I__8006 (
            .O(N__43031),
            .I(\ALU.a_15_sZ0Z_11 ));
    Odrv4 I__8005 (
            .O(N__43024),
            .I(\ALU.a_15_sZ0Z_11 ));
    LocalMux I__8004 (
            .O(N__43021),
            .I(\ALU.a_15_sZ0Z_11 ));
    LocalMux I__8003 (
            .O(N__43018),
            .I(\ALU.a_15_sZ0Z_11 ));
    LocalMux I__8002 (
            .O(N__43015),
            .I(\ALU.a_15_sZ0Z_11 ));
    LocalMux I__8001 (
            .O(N__43010),
            .I(\ALU.a_15_sZ0Z_11 ));
    CascadeMux I__8000 (
            .O(N__42995),
            .I(\ALU.d_RNIK8M6K5Z0Z_6_cascade_ ));
    InMux I__7999 (
            .O(N__42992),
            .I(N__42987));
    InMux I__7998 (
            .O(N__42991),
            .I(N__42984));
    InMux I__7997 (
            .O(N__42990),
            .I(N__42979));
    LocalMux I__7996 (
            .O(N__42987),
            .I(N__42974));
    LocalMux I__7995 (
            .O(N__42984),
            .I(N__42971));
    InMux I__7994 (
            .O(N__42983),
            .I(N__42968));
    InMux I__7993 (
            .O(N__42982),
            .I(N__42965));
    LocalMux I__7992 (
            .O(N__42979),
            .I(N__42962));
    InMux I__7991 (
            .O(N__42978),
            .I(N__42959));
    InMux I__7990 (
            .O(N__42977),
            .I(N__42956));
    Odrv4 I__7989 (
            .O(N__42974),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0 ));
    Odrv4 I__7988 (
            .O(N__42971),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0 ));
    LocalMux I__7987 (
            .O(N__42968),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0 ));
    LocalMux I__7986 (
            .O(N__42965),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0 ));
    Odrv12 I__7985 (
            .O(N__42962),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0 ));
    LocalMux I__7984 (
            .O(N__42959),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0 ));
    LocalMux I__7983 (
            .O(N__42956),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0 ));
    InMux I__7982 (
            .O(N__42941),
            .I(N__42938));
    LocalMux I__7981 (
            .O(N__42938),
            .I(N__42934));
    InMux I__7980 (
            .O(N__42937),
            .I(N__42931));
    Span4Mux_v I__7979 (
            .O(N__42934),
            .I(N__42928));
    LocalMux I__7978 (
            .O(N__42931),
            .I(N__42925));
    Span4Mux_h I__7977 (
            .O(N__42928),
            .I(N__42922));
    Span4Mux_v I__7976 (
            .O(N__42925),
            .I(N__42919));
    Span4Mux_h I__7975 (
            .O(N__42922),
            .I(N__42916));
    Span4Mux_h I__7974 (
            .O(N__42919),
            .I(N__42913));
    Odrv4 I__7973 (
            .O(N__42916),
            .I(\ALU.aZ0Z_6 ));
    Odrv4 I__7972 (
            .O(N__42913),
            .I(\ALU.aZ0Z_6 ));
    InMux I__7971 (
            .O(N__42908),
            .I(N__42905));
    LocalMux I__7970 (
            .O(N__42905),
            .I(\ALU.N_766 ));
    CascadeMux I__7969 (
            .O(N__42902),
            .I(\ALU.N_606_cascade_ ));
    InMux I__7968 (
            .O(N__42899),
            .I(N__42896));
    LocalMux I__7967 (
            .O(N__42896),
            .I(N__42893));
    Span4Mux_h I__7966 (
            .O(N__42893),
            .I(N__42890));
    Odrv4 I__7965 (
            .O(N__42890),
            .I(\ALU.addsub_axb_1_1 ));
    InMux I__7964 (
            .O(N__42887),
            .I(N__42884));
    LocalMux I__7963 (
            .O(N__42884),
            .I(\ALU.N_1026 ));
    InMux I__7962 (
            .O(N__42881),
            .I(N__42878));
    LocalMux I__7961 (
            .O(N__42878),
            .I(N__42875));
    Odrv4 I__7960 (
            .O(N__42875),
            .I(\ALU.mult_293_c_RNOZ0Z_0 ));
    CascadeMux I__7959 (
            .O(N__42872),
            .I(N__42869));
    InMux I__7958 (
            .O(N__42869),
            .I(N__42865));
    InMux I__7957 (
            .O(N__42868),
            .I(N__42862));
    LocalMux I__7956 (
            .O(N__42865),
            .I(N__42859));
    LocalMux I__7955 (
            .O(N__42862),
            .I(\ALU.N_1011 ));
    Odrv4 I__7954 (
            .O(N__42859),
            .I(\ALU.N_1011 ));
    InMux I__7953 (
            .O(N__42854),
            .I(N__42851));
    LocalMux I__7952 (
            .O(N__42851),
            .I(\ALU.mult_323_c_RNIAA0BZ0Z82 ));
    InMux I__7951 (
            .O(N__42848),
            .I(N__42845));
    LocalMux I__7950 (
            .O(N__42845),
            .I(\ALU.d_RNIGD2441Z0Z_8 ));
    CascadeMux I__7949 (
            .O(N__42842),
            .I(\ALU.N_639_cascade_ ));
    InMux I__7948 (
            .O(N__42839),
            .I(N__42836));
    LocalMux I__7947 (
            .O(N__42836),
            .I(N__42833));
    Span4Mux_v I__7946 (
            .O(N__42833),
            .I(N__42830));
    Sp12to4 I__7945 (
            .O(N__42830),
            .I(N__42827));
    Odrv12 I__7944 (
            .O(N__42827),
            .I(\ALU.d_RNIC6EBM2Z0Z_2 ));
    CascadeMux I__7943 (
            .O(N__42824),
            .I(\ALU.d_RNIFVCT15Z0Z_8_cascade_ ));
    InMux I__7942 (
            .O(N__42821),
            .I(N__42818));
    LocalMux I__7941 (
            .O(N__42818),
            .I(\ALU.lshift_11 ));
    InMux I__7940 (
            .O(N__42815),
            .I(N__42812));
    LocalMux I__7939 (
            .O(N__42812),
            .I(N__42807));
    InMux I__7938 (
            .O(N__42811),
            .I(N__42802));
    InMux I__7937 (
            .O(N__42810),
            .I(N__42802));
    Odrv4 I__7936 (
            .O(N__42807),
            .I(\ALU.N_851 ));
    LocalMux I__7935 (
            .O(N__42802),
            .I(\ALU.N_851 ));
    CascadeMux I__7934 (
            .O(N__42797),
            .I(\ALU.N_851_cascade_ ));
    InMux I__7933 (
            .O(N__42794),
            .I(N__42791));
    LocalMux I__7932 (
            .O(N__42791),
            .I(\ALU.c_RNINT9PO2_0Z0Z_10 ));
    InMux I__7931 (
            .O(N__42788),
            .I(N__42782));
    InMux I__7930 (
            .O(N__42787),
            .I(N__42782));
    LocalMux I__7929 (
            .O(N__42782),
            .I(\ALU.N_978 ));
    CascadeMux I__7928 (
            .O(N__42779),
            .I(\ALU.N_978_cascade_ ));
    InMux I__7927 (
            .O(N__42776),
            .I(N__42773));
    LocalMux I__7926 (
            .O(N__42773),
            .I(N__42769));
    InMux I__7925 (
            .O(N__42772),
            .I(N__42766));
    Span4Mux_h I__7924 (
            .O(N__42769),
            .I(N__42763));
    LocalMux I__7923 (
            .O(N__42766),
            .I(N__42758));
    Span4Mux_h I__7922 (
            .O(N__42763),
            .I(N__42758));
    Odrv4 I__7921 (
            .O(N__42758),
            .I(\ALU.N_836 ));
    CascadeMux I__7920 (
            .O(N__42755),
            .I(N__42752));
    InMux I__7919 (
            .O(N__42752),
            .I(N__42749));
    LocalMux I__7918 (
            .O(N__42749),
            .I(N__42746));
    Span4Mux_v I__7917 (
            .O(N__42746),
            .I(N__42743));
    Odrv4 I__7916 (
            .O(N__42743),
            .I(\ALU.mult_293_c_RNOZ0 ));
    InMux I__7915 (
            .O(N__42740),
            .I(N__42737));
    LocalMux I__7914 (
            .O(N__42737),
            .I(N__42734));
    Span4Mux_v I__7913 (
            .O(N__42734),
            .I(N__42731));
    Odrv4 I__7912 (
            .O(N__42731),
            .I(\ALU.d_RNI34ECOZ0Z_9 ));
    CascadeMux I__7911 (
            .O(N__42728),
            .I(N__42725));
    InMux I__7910 (
            .O(N__42725),
            .I(N__42722));
    LocalMux I__7909 (
            .O(N__42722),
            .I(N__42719));
    Span4Mux_h I__7908 (
            .O(N__42719),
            .I(N__42716));
    Span4Mux_h I__7907 (
            .O(N__42716),
            .I(N__42713));
    Odrv4 I__7906 (
            .O(N__42713),
            .I(\ALU.d_RNI0PI3E1Z0Z_8 ));
    InMux I__7905 (
            .O(N__42710),
            .I(N__42707));
    LocalMux I__7904 (
            .O(N__42707),
            .I(\ALU.mult_9_10 ));
    InMux I__7903 (
            .O(N__42704),
            .I(\ALU.mult_9_c9 ));
    InMux I__7902 (
            .O(N__42701),
            .I(N__42698));
    LocalMux I__7901 (
            .O(N__42698),
            .I(\ALU.d_RNIFCNKLZ0Z_9 ));
    CascadeMux I__7900 (
            .O(N__42695),
            .I(N__42692));
    InMux I__7899 (
            .O(N__42692),
            .I(N__42689));
    LocalMux I__7898 (
            .O(N__42689),
            .I(N__42686));
    Odrv4 I__7897 (
            .O(N__42686),
            .I(\ALU.d_RNIDR5C61Z0Z_8 ));
    InMux I__7896 (
            .O(N__42683),
            .I(N__42680));
    LocalMux I__7895 (
            .O(N__42680),
            .I(\ALU.mult_9_11 ));
    InMux I__7894 (
            .O(N__42677),
            .I(\ALU.mult_9_c10 ));
    CascadeMux I__7893 (
            .O(N__42674),
            .I(N__42671));
    InMux I__7892 (
            .O(N__42671),
            .I(N__42668));
    LocalMux I__7891 (
            .O(N__42668),
            .I(\ALU.d_RNIG61LGZ0Z_9 ));
    InMux I__7890 (
            .O(N__42665),
            .I(N__42662));
    LocalMux I__7889 (
            .O(N__42662),
            .I(\ALU.mult_9_12 ));
    InMux I__7888 (
            .O(N__42659),
            .I(\ALU.mult_9_c11 ));
    CascadeMux I__7887 (
            .O(N__42656),
            .I(N__42653));
    InMux I__7886 (
            .O(N__42653),
            .I(N__42650));
    LocalMux I__7885 (
            .O(N__42650),
            .I(N__42647));
    Span4Mux_h I__7884 (
            .O(N__42647),
            .I(N__42644));
    Odrv4 I__7883 (
            .O(N__42644),
            .I(\ALU.d_RNI68LSHZ0Z_9 ));
    InMux I__7882 (
            .O(N__42641),
            .I(N__42638));
    LocalMux I__7881 (
            .O(N__42638),
            .I(\ALU.mult_9_13 ));
    InMux I__7880 (
            .O(N__42635),
            .I(\ALU.mult_9_c12 ));
    InMux I__7879 (
            .O(N__42632),
            .I(N__42629));
    LocalMux I__7878 (
            .O(N__42629),
            .I(N__42626));
    Span4Mux_v I__7877 (
            .O(N__42626),
            .I(N__42623));
    Sp12to4 I__7876 (
            .O(N__42623),
            .I(N__42620));
    Odrv12 I__7875 (
            .O(N__42620),
            .I(\ALU.d_RNISSV4IZ0Z_9 ));
    CascadeMux I__7874 (
            .O(N__42617),
            .I(N__42614));
    InMux I__7873 (
            .O(N__42614),
            .I(N__42611));
    LocalMux I__7872 (
            .O(N__42611),
            .I(N__42608));
    Span12Mux_h I__7871 (
            .O(N__42608),
            .I(N__42605));
    Odrv12 I__7870 (
            .O(N__42605),
            .I(\ALU.d_RNI371041Z0Z_8 ));
    InMux I__7869 (
            .O(N__42602),
            .I(N__42599));
    LocalMux I__7868 (
            .O(N__42599),
            .I(\ALU.mult_9_14 ));
    InMux I__7867 (
            .O(N__42596),
            .I(\ALU.mult_9_c13 ));
    InMux I__7866 (
            .O(N__42593),
            .I(N__42590));
    LocalMux I__7865 (
            .O(N__42590),
            .I(N__42587));
    Span4Mux_h I__7864 (
            .O(N__42587),
            .I(N__42584));
    Span4Mux_h I__7863 (
            .O(N__42584),
            .I(N__42581));
    Odrv4 I__7862 (
            .O(N__42581),
            .I(\ALU.c_RNI0QV651Z0Z_10 ));
    InMux I__7861 (
            .O(N__42578),
            .I(\ALU.mult_9_c14 ));
    InMux I__7860 (
            .O(N__42575),
            .I(N__42572));
    LocalMux I__7859 (
            .O(N__42572),
            .I(\ALU.N_862 ));
    CascadeMux I__7858 (
            .O(N__42569),
            .I(\ALU.N_862_cascade_ ));
    CascadeMux I__7857 (
            .O(N__42566),
            .I(\ALU.N_922_cascade_ ));
    InMux I__7856 (
            .O(N__42563),
            .I(N__42560));
    LocalMux I__7855 (
            .O(N__42560),
            .I(N__42557));
    Span4Mux_h I__7854 (
            .O(N__42557),
            .I(N__42554));
    Odrv4 I__7853 (
            .O(N__42554),
            .I(\ALU.d_RNIR6J013Z0Z_2 ));
    InMux I__7852 (
            .O(N__42551),
            .I(N__42543));
    InMux I__7851 (
            .O(N__42550),
            .I(N__42540));
    InMux I__7850 (
            .O(N__42549),
            .I(N__42537));
    InMux I__7849 (
            .O(N__42548),
            .I(N__42533));
    InMux I__7848 (
            .O(N__42547),
            .I(N__42530));
    InMux I__7847 (
            .O(N__42546),
            .I(N__42526));
    LocalMux I__7846 (
            .O(N__42543),
            .I(N__42523));
    LocalMux I__7845 (
            .O(N__42540),
            .I(N__42520));
    LocalMux I__7844 (
            .O(N__42537),
            .I(N__42517));
    InMux I__7843 (
            .O(N__42536),
            .I(N__42514));
    LocalMux I__7842 (
            .O(N__42533),
            .I(N__42509));
    LocalMux I__7841 (
            .O(N__42530),
            .I(N__42509));
    InMux I__7840 (
            .O(N__42529),
            .I(N__42506));
    LocalMux I__7839 (
            .O(N__42526),
            .I(N__42501));
    Span4Mux_h I__7838 (
            .O(N__42523),
            .I(N__42501));
    Span4Mux_v I__7837 (
            .O(N__42520),
            .I(N__42498));
    Span4Mux_v I__7836 (
            .O(N__42517),
            .I(N__42495));
    LocalMux I__7835 (
            .O(N__42514),
            .I(N__42490));
    Span4Mux_v I__7834 (
            .O(N__42509),
            .I(N__42490));
    LocalMux I__7833 (
            .O(N__42506),
            .I(N__42485));
    Span4Mux_h I__7832 (
            .O(N__42501),
            .I(N__42485));
    Span4Mux_h I__7831 (
            .O(N__42498),
            .I(N__42482));
    Span4Mux_h I__7830 (
            .O(N__42495),
            .I(N__42477));
    Span4Mux_v I__7829 (
            .O(N__42490),
            .I(N__42477));
    Span4Mux_v I__7828 (
            .O(N__42485),
            .I(N__42474));
    Span4Mux_h I__7827 (
            .O(N__42482),
            .I(N__42471));
    Odrv4 I__7826 (
            .O(N__42477),
            .I(\ALU.d_RNI1AHUF8Z0Z_2 ));
    Odrv4 I__7825 (
            .O(N__42474),
            .I(\ALU.d_RNI1AHUF8Z0Z_2 ));
    Odrv4 I__7824 (
            .O(N__42471),
            .I(\ALU.d_RNI1AHUF8Z0Z_2 ));
    InMux I__7823 (
            .O(N__42464),
            .I(N__42460));
    CascadeMux I__7822 (
            .O(N__42463),
            .I(N__42457));
    LocalMux I__7821 (
            .O(N__42460),
            .I(N__42454));
    InMux I__7820 (
            .O(N__42457),
            .I(N__42451));
    Odrv12 I__7819 (
            .O(N__42454),
            .I(\ALU.mult_25_10 ));
    LocalMux I__7818 (
            .O(N__42451),
            .I(\ALU.mult_25_10 ));
    CascadeMux I__7817 (
            .O(N__42446),
            .I(N__42443));
    InMux I__7816 (
            .O(N__42443),
            .I(N__42440));
    LocalMux I__7815 (
            .O(N__42440),
            .I(\ALU.mult_11_10 ));
    InMux I__7814 (
            .O(N__42437),
            .I(N__42434));
    LocalMux I__7813 (
            .O(N__42434),
            .I(N__42431));
    Span4Mux_h I__7812 (
            .O(N__42431),
            .I(N__42428));
    Odrv4 I__7811 (
            .O(N__42428),
            .I(\ALU.mult_293_c_RNIOCJMDZ0Z9 ));
    CascadeMux I__7810 (
            .O(N__42425),
            .I(N__42422));
    InMux I__7809 (
            .O(N__42422),
            .I(N__42419));
    LocalMux I__7808 (
            .O(N__42419),
            .I(\ALU.mult_11_11 ));
    InMux I__7807 (
            .O(N__42416),
            .I(N__42413));
    LocalMux I__7806 (
            .O(N__42413),
            .I(N__42410));
    Span4Mux_h I__7805 (
            .O(N__42410),
            .I(N__42407));
    Odrv4 I__7804 (
            .O(N__42407),
            .I(\ALU.mult_21_11 ));
    InMux I__7803 (
            .O(N__42404),
            .I(\ALU.mult_21_c10 ));
    InMux I__7802 (
            .O(N__42401),
            .I(N__42397));
    InMux I__7801 (
            .O(N__42400),
            .I(N__42394));
    LocalMux I__7800 (
            .O(N__42397),
            .I(\ALU.mult_21_12 ));
    LocalMux I__7799 (
            .O(N__42394),
            .I(\ALU.mult_21_12 ));
    InMux I__7798 (
            .O(N__42389),
            .I(\ALU.mult_21_c11 ));
    InMux I__7797 (
            .O(N__42386),
            .I(N__42383));
    LocalMux I__7796 (
            .O(N__42383),
            .I(\ALU.mult_21_13 ));
    InMux I__7795 (
            .O(N__42380),
            .I(\ALU.mult_21_c12 ));
    CascadeMux I__7794 (
            .O(N__42377),
            .I(N__42374));
    InMux I__7793 (
            .O(N__42374),
            .I(N__42371));
    LocalMux I__7792 (
            .O(N__42371),
            .I(N__42367));
    InMux I__7791 (
            .O(N__42370),
            .I(N__42364));
    Odrv4 I__7790 (
            .O(N__42367),
            .I(\ALU.mult_21_14 ));
    LocalMux I__7789 (
            .O(N__42364),
            .I(\ALU.mult_21_14 ));
    InMux I__7788 (
            .O(N__42359),
            .I(\ALU.mult_21_c13 ));
    InMux I__7787 (
            .O(N__42356),
            .I(N__42353));
    LocalMux I__7786 (
            .O(N__42353),
            .I(\ALU.mult_23_15 ));
    InMux I__7785 (
            .O(N__42350),
            .I(\ALU.mult_21_c14 ));
    InMux I__7784 (
            .O(N__42347),
            .I(N__42344));
    LocalMux I__7783 (
            .O(N__42344),
            .I(N__42341));
    Span4Mux_v I__7782 (
            .O(N__42341),
            .I(N__42338));
    Odrv4 I__7781 (
            .O(N__42338),
            .I(\ALU.mult_476_c_RNIFLP0OZ0Z7 ));
    InMux I__7780 (
            .O(N__42335),
            .I(N__42329));
    InMux I__7779 (
            .O(N__42334),
            .I(N__42329));
    LocalMux I__7778 (
            .O(N__42329),
            .I(N__42326));
    Span4Mux_h I__7777 (
            .O(N__42326),
            .I(N__42323));
    Span4Mux_h I__7776 (
            .O(N__42323),
            .I(N__42319));
    CascadeMux I__7775 (
            .O(N__42322),
            .I(N__42316));
    Span4Mux_h I__7774 (
            .O(N__42319),
            .I(N__42313));
    InMux I__7773 (
            .O(N__42316),
            .I(N__42310));
    Odrv4 I__7772 (
            .O(N__42313),
            .I(\CONTROL.addrstack_1_7 ));
    LocalMux I__7771 (
            .O(N__42310),
            .I(\CONTROL.addrstack_1_7 ));
    InMux I__7770 (
            .O(N__42305),
            .I(N__42299));
    InMux I__7769 (
            .O(N__42304),
            .I(N__42299));
    LocalMux I__7768 (
            .O(N__42299),
            .I(\CONTROL.g0_4Z0Z_2 ));
    CascadeMux I__7767 (
            .O(N__42296),
            .I(\CONTROL.g0_i_m2_1_cascade_ ));
    InMux I__7766 (
            .O(N__42293),
            .I(N__42290));
    LocalMux I__7765 (
            .O(N__42290),
            .I(\CONTROL.g1_1 ));
    InMux I__7764 (
            .O(N__42287),
            .I(N__42284));
    LocalMux I__7763 (
            .O(N__42284),
            .I(N__42281));
    Span4Mux_v I__7762 (
            .O(N__42281),
            .I(N__42277));
    InMux I__7761 (
            .O(N__42280),
            .I(N__42274));
    Sp12to4 I__7760 (
            .O(N__42277),
            .I(N__42271));
    LocalMux I__7759 (
            .O(N__42274),
            .I(\CONTROL.addrstackptrZ0Z_7 ));
    Odrv12 I__7758 (
            .O(N__42271),
            .I(\CONTROL.addrstackptrZ0Z_7 ));
    InMux I__7757 (
            .O(N__42266),
            .I(N__42258));
    InMux I__7756 (
            .O(N__42265),
            .I(N__42255));
    InMux I__7755 (
            .O(N__42264),
            .I(N__42250));
    InMux I__7754 (
            .O(N__42263),
            .I(N__42250));
    CascadeMux I__7753 (
            .O(N__42262),
            .I(N__42245));
    InMux I__7752 (
            .O(N__42261),
            .I(N__42241));
    LocalMux I__7751 (
            .O(N__42258),
            .I(N__42236));
    LocalMux I__7750 (
            .O(N__42255),
            .I(N__42236));
    LocalMux I__7749 (
            .O(N__42250),
            .I(N__42232));
    InMux I__7748 (
            .O(N__42249),
            .I(N__42225));
    InMux I__7747 (
            .O(N__42248),
            .I(N__42225));
    InMux I__7746 (
            .O(N__42245),
            .I(N__42225));
    InMux I__7745 (
            .O(N__42244),
            .I(N__42222));
    LocalMux I__7744 (
            .O(N__42241),
            .I(N__42217));
    Span4Mux_h I__7743 (
            .O(N__42236),
            .I(N__42213));
    CascadeMux I__7742 (
            .O(N__42235),
            .I(N__42209));
    Span4Mux_h I__7741 (
            .O(N__42232),
            .I(N__42203));
    LocalMux I__7740 (
            .O(N__42225),
            .I(N__42203));
    LocalMux I__7739 (
            .O(N__42222),
            .I(N__42200));
    InMux I__7738 (
            .O(N__42221),
            .I(N__42197));
    CascadeMux I__7737 (
            .O(N__42220),
            .I(N__42192));
    Span4Mux_h I__7736 (
            .O(N__42217),
            .I(N__42189));
    InMux I__7735 (
            .O(N__42216),
            .I(N__42186));
    Span4Mux_h I__7734 (
            .O(N__42213),
            .I(N__42183));
    InMux I__7733 (
            .O(N__42212),
            .I(N__42176));
    InMux I__7732 (
            .O(N__42209),
            .I(N__42176));
    InMux I__7731 (
            .O(N__42208),
            .I(N__42176));
    Span4Mux_h I__7730 (
            .O(N__42203),
            .I(N__42169));
    Span4Mux_h I__7729 (
            .O(N__42200),
            .I(N__42169));
    LocalMux I__7728 (
            .O(N__42197),
            .I(N__42169));
    InMux I__7727 (
            .O(N__42196),
            .I(N__42162));
    InMux I__7726 (
            .O(N__42195),
            .I(N__42162));
    InMux I__7725 (
            .O(N__42192),
            .I(N__42162));
    Odrv4 I__7724 (
            .O(N__42189),
            .I(PROM_ROMDATA_dintern_5ro));
    LocalMux I__7723 (
            .O(N__42186),
            .I(PROM_ROMDATA_dintern_5ro));
    Odrv4 I__7722 (
            .O(N__42183),
            .I(PROM_ROMDATA_dintern_5ro));
    LocalMux I__7721 (
            .O(N__42176),
            .I(PROM_ROMDATA_dintern_5ro));
    Odrv4 I__7720 (
            .O(N__42169),
            .I(PROM_ROMDATA_dintern_5ro));
    LocalMux I__7719 (
            .O(N__42162),
            .I(PROM_ROMDATA_dintern_5ro));
    InMux I__7718 (
            .O(N__42149),
            .I(N__42146));
    LocalMux I__7717 (
            .O(N__42146),
            .I(N__42143));
    Span4Mux_h I__7716 (
            .O(N__42143),
            .I(N__42140));
    Odrv4 I__7715 (
            .O(N__42140),
            .I(\CONTROL.g0_2_iZ0Z_1 ));
    InMux I__7714 (
            .O(N__42137),
            .I(N__42134));
    LocalMux I__7713 (
            .O(N__42134),
            .I(\PROM.ROMDATA.m381_am ));
    InMux I__7712 (
            .O(N__42131),
            .I(N__42128));
    LocalMux I__7711 (
            .O(N__42128),
            .I(N__42125));
    Span4Mux_h I__7710 (
            .O(N__42125),
            .I(N__42122));
    Odrv4 I__7709 (
            .O(N__42122),
            .I(\PROM.ROMDATA.m375_am ));
    InMux I__7708 (
            .O(N__42119),
            .I(N__42116));
    LocalMux I__7707 (
            .O(N__42116),
            .I(\PROM.ROMDATA.m382_ns_1 ));
    CascadeMux I__7706 (
            .O(N__42113),
            .I(N__42110));
    InMux I__7705 (
            .O(N__42110),
            .I(N__42107));
    LocalMux I__7704 (
            .O(N__42107),
            .I(N__42104));
    Span4Mux_h I__7703 (
            .O(N__42104),
            .I(N__42101));
    Span4Mux_h I__7702 (
            .O(N__42101),
            .I(N__42098));
    Odrv4 I__7701 (
            .O(N__42098),
            .I(\ALU.rshift_3_ns_1_0 ));
    CascadeMux I__7700 (
            .O(N__42095),
            .I(\ALU.N_858_cascade_ ));
    CascadeMux I__7699 (
            .O(N__42092),
            .I(\ALU.rshift_15_ns_1_0_cascade_ ));
    CascadeMux I__7698 (
            .O(N__42089),
            .I(\ALU.rshift_3_ns_1_4_cascade_ ));
    InMux I__7697 (
            .O(N__42086),
            .I(N__42083));
    LocalMux I__7696 (
            .O(N__42083),
            .I(N__42077));
    InMux I__7695 (
            .O(N__42082),
            .I(N__42074));
    InMux I__7694 (
            .O(N__42081),
            .I(N__42071));
    InMux I__7693 (
            .O(N__42080),
            .I(N__42067));
    Span4Mux_v I__7692 (
            .O(N__42077),
            .I(N__42060));
    LocalMux I__7691 (
            .O(N__42074),
            .I(N__42060));
    LocalMux I__7690 (
            .O(N__42071),
            .I(N__42060));
    InMux I__7689 (
            .O(N__42070),
            .I(N__42057));
    LocalMux I__7688 (
            .O(N__42067),
            .I(N__42054));
    Span4Mux_h I__7687 (
            .O(N__42060),
            .I(N__42049));
    LocalMux I__7686 (
            .O(N__42057),
            .I(N__42049));
    Odrv12 I__7685 (
            .O(N__42054),
            .I(\CONTROL.un1_programCounter9_reto_rep1 ));
    Odrv4 I__7684 (
            .O(N__42049),
            .I(\CONTROL.un1_programCounter9_reto_rep1 ));
    InMux I__7683 (
            .O(N__42044),
            .I(N__42041));
    LocalMux I__7682 (
            .O(N__42041),
            .I(N__42038));
    Span4Mux_v I__7681 (
            .O(N__42038),
            .I(N__42035));
    Span4Mux_h I__7680 (
            .O(N__42035),
            .I(N__42032));
    Span4Mux_h I__7679 (
            .O(N__42032),
            .I(N__42029));
    Odrv4 I__7678 (
            .O(N__42029),
            .I(\CONTROL.g0_2Z0Z_1 ));
    InMux I__7677 (
            .O(N__42026),
            .I(N__42023));
    LocalMux I__7676 (
            .O(N__42023),
            .I(N__42020));
    Odrv4 I__7675 (
            .O(N__42020),
            .I(\CONTROL.N_133_0_0 ));
    InMux I__7674 (
            .O(N__42017),
            .I(N__42014));
    LocalMux I__7673 (
            .O(N__42014),
            .I(\CONTROL.N_114_i ));
    CascadeMux I__7672 (
            .O(N__42011),
            .I(N__42008));
    InMux I__7671 (
            .O(N__42008),
            .I(N__42005));
    LocalMux I__7670 (
            .O(N__42005),
            .I(N__42002));
    Span4Mux_v I__7669 (
            .O(N__42002),
            .I(N__41999));
    Span4Mux_h I__7668 (
            .O(N__41999),
            .I(N__41996));
    Span4Mux_h I__7667 (
            .O(N__41996),
            .I(N__41993));
    Odrv4 I__7666 (
            .O(N__41993),
            .I(\CONTROL.g1_1_4 ));
    InMux I__7665 (
            .O(N__41990),
            .I(N__41987));
    LocalMux I__7664 (
            .O(N__41987),
            .I(N__41983));
    InMux I__7663 (
            .O(N__41986),
            .I(N__41978));
    Span4Mux_v I__7662 (
            .O(N__41983),
            .I(N__41973));
    InMux I__7661 (
            .O(N__41982),
            .I(N__41970));
    InMux I__7660 (
            .O(N__41981),
            .I(N__41967));
    LocalMux I__7659 (
            .O(N__41978),
            .I(N__41964));
    InMux I__7658 (
            .O(N__41977),
            .I(N__41961));
    InMux I__7657 (
            .O(N__41976),
            .I(N__41955));
    Span4Mux_v I__7656 (
            .O(N__41973),
            .I(N__41952));
    LocalMux I__7655 (
            .O(N__41970),
            .I(N__41949));
    LocalMux I__7654 (
            .O(N__41967),
            .I(N__41946));
    Span4Mux_h I__7653 (
            .O(N__41964),
            .I(N__41941));
    LocalMux I__7652 (
            .O(N__41961),
            .I(N__41941));
    InMux I__7651 (
            .O(N__41960),
            .I(N__41938));
    InMux I__7650 (
            .O(N__41959),
            .I(N__41933));
    InMux I__7649 (
            .O(N__41958),
            .I(N__41933));
    LocalMux I__7648 (
            .O(N__41955),
            .I(N__41930));
    Span4Mux_v I__7647 (
            .O(N__41952),
            .I(N__41927));
    Span4Mux_h I__7646 (
            .O(N__41949),
            .I(N__41924));
    Sp12to4 I__7645 (
            .O(N__41946),
            .I(N__41916));
    Sp12to4 I__7644 (
            .O(N__41941),
            .I(N__41916));
    LocalMux I__7643 (
            .O(N__41938),
            .I(N__41916));
    LocalMux I__7642 (
            .O(N__41933),
            .I(N__41913));
    Span4Mux_v I__7641 (
            .O(N__41930),
            .I(N__41910));
    Span4Mux_h I__7640 (
            .O(N__41927),
            .I(N__41905));
    Span4Mux_h I__7639 (
            .O(N__41924),
            .I(N__41905));
    InMux I__7638 (
            .O(N__41923),
            .I(N__41902));
    Span12Mux_v I__7637 (
            .O(N__41916),
            .I(N__41899));
    Odrv4 I__7636 (
            .O(N__41913),
            .I(\CONTROL.un1_busState114_2_0_0 ));
    Odrv4 I__7635 (
            .O(N__41910),
            .I(\CONTROL.un1_busState114_2_0_0 ));
    Odrv4 I__7634 (
            .O(N__41905),
            .I(\CONTROL.un1_busState114_2_0_0 ));
    LocalMux I__7633 (
            .O(N__41902),
            .I(\CONTROL.un1_busState114_2_0_0 ));
    Odrv12 I__7632 (
            .O(N__41899),
            .I(\CONTROL.un1_busState114_2_0_0 ));
    CascadeMux I__7631 (
            .O(N__41888),
            .I(\CONTROL.g1_1_cascade_ ));
    CascadeMux I__7630 (
            .O(N__41885),
            .I(N__41882));
    InMux I__7629 (
            .O(N__41882),
            .I(N__41879));
    LocalMux I__7628 (
            .O(N__41879),
            .I(N__41876));
    Span4Mux_v I__7627 (
            .O(N__41876),
            .I(N__41873));
    Span4Mux_h I__7626 (
            .O(N__41873),
            .I(N__41870));
    Span4Mux_h I__7625 (
            .O(N__41870),
            .I(N__41867));
    Odrv4 I__7624 (
            .O(N__41867),
            .I(\CONTROL.addrstackptr_N_7_i ));
    CascadeMux I__7623 (
            .O(N__41864),
            .I(N__41861));
    InMux I__7622 (
            .O(N__41861),
            .I(N__41858));
    LocalMux I__7621 (
            .O(N__41858),
            .I(N__41855));
    Odrv4 I__7620 (
            .O(N__41855),
            .I(\CONTROL.g1_0_0 ));
    InMux I__7619 (
            .O(N__41852),
            .I(N__41849));
    LocalMux I__7618 (
            .O(N__41849),
            .I(\CONTROL.g0_i_m2_1 ));
    InMux I__7617 (
            .O(N__41846),
            .I(N__41843));
    LocalMux I__7616 (
            .O(N__41843),
            .I(N__41840));
    Odrv4 I__7615 (
            .O(N__41840),
            .I(\PROM.ROMDATA.m31 ));
    CascadeMux I__7614 (
            .O(N__41837),
            .I(m125_e_cascade_));
    InMux I__7613 (
            .O(N__41834),
            .I(N__41830));
    InMux I__7612 (
            .O(N__41833),
            .I(N__41827));
    LocalMux I__7611 (
            .O(N__41830),
            .I(N__41824));
    LocalMux I__7610 (
            .O(N__41827),
            .I(\PROM.ROMDATA.N_557_mux ));
    Odrv4 I__7609 (
            .O(N__41824),
            .I(\PROM.ROMDATA.N_557_mux ));
    InMux I__7608 (
            .O(N__41819),
            .I(N__41816));
    LocalMux I__7607 (
            .O(N__41816),
            .I(N__41813));
    Odrv4 I__7606 (
            .O(N__41813),
            .I(\PROM.ROMDATA.m77 ));
    InMux I__7605 (
            .O(N__41810),
            .I(N__41807));
    LocalMux I__7604 (
            .O(N__41807),
            .I(N__41802));
    InMux I__7603 (
            .O(N__41806),
            .I(N__41797));
    InMux I__7602 (
            .O(N__41805),
            .I(N__41797));
    Odrv4 I__7601 (
            .O(N__41802),
            .I(m93_ns));
    LocalMux I__7600 (
            .O(N__41797),
            .I(m93_ns));
    CascadeMux I__7599 (
            .O(N__41792),
            .I(m93_ns_cascade_));
    InMux I__7598 (
            .O(N__41789),
            .I(N__41786));
    LocalMux I__7597 (
            .O(N__41786),
            .I(N__41783));
    Span4Mux_v I__7596 (
            .O(N__41783),
            .I(N__41780));
    Span4Mux_h I__7595 (
            .O(N__41780),
            .I(N__41777));
    Span4Mux_h I__7594 (
            .O(N__41777),
            .I(N__41774));
    Odrv4 I__7593 (
            .O(N__41774),
            .I(\CONTROL.addrstack_5 ));
    InMux I__7592 (
            .O(N__41771),
            .I(N__41768));
    LocalMux I__7591 (
            .O(N__41768),
            .I(N__41765));
    Span4Mux_h I__7590 (
            .O(N__41765),
            .I(N__41760));
    InMux I__7589 (
            .O(N__41764),
            .I(N__41757));
    InMux I__7588 (
            .O(N__41763),
            .I(N__41754));
    Odrv4 I__7587 (
            .O(N__41760),
            .I(\CONTROL.addrstack_reto_5 ));
    LocalMux I__7586 (
            .O(N__41757),
            .I(\CONTROL.addrstack_reto_5 ));
    LocalMux I__7585 (
            .O(N__41754),
            .I(\CONTROL.addrstack_reto_5 ));
    InMux I__7584 (
            .O(N__41747),
            .I(N__41744));
    LocalMux I__7583 (
            .O(N__41744),
            .I(N__41741));
    Span4Mux_v I__7582 (
            .O(N__41741),
            .I(N__41737));
    InMux I__7581 (
            .O(N__41740),
            .I(N__41734));
    Span4Mux_h I__7580 (
            .O(N__41737),
            .I(N__41729));
    LocalMux I__7579 (
            .O(N__41734),
            .I(N__41729));
    Span4Mux_h I__7578 (
            .O(N__41729),
            .I(N__41726));
    Odrv4 I__7577 (
            .O(N__41726),
            .I(\CONTROL.programCounter_1_5 ));
    InMux I__7576 (
            .O(N__41723),
            .I(N__41720));
    LocalMux I__7575 (
            .O(N__41720),
            .I(N__41717));
    Span4Mux_h I__7574 (
            .O(N__41717),
            .I(N__41713));
    InMux I__7573 (
            .O(N__41716),
            .I(N__41710));
    Odrv4 I__7572 (
            .O(N__41713),
            .I(\CONTROL.programCounter_1_reto_5 ));
    LocalMux I__7571 (
            .O(N__41710),
            .I(\CONTROL.programCounter_1_reto_5 ));
    CascadeMux I__7570 (
            .O(N__41705),
            .I(\CONTROL.N_86_0_cascade_ ));
    CascadeMux I__7569 (
            .O(N__41702),
            .I(N__41699));
    InMux I__7568 (
            .O(N__41699),
            .I(N__41693));
    CascadeMux I__7567 (
            .O(N__41698),
            .I(N__41690));
    InMux I__7566 (
            .O(N__41697),
            .I(N__41685));
    CascadeMux I__7565 (
            .O(N__41696),
            .I(N__41682));
    LocalMux I__7564 (
            .O(N__41693),
            .I(N__41679));
    InMux I__7563 (
            .O(N__41690),
            .I(N__41676));
    InMux I__7562 (
            .O(N__41689),
            .I(N__41671));
    InMux I__7561 (
            .O(N__41688),
            .I(N__41671));
    LocalMux I__7560 (
            .O(N__41685),
            .I(N__41667));
    InMux I__7559 (
            .O(N__41682),
            .I(N__41664));
    Span4Mux_v I__7558 (
            .O(N__41679),
            .I(N__41659));
    LocalMux I__7557 (
            .O(N__41676),
            .I(N__41659));
    LocalMux I__7556 (
            .O(N__41671),
            .I(N__41656));
    CascadeMux I__7555 (
            .O(N__41670),
            .I(N__41652));
    Span4Mux_v I__7554 (
            .O(N__41667),
            .I(N__41647));
    LocalMux I__7553 (
            .O(N__41664),
            .I(N__41642));
    Span4Mux_h I__7552 (
            .O(N__41659),
            .I(N__41642));
    Span4Mux_h I__7551 (
            .O(N__41656),
            .I(N__41639));
    InMux I__7550 (
            .O(N__41655),
            .I(N__41636));
    InMux I__7549 (
            .O(N__41652),
            .I(N__41633));
    InMux I__7548 (
            .O(N__41651),
            .I(N__41628));
    InMux I__7547 (
            .O(N__41650),
            .I(N__41628));
    Odrv4 I__7546 (
            .O(N__41647),
            .I(controlWord_1));
    Odrv4 I__7545 (
            .O(N__41642),
            .I(controlWord_1));
    Odrv4 I__7544 (
            .O(N__41639),
            .I(controlWord_1));
    LocalMux I__7543 (
            .O(N__41636),
            .I(controlWord_1));
    LocalMux I__7542 (
            .O(N__41633),
            .I(controlWord_1));
    LocalMux I__7541 (
            .O(N__41628),
            .I(controlWord_1));
    InMux I__7540 (
            .O(N__41615),
            .I(N__41612));
    LocalMux I__7539 (
            .O(N__41612),
            .I(N__41609));
    Span4Mux_h I__7538 (
            .O(N__41609),
            .I(N__41606));
    Odrv4 I__7537 (
            .O(N__41606),
            .I(\CONTROL.N_135 ));
    InMux I__7536 (
            .O(N__41603),
            .I(N__41597));
    InMux I__7535 (
            .O(N__41602),
            .I(N__41597));
    LocalMux I__7534 (
            .O(N__41597),
            .I(N__41591));
    InMux I__7533 (
            .O(N__41596),
            .I(N__41586));
    InMux I__7532 (
            .O(N__41595),
            .I(N__41586));
    InMux I__7531 (
            .O(N__41594),
            .I(N__41583));
    Span4Mux_v I__7530 (
            .O(N__41591),
            .I(N__41577));
    LocalMux I__7529 (
            .O(N__41586),
            .I(N__41572));
    LocalMux I__7528 (
            .O(N__41583),
            .I(N__41569));
    InMux I__7527 (
            .O(N__41582),
            .I(N__41566));
    InMux I__7526 (
            .O(N__41581),
            .I(N__41563));
    InMux I__7525 (
            .O(N__41580),
            .I(N__41560));
    Span4Mux_h I__7524 (
            .O(N__41577),
            .I(N__41555));
    InMux I__7523 (
            .O(N__41576),
            .I(N__41550));
    InMux I__7522 (
            .O(N__41575),
            .I(N__41550));
    Span4Mux_h I__7521 (
            .O(N__41572),
            .I(N__41545));
    Span4Mux_h I__7520 (
            .O(N__41569),
            .I(N__41545));
    LocalMux I__7519 (
            .O(N__41566),
            .I(N__41542));
    LocalMux I__7518 (
            .O(N__41563),
            .I(N__41539));
    LocalMux I__7517 (
            .O(N__41560),
            .I(N__41536));
    InMux I__7516 (
            .O(N__41559),
            .I(N__41531));
    InMux I__7515 (
            .O(N__41558),
            .I(N__41531));
    Span4Mux_h I__7514 (
            .O(N__41555),
            .I(N__41526));
    LocalMux I__7513 (
            .O(N__41550),
            .I(N__41526));
    Span4Mux_h I__7512 (
            .O(N__41545),
            .I(N__41523));
    Span4Mux_h I__7511 (
            .O(N__41542),
            .I(N__41518));
    Span4Mux_h I__7510 (
            .O(N__41539),
            .I(N__41518));
    Span12Mux_h I__7509 (
            .O(N__41536),
            .I(N__41515));
    LocalMux I__7508 (
            .O(N__41531),
            .I(\CONTROL.N_74_0 ));
    Odrv4 I__7507 (
            .O(N__41526),
            .I(\CONTROL.N_74_0 ));
    Odrv4 I__7506 (
            .O(N__41523),
            .I(\CONTROL.N_74_0 ));
    Odrv4 I__7505 (
            .O(N__41518),
            .I(\CONTROL.N_74_0 ));
    Odrv12 I__7504 (
            .O(N__41515),
            .I(\CONTROL.N_74_0 ));
    InMux I__7503 (
            .O(N__41504),
            .I(N__41500));
    InMux I__7502 (
            .O(N__41503),
            .I(N__41497));
    LocalMux I__7501 (
            .O(N__41500),
            .I(N__41493));
    LocalMux I__7500 (
            .O(N__41497),
            .I(N__41490));
    InMux I__7499 (
            .O(N__41496),
            .I(N__41485));
    Span4Mux_v I__7498 (
            .O(N__41493),
            .I(N__41480));
    Span4Mux_v I__7497 (
            .O(N__41490),
            .I(N__41480));
    InMux I__7496 (
            .O(N__41489),
            .I(N__41477));
    InMux I__7495 (
            .O(N__41488),
            .I(N__41473));
    LocalMux I__7494 (
            .O(N__41485),
            .I(N__41470));
    Span4Mux_h I__7493 (
            .O(N__41480),
            .I(N__41465));
    LocalMux I__7492 (
            .O(N__41477),
            .I(N__41465));
    InMux I__7491 (
            .O(N__41476),
            .I(N__41460));
    LocalMux I__7490 (
            .O(N__41473),
            .I(N__41457));
    Span4Mux_h I__7489 (
            .O(N__41470),
            .I(N__41452));
    Span4Mux_h I__7488 (
            .O(N__41465),
            .I(N__41452));
    InMux I__7487 (
            .O(N__41464),
            .I(N__41449));
    InMux I__7486 (
            .O(N__41463),
            .I(N__41446));
    LocalMux I__7485 (
            .O(N__41460),
            .I(\CONTROL.N_249 ));
    Odrv12 I__7484 (
            .O(N__41457),
            .I(\CONTROL.N_249 ));
    Odrv4 I__7483 (
            .O(N__41452),
            .I(\CONTROL.N_249 ));
    LocalMux I__7482 (
            .O(N__41449),
            .I(\CONTROL.N_249 ));
    LocalMux I__7481 (
            .O(N__41446),
            .I(\CONTROL.N_249 ));
    CascadeMux I__7480 (
            .O(N__41435),
            .I(N__41425));
    InMux I__7479 (
            .O(N__41434),
            .I(N__41420));
    CascadeMux I__7478 (
            .O(N__41433),
            .I(N__41417));
    InMux I__7477 (
            .O(N__41432),
            .I(N__41412));
    InMux I__7476 (
            .O(N__41431),
            .I(N__41409));
    InMux I__7475 (
            .O(N__41430),
            .I(N__41405));
    InMux I__7474 (
            .O(N__41429),
            .I(N__41398));
    InMux I__7473 (
            .O(N__41428),
            .I(N__41398));
    InMux I__7472 (
            .O(N__41425),
            .I(N__41398));
    InMux I__7471 (
            .O(N__41424),
            .I(N__41388));
    InMux I__7470 (
            .O(N__41423),
            .I(N__41385));
    LocalMux I__7469 (
            .O(N__41420),
            .I(N__41382));
    InMux I__7468 (
            .O(N__41417),
            .I(N__41379));
    CascadeMux I__7467 (
            .O(N__41416),
            .I(N__41376));
    CascadeMux I__7466 (
            .O(N__41415),
            .I(N__41373));
    LocalMux I__7465 (
            .O(N__41412),
            .I(N__41366));
    LocalMux I__7464 (
            .O(N__41409),
            .I(N__41366));
    InMux I__7463 (
            .O(N__41408),
            .I(N__41363));
    LocalMux I__7462 (
            .O(N__41405),
            .I(N__41358));
    LocalMux I__7461 (
            .O(N__41398),
            .I(N__41358));
    CascadeMux I__7460 (
            .O(N__41397),
            .I(N__41353));
    InMux I__7459 (
            .O(N__41396),
            .I(N__41350));
    CascadeMux I__7458 (
            .O(N__41395),
            .I(N__41347));
    InMux I__7457 (
            .O(N__41394),
            .I(N__41340));
    InMux I__7456 (
            .O(N__41393),
            .I(N__41340));
    InMux I__7455 (
            .O(N__41392),
            .I(N__41340));
    InMux I__7454 (
            .O(N__41391),
            .I(N__41337));
    LocalMux I__7453 (
            .O(N__41388),
            .I(N__41328));
    LocalMux I__7452 (
            .O(N__41385),
            .I(N__41328));
    Span4Mux_v I__7451 (
            .O(N__41382),
            .I(N__41328));
    LocalMux I__7450 (
            .O(N__41379),
            .I(N__41328));
    InMux I__7449 (
            .O(N__41376),
            .I(N__41319));
    InMux I__7448 (
            .O(N__41373),
            .I(N__41319));
    InMux I__7447 (
            .O(N__41372),
            .I(N__41319));
    InMux I__7446 (
            .O(N__41371),
            .I(N__41319));
    Span4Mux_h I__7445 (
            .O(N__41366),
            .I(N__41312));
    LocalMux I__7444 (
            .O(N__41363),
            .I(N__41312));
    Span4Mux_v I__7443 (
            .O(N__41358),
            .I(N__41312));
    CascadeMux I__7442 (
            .O(N__41357),
            .I(N__41309));
    CascadeMux I__7441 (
            .O(N__41356),
            .I(N__41306));
    InMux I__7440 (
            .O(N__41353),
            .I(N__41302));
    LocalMux I__7439 (
            .O(N__41350),
            .I(N__41299));
    InMux I__7438 (
            .O(N__41347),
            .I(N__41296));
    LocalMux I__7437 (
            .O(N__41340),
            .I(N__41289));
    LocalMux I__7436 (
            .O(N__41337),
            .I(N__41289));
    Span4Mux_v I__7435 (
            .O(N__41328),
            .I(N__41289));
    LocalMux I__7434 (
            .O(N__41319),
            .I(N__41284));
    Span4Mux_h I__7433 (
            .O(N__41312),
            .I(N__41284));
    InMux I__7432 (
            .O(N__41309),
            .I(N__41277));
    InMux I__7431 (
            .O(N__41306),
            .I(N__41277));
    InMux I__7430 (
            .O(N__41305),
            .I(N__41277));
    LocalMux I__7429 (
            .O(N__41302),
            .I(controlWord_5));
    Odrv4 I__7428 (
            .O(N__41299),
            .I(controlWord_5));
    LocalMux I__7427 (
            .O(N__41296),
            .I(controlWord_5));
    Odrv4 I__7426 (
            .O(N__41289),
            .I(controlWord_5));
    Odrv4 I__7425 (
            .O(N__41284),
            .I(controlWord_5));
    LocalMux I__7424 (
            .O(N__41277),
            .I(controlWord_5));
    CascadeMux I__7423 (
            .O(N__41264),
            .I(\CONTROL.N_74_0_cascade_ ));
    CascadeMux I__7422 (
            .O(N__41261),
            .I(N__41253));
    InMux I__7421 (
            .O(N__41260),
            .I(N__41250));
    CascadeMux I__7420 (
            .O(N__41259),
            .I(N__41242));
    InMux I__7419 (
            .O(N__41258),
            .I(N__41236));
    InMux I__7418 (
            .O(N__41257),
            .I(N__41236));
    InMux I__7417 (
            .O(N__41256),
            .I(N__41230));
    InMux I__7416 (
            .O(N__41253),
            .I(N__41227));
    LocalMux I__7415 (
            .O(N__41250),
            .I(N__41224));
    InMux I__7414 (
            .O(N__41249),
            .I(N__41211));
    InMux I__7413 (
            .O(N__41248),
            .I(N__41211));
    InMux I__7412 (
            .O(N__41247),
            .I(N__41211));
    InMux I__7411 (
            .O(N__41246),
            .I(N__41211));
    InMux I__7410 (
            .O(N__41245),
            .I(N__41211));
    InMux I__7409 (
            .O(N__41242),
            .I(N__41211));
    InMux I__7408 (
            .O(N__41241),
            .I(N__41207));
    LocalMux I__7407 (
            .O(N__41236),
            .I(N__41204));
    CascadeMux I__7406 (
            .O(N__41235),
            .I(N__41198));
    InMux I__7405 (
            .O(N__41234),
            .I(N__41195));
    InMux I__7404 (
            .O(N__41233),
            .I(N__41188));
    LocalMux I__7403 (
            .O(N__41230),
            .I(N__41185));
    LocalMux I__7402 (
            .O(N__41227),
            .I(N__41182));
    Span4Mux_h I__7401 (
            .O(N__41224),
            .I(N__41177));
    LocalMux I__7400 (
            .O(N__41211),
            .I(N__41177));
    InMux I__7399 (
            .O(N__41210),
            .I(N__41174));
    LocalMux I__7398 (
            .O(N__41207),
            .I(N__41171));
    Span4Mux_h I__7397 (
            .O(N__41204),
            .I(N__41168));
    InMux I__7396 (
            .O(N__41203),
            .I(N__41163));
    InMux I__7395 (
            .O(N__41202),
            .I(N__41163));
    InMux I__7394 (
            .O(N__41201),
            .I(N__41158));
    InMux I__7393 (
            .O(N__41198),
            .I(N__41158));
    LocalMux I__7392 (
            .O(N__41195),
            .I(N__41155));
    InMux I__7391 (
            .O(N__41194),
            .I(N__41146));
    InMux I__7390 (
            .O(N__41193),
            .I(N__41146));
    InMux I__7389 (
            .O(N__41192),
            .I(N__41146));
    InMux I__7388 (
            .O(N__41191),
            .I(N__41146));
    LocalMux I__7387 (
            .O(N__41188),
            .I(N__41137));
    Span4Mux_v I__7386 (
            .O(N__41185),
            .I(N__41137));
    Span4Mux_h I__7385 (
            .O(N__41182),
            .I(N__41137));
    Span4Mux_h I__7384 (
            .O(N__41177),
            .I(N__41137));
    LocalMux I__7383 (
            .O(N__41174),
            .I(controlWord_6));
    Odrv12 I__7382 (
            .O(N__41171),
            .I(controlWord_6));
    Odrv4 I__7381 (
            .O(N__41168),
            .I(controlWord_6));
    LocalMux I__7380 (
            .O(N__41163),
            .I(controlWord_6));
    LocalMux I__7379 (
            .O(N__41158),
            .I(controlWord_6));
    Odrv4 I__7378 (
            .O(N__41155),
            .I(controlWord_6));
    LocalMux I__7377 (
            .O(N__41146),
            .I(controlWord_6));
    Odrv4 I__7376 (
            .O(N__41137),
            .I(controlWord_6));
    CascadeMux I__7375 (
            .O(N__41120),
            .I(\CONTROL.un1_busState96_1_i_i_232_1_cascade_ ));
    InMux I__7374 (
            .O(N__41117),
            .I(N__41114));
    LocalMux I__7373 (
            .O(N__41114),
            .I(\CONTROL.programCounter_ret_36_RNINU4NARZ0Z_7 ));
    CascadeMux I__7372 (
            .O(N__41111),
            .I(\PROM.ROMDATA.m23_cascade_ ));
    InMux I__7371 (
            .O(N__41108),
            .I(N__41105));
    LocalMux I__7370 (
            .O(N__41105),
            .I(N__41102));
    Span4Mux_v I__7369 (
            .O(N__41102),
            .I(N__41097));
    InMux I__7368 (
            .O(N__41101),
            .I(N__41092));
    InMux I__7367 (
            .O(N__41100),
            .I(N__41092));
    Span4Mux_h I__7366 (
            .O(N__41097),
            .I(N__41089));
    LocalMux I__7365 (
            .O(N__41092),
            .I(N__41086));
    Odrv4 I__7364 (
            .O(N__41089),
            .I(PROM_ROMDATA_dintern_31_0__N_556_mux));
    Odrv4 I__7363 (
            .O(N__41086),
            .I(PROM_ROMDATA_dintern_31_0__N_556_mux));
    InMux I__7362 (
            .O(N__41081),
            .I(N__41078));
    LocalMux I__7361 (
            .O(N__41078),
            .I(N__41075));
    Odrv4 I__7360 (
            .O(N__41075),
            .I(\PROM.ROMDATA.m294_am ));
    CascadeMux I__7359 (
            .O(N__41072),
            .I(N__41069));
    InMux I__7358 (
            .O(N__41069),
            .I(N__41066));
    LocalMux I__7357 (
            .O(N__41066),
            .I(N__41063));
    Span4Mux_h I__7356 (
            .O(N__41063),
            .I(N__41060));
    Odrv4 I__7355 (
            .O(N__41060),
            .I(\PROM.ROMDATA.m271_1 ));
    CascadeMux I__7354 (
            .O(N__41057),
            .I(\PROM.ROMDATA.m271_1_cascade_ ));
    InMux I__7353 (
            .O(N__41054),
            .I(N__41046));
    InMux I__7352 (
            .O(N__41053),
            .I(N__41046));
    InMux I__7351 (
            .O(N__41052),
            .I(N__41041));
    InMux I__7350 (
            .O(N__41051),
            .I(N__41041));
    LocalMux I__7349 (
            .O(N__41046),
            .I(N__41036));
    LocalMux I__7348 (
            .O(N__41041),
            .I(N__41036));
    Span4Mux_v I__7347 (
            .O(N__41036),
            .I(N__41033));
    Span4Mux_v I__7346 (
            .O(N__41033),
            .I(N__41030));
    Span4Mux_h I__7345 (
            .O(N__41030),
            .I(N__41027));
    Odrv4 I__7344 (
            .O(N__41027),
            .I(\PROM.ROMDATA.m258_ns ));
    CascadeMux I__7343 (
            .O(N__41024),
            .I(\PROM.ROMDATA.m258_ns_cascade_ ));
    CascadeMux I__7342 (
            .O(N__41021),
            .I(PROM_ROMDATA_dintern_9ro_cascade_));
    InMux I__7341 (
            .O(N__41018),
            .I(N__41015));
    LocalMux I__7340 (
            .O(N__41015),
            .I(\CONTROL.increment28lto5_1Z0Z_0 ));
    CascadeMux I__7339 (
            .O(N__41012),
            .I(N__41009));
    InMux I__7338 (
            .O(N__41009),
            .I(N__41005));
    InMux I__7337 (
            .O(N__41008),
            .I(N__41002));
    LocalMux I__7336 (
            .O(N__41005),
            .I(N__40999));
    LocalMux I__7335 (
            .O(N__41002),
            .I(N__40996));
    Span4Mux_v I__7334 (
            .O(N__40999),
            .I(N__40993));
    Span4Mux_v I__7333 (
            .O(N__40996),
            .I(N__40988));
    Span4Mux_h I__7332 (
            .O(N__40993),
            .I(N__40988));
    Odrv4 I__7331 (
            .O(N__40988),
            .I(\PROM.ROMDATA.N_566_mux ));
    InMux I__7330 (
            .O(N__40985),
            .I(N__40982));
    LocalMux I__7329 (
            .O(N__40982),
            .I(N__40979));
    Span4Mux_v I__7328 (
            .O(N__40979),
            .I(N__40976));
    Span4Mux_h I__7327 (
            .O(N__40976),
            .I(N__40973));
    Span4Mux_h I__7326 (
            .O(N__40973),
            .I(N__40970));
    Odrv4 I__7325 (
            .O(N__40970),
            .I(\PROM.ROMDATA.m470_bm ));
    CascadeMux I__7324 (
            .O(N__40967),
            .I(N__40964));
    InMux I__7323 (
            .O(N__40964),
            .I(N__40959));
    InMux I__7322 (
            .O(N__40963),
            .I(N__40955));
    CascadeMux I__7321 (
            .O(N__40962),
            .I(N__40952));
    LocalMux I__7320 (
            .O(N__40959),
            .I(N__40949));
    InMux I__7319 (
            .O(N__40958),
            .I(N__40946));
    LocalMux I__7318 (
            .O(N__40955),
            .I(N__40943));
    InMux I__7317 (
            .O(N__40952),
            .I(N__40940));
    Span12Mux_h I__7316 (
            .O(N__40949),
            .I(N__40935));
    LocalMux I__7315 (
            .O(N__40946),
            .I(N__40935));
    Span4Mux_v I__7314 (
            .O(N__40943),
            .I(N__40930));
    LocalMux I__7313 (
            .O(N__40940),
            .I(N__40930));
    Odrv12 I__7312 (
            .O(N__40935),
            .I(\CONTROL.N_215 ));
    Odrv4 I__7311 (
            .O(N__40930),
            .I(\CONTROL.N_215 ));
    CascadeMux I__7310 (
            .O(N__40925),
            .I(N__40921));
    CascadeMux I__7309 (
            .O(N__40924),
            .I(N__40917));
    InMux I__7308 (
            .O(N__40921),
            .I(N__40906));
    InMux I__7307 (
            .O(N__40920),
            .I(N__40906));
    InMux I__7306 (
            .O(N__40917),
            .I(N__40901));
    InMux I__7305 (
            .O(N__40916),
            .I(N__40901));
    InMux I__7304 (
            .O(N__40915),
            .I(N__40896));
    InMux I__7303 (
            .O(N__40914),
            .I(N__40896));
    InMux I__7302 (
            .O(N__40913),
            .I(N__40893));
    InMux I__7301 (
            .O(N__40912),
            .I(N__40884));
    InMux I__7300 (
            .O(N__40911),
            .I(N__40884));
    LocalMux I__7299 (
            .O(N__40906),
            .I(N__40881));
    LocalMux I__7298 (
            .O(N__40901),
            .I(N__40878));
    LocalMux I__7297 (
            .O(N__40896),
            .I(N__40875));
    LocalMux I__7296 (
            .O(N__40893),
            .I(N__40872));
    InMux I__7295 (
            .O(N__40892),
            .I(N__40863));
    InMux I__7294 (
            .O(N__40891),
            .I(N__40863));
    InMux I__7293 (
            .O(N__40890),
            .I(N__40863));
    InMux I__7292 (
            .O(N__40889),
            .I(N__40863));
    LocalMux I__7291 (
            .O(N__40884),
            .I(N__40860));
    Span4Mux_v I__7290 (
            .O(N__40881),
            .I(N__40857));
    Span4Mux_v I__7289 (
            .O(N__40878),
            .I(N__40850));
    Span4Mux_v I__7288 (
            .O(N__40875),
            .I(N__40850));
    Span4Mux_v I__7287 (
            .O(N__40872),
            .I(N__40850));
    LocalMux I__7286 (
            .O(N__40863),
            .I(N__40847));
    Span4Mux_h I__7285 (
            .O(N__40860),
            .I(N__40844));
    Sp12to4 I__7284 (
            .O(N__40857),
            .I(N__40839));
    Sp12to4 I__7283 (
            .O(N__40850),
            .I(N__40839));
    Odrv4 I__7282 (
            .O(N__40847),
            .I(\PROM.ROMDATA.dintern_12dfltZ0Z_0 ));
    Odrv4 I__7281 (
            .O(N__40844),
            .I(\PROM.ROMDATA.dintern_12dfltZ0Z_0 ));
    Odrv12 I__7280 (
            .O(N__40839),
            .I(\PROM.ROMDATA.dintern_12dfltZ0Z_0 ));
    CascadeMux I__7279 (
            .O(N__40832),
            .I(\PROM.ROMDATA.m284_cascade_ ));
    CascadeMux I__7278 (
            .O(N__40829),
            .I(controlWord_12_cascade_));
    InMux I__7277 (
            .O(N__40826),
            .I(N__40823));
    LocalMux I__7276 (
            .O(N__40823),
            .I(N__40820));
    Span4Mux_h I__7275 (
            .O(N__40820),
            .I(N__40815));
    InMux I__7274 (
            .O(N__40819),
            .I(N__40812));
    InMux I__7273 (
            .O(N__40818),
            .I(N__40809));
    Odrv4 I__7272 (
            .O(N__40815),
            .I(\CONTROL.increment28lto5_0 ));
    LocalMux I__7271 (
            .O(N__40812),
            .I(\CONTROL.increment28lto5_0 ));
    LocalMux I__7270 (
            .O(N__40809),
            .I(\CONTROL.increment28lto5_0 ));
    CascadeMux I__7269 (
            .O(N__40802),
            .I(N__40797));
    InMux I__7268 (
            .O(N__40801),
            .I(N__40787));
    InMux I__7267 (
            .O(N__40800),
            .I(N__40787));
    InMux I__7266 (
            .O(N__40797),
            .I(N__40787));
    InMux I__7265 (
            .O(N__40796),
            .I(N__40787));
    LocalMux I__7264 (
            .O(N__40787),
            .I(N__40784));
    Odrv12 I__7263 (
            .O(N__40784),
            .I(\PROM.ROMDATA.m273 ));
    CascadeMux I__7262 (
            .O(N__40781),
            .I(\PROM.ROMDATA.m273_cascade_ ));
    CascadeMux I__7261 (
            .O(N__40778),
            .I(PROM_ROMDATA_dintern_11ro_cascade_));
    InMux I__7260 (
            .O(N__40775),
            .I(N__40772));
    LocalMux I__7259 (
            .O(N__40772),
            .I(\CONTROL.increment28lto5_0_xZ0Z1 ));
    InMux I__7258 (
            .O(N__40769),
            .I(N__40766));
    LocalMux I__7257 (
            .O(N__40766),
            .I(\CONTROL.increment28lto5_0_xZ0Z0 ));
    InMux I__7256 (
            .O(N__40763),
            .I(N__40757));
    InMux I__7255 (
            .O(N__40762),
            .I(N__40757));
    LocalMux I__7254 (
            .O(N__40757),
            .I(PROM_ROMDATA_dintern_11ro));
    CascadeMux I__7253 (
            .O(N__40754),
            .I(N__40751));
    InMux I__7252 (
            .O(N__40751),
            .I(N__40746));
    InMux I__7251 (
            .O(N__40750),
            .I(N__40741));
    InMux I__7250 (
            .O(N__40749),
            .I(N__40741));
    LocalMux I__7249 (
            .O(N__40746),
            .I(N__40736));
    LocalMux I__7248 (
            .O(N__40741),
            .I(N__40736));
    Span4Mux_h I__7247 (
            .O(N__40736),
            .I(N__40733));
    Span4Mux_h I__7246 (
            .O(N__40733),
            .I(N__40730));
    Span4Mux_h I__7245 (
            .O(N__40730),
            .I(N__40726));
    InMux I__7244 (
            .O(N__40729),
            .I(N__40723));
    Span4Mux_v I__7243 (
            .O(N__40726),
            .I(N__40720));
    LocalMux I__7242 (
            .O(N__40723),
            .I(aluStatus_4));
    Odrv4 I__7241 (
            .O(N__40720),
            .I(aluStatus_4));
    InMux I__7240 (
            .O(N__40715),
            .I(N__40712));
    LocalMux I__7239 (
            .O(N__40712),
            .I(controlWord_12));
    InMux I__7238 (
            .O(N__40709),
            .I(N__40706));
    LocalMux I__7237 (
            .O(N__40706),
            .I(N__40703));
    Span4Mux_h I__7236 (
            .O(N__40703),
            .I(N__40700));
    Sp12to4 I__7235 (
            .O(N__40700),
            .I(N__40697));
    Span12Mux_v I__7234 (
            .O(N__40697),
            .I(N__40694));
    Odrv12 I__7233 (
            .O(N__40694),
            .I(\CONTROL.g0_1_i_a6Z0Z_0 ));
    InMux I__7232 (
            .O(N__40691),
            .I(N__40688));
    LocalMux I__7231 (
            .O(N__40688),
            .I(N__40685));
    Span4Mux_h I__7230 (
            .O(N__40685),
            .I(N__40682));
    Span4Mux_v I__7229 (
            .O(N__40682),
            .I(N__40679));
    Odrv4 I__7228 (
            .O(N__40679),
            .I(\CONTROL.g0_1_i_a6Z0Z_1 ));
    InMux I__7227 (
            .O(N__40676),
            .I(N__40673));
    LocalMux I__7226 (
            .O(N__40673),
            .I(N__40670));
    Span4Mux_v I__7225 (
            .O(N__40670),
            .I(N__40667));
    Span4Mux_h I__7224 (
            .O(N__40667),
            .I(N__40664));
    Span4Mux_h I__7223 (
            .O(N__40664),
            .I(N__40661));
    Odrv4 I__7222 (
            .O(N__40661),
            .I(\CONTROL.g0_3_i_a7Z0Z_0 ));
    CEMux I__7221 (
            .O(N__40658),
            .I(N__40654));
    CEMux I__7220 (
            .O(N__40657),
            .I(N__40651));
    LocalMux I__7219 (
            .O(N__40654),
            .I(N__40648));
    LocalMux I__7218 (
            .O(N__40651),
            .I(N__40644));
    Span4Mux_v I__7217 (
            .O(N__40648),
            .I(N__40641));
    CEMux I__7216 (
            .O(N__40647),
            .I(N__40638));
    Span4Mux_v I__7215 (
            .O(N__40644),
            .I(N__40629));
    Span4Mux_h I__7214 (
            .O(N__40641),
            .I(N__40629));
    LocalMux I__7213 (
            .O(N__40638),
            .I(N__40629));
    InMux I__7212 (
            .O(N__40637),
            .I(N__40626));
    InMux I__7211 (
            .O(N__40636),
            .I(N__40622));
    Span4Mux_h I__7210 (
            .O(N__40629),
            .I(N__40619));
    LocalMux I__7209 (
            .O(N__40626),
            .I(N__40616));
    InMux I__7208 (
            .O(N__40625),
            .I(N__40613));
    LocalMux I__7207 (
            .O(N__40622),
            .I(N__40610));
    Odrv4 I__7206 (
            .O(N__40619),
            .I(\CONTROL.aluReadBus_1_sqmuxa ));
    Odrv4 I__7205 (
            .O(N__40616),
            .I(\CONTROL.aluReadBus_1_sqmuxa ));
    LocalMux I__7204 (
            .O(N__40613),
            .I(\CONTROL.aluReadBus_1_sqmuxa ));
    Odrv4 I__7203 (
            .O(N__40610),
            .I(\CONTROL.aluReadBus_1_sqmuxa ));
    InMux I__7202 (
            .O(N__40601),
            .I(N__40598));
    LocalMux I__7201 (
            .O(N__40598),
            .I(N__40595));
    Span4Mux_v I__7200 (
            .O(N__40595),
            .I(N__40589));
    InMux I__7199 (
            .O(N__40594),
            .I(N__40586));
    InMux I__7198 (
            .O(N__40593),
            .I(N__40582));
    CascadeMux I__7197 (
            .O(N__40592),
            .I(N__40577));
    Span4Mux_h I__7196 (
            .O(N__40589),
            .I(N__40571));
    LocalMux I__7195 (
            .O(N__40586),
            .I(N__40571));
    InMux I__7194 (
            .O(N__40585),
            .I(N__40568));
    LocalMux I__7193 (
            .O(N__40582),
            .I(N__40565));
    InMux I__7192 (
            .O(N__40581),
            .I(N__40560));
    InMux I__7191 (
            .O(N__40580),
            .I(N__40560));
    InMux I__7190 (
            .O(N__40577),
            .I(N__40555));
    InMux I__7189 (
            .O(N__40576),
            .I(N__40555));
    Span4Mux_h I__7188 (
            .O(N__40571),
            .I(N__40550));
    LocalMux I__7187 (
            .O(N__40568),
            .I(N__40550));
    Odrv4 I__7186 (
            .O(N__40565),
            .I(\ALU.un14_log_a0_2Z0Z_15 ));
    LocalMux I__7185 (
            .O(N__40560),
            .I(\ALU.un14_log_a0_2Z0Z_15 ));
    LocalMux I__7184 (
            .O(N__40555),
            .I(\ALU.un14_log_a0_2Z0Z_15 ));
    Odrv4 I__7183 (
            .O(N__40550),
            .I(\ALU.un14_log_a0_2Z0Z_15 ));
    InMux I__7182 (
            .O(N__40541),
            .I(N__40537));
    InMux I__7181 (
            .O(N__40540),
            .I(N__40534));
    LocalMux I__7180 (
            .O(N__40537),
            .I(N__40531));
    LocalMux I__7179 (
            .O(N__40534),
            .I(N__40528));
    Span4Mux_v I__7178 (
            .O(N__40531),
            .I(N__40523));
    Span4Mux_h I__7177 (
            .O(N__40528),
            .I(N__40523));
    Odrv4 I__7176 (
            .O(N__40523),
            .I(\ALU.d_RNIN8NU4Z0Z_9 ));
    InMux I__7175 (
            .O(N__40520),
            .I(N__40517));
    LocalMux I__7174 (
            .O(N__40517),
            .I(N__40514));
    Span4Mux_v I__7173 (
            .O(N__40514),
            .I(N__40510));
    InMux I__7172 (
            .O(N__40513),
            .I(N__40507));
    Span4Mux_h I__7171 (
            .O(N__40510),
            .I(N__40504));
    LocalMux I__7170 (
            .O(N__40507),
            .I(\ALU.combOperand2_0_0_9 ));
    Odrv4 I__7169 (
            .O(N__40504),
            .I(\ALU.combOperand2_0_0_9 ));
    CascadeMux I__7168 (
            .O(N__40499),
            .I(N__40495));
    InMux I__7167 (
            .O(N__40498),
            .I(N__40491));
    InMux I__7166 (
            .O(N__40495),
            .I(N__40488));
    CascadeMux I__7165 (
            .O(N__40494),
            .I(N__40485));
    LocalMux I__7164 (
            .O(N__40491),
            .I(N__40480));
    LocalMux I__7163 (
            .O(N__40488),
            .I(N__40480));
    InMux I__7162 (
            .O(N__40485),
            .I(N__40477));
    Span4Mux_h I__7161 (
            .O(N__40480),
            .I(N__40474));
    LocalMux I__7160 (
            .O(N__40477),
            .I(N__40471));
    Span4Mux_h I__7159 (
            .O(N__40474),
            .I(N__40466));
    Span4Mux_v I__7158 (
            .O(N__40471),
            .I(N__40466));
    Odrv4 I__7157 (
            .O(N__40466),
            .I(DROM_ROMDATA_dintern_9ro));
    InMux I__7156 (
            .O(N__40463),
            .I(N__40460));
    LocalMux I__7155 (
            .O(N__40460),
            .I(N__40457));
    Span4Mux_h I__7154 (
            .O(N__40457),
            .I(N__40454));
    Span4Mux_v I__7153 (
            .O(N__40454),
            .I(N__40451));
    Span4Mux_v I__7152 (
            .O(N__40451),
            .I(N__40448));
    Span4Mux_v I__7151 (
            .O(N__40448),
            .I(N__40445));
    Span4Mux_h I__7150 (
            .O(N__40445),
            .I(N__40442));
    Span4Mux_h I__7149 (
            .O(N__40442),
            .I(N__40439));
    Span4Mux_h I__7148 (
            .O(N__40439),
            .I(N__40436));
    Odrv4 I__7147 (
            .O(N__40436),
            .I(gpuOut_c_9));
    InMux I__7146 (
            .O(N__40433),
            .I(N__40430));
    LocalMux I__7145 (
            .O(N__40430),
            .I(N__40427));
    Span4Mux_h I__7144 (
            .O(N__40427),
            .I(N__40424));
    Span4Mux_h I__7143 (
            .O(N__40424),
            .I(N__40421));
    Span4Mux_h I__7142 (
            .O(N__40421),
            .I(N__40418));
    Span4Mux_v I__7141 (
            .O(N__40418),
            .I(N__40415));
    Span4Mux_v I__7140 (
            .O(N__40415),
            .I(N__40412));
    Span4Mux_v I__7139 (
            .O(N__40412),
            .I(N__40409));
    IoSpan4Mux I__7138 (
            .O(N__40409),
            .I(N__40406));
    Odrv4 I__7137 (
            .O(N__40406),
            .I(D9_in_c));
    CascadeMux I__7136 (
            .O(N__40403),
            .I(\CONTROL.N_170_cascade_ ));
    InMux I__7135 (
            .O(N__40400),
            .I(N__40397));
    LocalMux I__7134 (
            .O(N__40397),
            .I(N_186));
    InMux I__7133 (
            .O(N__40394),
            .I(N__40391));
    LocalMux I__7132 (
            .O(N__40391),
            .I(\CONTROL.N_202 ));
    CascadeMux I__7131 (
            .O(N__40388),
            .I(N_186_cascade_));
    IoInMux I__7130 (
            .O(N__40385),
            .I(N__40381));
    IoInMux I__7129 (
            .O(N__40384),
            .I(N__40378));
    LocalMux I__7128 (
            .O(N__40381),
            .I(N__40375));
    LocalMux I__7127 (
            .O(N__40378),
            .I(N__40372));
    IoSpan4Mux I__7126 (
            .O(N__40375),
            .I(N__40369));
    IoSpan4Mux I__7125 (
            .O(N__40372),
            .I(N__40366));
    Span4Mux_s1_h I__7124 (
            .O(N__40369),
            .I(N__40363));
    Span4Mux_s2_h I__7123 (
            .O(N__40366),
            .I(N__40360));
    Span4Mux_h I__7122 (
            .O(N__40363),
            .I(N__40357));
    Span4Mux_h I__7121 (
            .O(N__40360),
            .I(N__40354));
    Span4Mux_h I__7120 (
            .O(N__40357),
            .I(N__40350));
    Span4Mux_h I__7119 (
            .O(N__40354),
            .I(N__40347));
    InMux I__7118 (
            .O(N__40353),
            .I(N__40344));
    Span4Mux_h I__7117 (
            .O(N__40350),
            .I(N__40341));
    Span4Mux_h I__7116 (
            .O(N__40347),
            .I(N__40336));
    LocalMux I__7115 (
            .O(N__40344),
            .I(N__40336));
    Span4Mux_h I__7114 (
            .O(N__40341),
            .I(N__40333));
    Span4Mux_v I__7113 (
            .O(N__40336),
            .I(N__40330));
    Span4Mux_v I__7112 (
            .O(N__40333),
            .I(N__40325));
    Span4Mux_v I__7111 (
            .O(N__40330),
            .I(N__40325));
    Odrv4 I__7110 (
            .O(N__40325),
            .I(bus_9));
    InMux I__7109 (
            .O(N__40322),
            .I(N__40319));
    LocalMux I__7108 (
            .O(N__40319),
            .I(N__40316));
    Span4Mux_h I__7107 (
            .O(N__40316),
            .I(N__40313));
    Span4Mux_v I__7106 (
            .O(N__40313),
            .I(N__40310));
    Span4Mux_h I__7105 (
            .O(N__40310),
            .I(N__40306));
    InMux I__7104 (
            .O(N__40309),
            .I(N__40303));
    Odrv4 I__7103 (
            .O(N__40306),
            .I(\CONTROL.ctrlOut_9 ));
    LocalMux I__7102 (
            .O(N__40303),
            .I(\CONTROL.ctrlOut_9 ));
    CascadeMux I__7101 (
            .O(N__40298),
            .I(N__40293));
    InMux I__7100 (
            .O(N__40297),
            .I(N__40287));
    InMux I__7099 (
            .O(N__40296),
            .I(N__40287));
    InMux I__7098 (
            .O(N__40293),
            .I(N__40282));
    InMux I__7097 (
            .O(N__40292),
            .I(N__40282));
    LocalMux I__7096 (
            .O(N__40287),
            .I(N__40279));
    LocalMux I__7095 (
            .O(N__40282),
            .I(N__40276));
    Span4Mux_v I__7094 (
            .O(N__40279),
            .I(N__40273));
    Odrv4 I__7093 (
            .O(N__40276),
            .I(\PROM.ROMDATA.m284 ));
    Odrv4 I__7092 (
            .O(N__40273),
            .I(\PROM.ROMDATA.m284 ));
    InMux I__7091 (
            .O(N__40268),
            .I(N__40264));
    CascadeMux I__7090 (
            .O(N__40267),
            .I(N__40261));
    LocalMux I__7089 (
            .O(N__40264),
            .I(N__40258));
    InMux I__7088 (
            .O(N__40261),
            .I(N__40255));
    Span4Mux_v I__7087 (
            .O(N__40258),
            .I(N__40252));
    LocalMux I__7086 (
            .O(N__40255),
            .I(N__40249));
    Span4Mux_h I__7085 (
            .O(N__40252),
            .I(N__40246));
    Span4Mux_v I__7084 (
            .O(N__40249),
            .I(N__40243));
    Span4Mux_v I__7083 (
            .O(N__40246),
            .I(N__40240));
    Span4Mux_v I__7082 (
            .O(N__40243),
            .I(N__40236));
    Span4Mux_v I__7081 (
            .O(N__40240),
            .I(N__40233));
    InMux I__7080 (
            .O(N__40239),
            .I(N__40230));
    Span4Mux_h I__7079 (
            .O(N__40236),
            .I(N__40227));
    Odrv4 I__7078 (
            .O(N__40233),
            .I(h_5));
    LocalMux I__7077 (
            .O(N__40230),
            .I(h_5));
    Odrv4 I__7076 (
            .O(N__40227),
            .I(h_5));
    InMux I__7075 (
            .O(N__40220),
            .I(N__40216));
    InMux I__7074 (
            .O(N__40219),
            .I(N__40213));
    LocalMux I__7073 (
            .O(N__40216),
            .I(N__40210));
    LocalMux I__7072 (
            .O(N__40213),
            .I(N__40207));
    Span12Mux_v I__7071 (
            .O(N__40210),
            .I(N__40204));
    Span4Mux_h I__7070 (
            .O(N__40207),
            .I(N__40201));
    Odrv12 I__7069 (
            .O(N__40204),
            .I(\ALU.dZ0Z_5 ));
    Odrv4 I__7068 (
            .O(N__40201),
            .I(\ALU.dZ0Z_5 ));
    InMux I__7067 (
            .O(N__40196),
            .I(N__40193));
    LocalMux I__7066 (
            .O(N__40193),
            .I(\ALU.d_RNIBT8EZ0Z_5 ));
    CascadeMux I__7065 (
            .O(N__40190),
            .I(\PROM.ROMDATA.m407_cascade_ ));
    CascadeMux I__7064 (
            .O(N__40187),
            .I(\PROM.ROMDATA.m488_ns_cascade_ ));
    InMux I__7063 (
            .O(N__40184),
            .I(N__40181));
    LocalMux I__7062 (
            .O(N__40181),
            .I(\ALU.lshift_15_0_1 ));
    CascadeMux I__7061 (
            .O(N__40178),
            .I(\ALU.mult_1_cascade_ ));
    InMux I__7060 (
            .O(N__40175),
            .I(N__40172));
    LocalMux I__7059 (
            .O(N__40172),
            .I(N__40169));
    Span4Mux_v I__7058 (
            .O(N__40169),
            .I(N__40166));
    Odrv4 I__7057 (
            .O(N__40166),
            .I(\ALU.a_15_m3_d_ns_1_1 ));
    InMux I__7056 (
            .O(N__40163),
            .I(N__40160));
    LocalMux I__7055 (
            .O(N__40160),
            .I(N__40157));
    Span4Mux_h I__7054 (
            .O(N__40157),
            .I(N__40154));
    Span4Mux_v I__7053 (
            .O(N__40154),
            .I(N__40151));
    Odrv4 I__7052 (
            .O(N__40151),
            .I(\ALU.d_RNIJOQE21Z0Z_0 ));
    InMux I__7051 (
            .O(N__40148),
            .I(N__40145));
    LocalMux I__7050 (
            .O(N__40145),
            .I(N__40141));
    InMux I__7049 (
            .O(N__40144),
            .I(N__40138));
    Span4Mux_v I__7048 (
            .O(N__40141),
            .I(N__40135));
    LocalMux I__7047 (
            .O(N__40138),
            .I(N__40131));
    Span4Mux_h I__7046 (
            .O(N__40135),
            .I(N__40128));
    InMux I__7045 (
            .O(N__40134),
            .I(N__40125));
    Span4Mux_v I__7044 (
            .O(N__40131),
            .I(N__40122));
    Span4Mux_v I__7043 (
            .O(N__40128),
            .I(N__40119));
    LocalMux I__7042 (
            .O(N__40125),
            .I(N__40116));
    Span4Mux_h I__7041 (
            .O(N__40122),
            .I(N__40113));
    Span4Mux_h I__7040 (
            .O(N__40119),
            .I(N__40108));
    Span4Mux_h I__7039 (
            .O(N__40116),
            .I(N__40108));
    Span4Mux_h I__7038 (
            .O(N__40113),
            .I(N__40105));
    Span4Mux_v I__7037 (
            .O(N__40108),
            .I(N__40102));
    Odrv4 I__7036 (
            .O(N__40105),
            .I(g_5));
    Odrv4 I__7035 (
            .O(N__40102),
            .I(g_5));
    InMux I__7034 (
            .O(N__40097),
            .I(N__40094));
    LocalMux I__7033 (
            .O(N__40094),
            .I(N__40091));
    Span4Mux_h I__7032 (
            .O(N__40091),
            .I(N__40087));
    InMux I__7031 (
            .O(N__40090),
            .I(N__40084));
    Span4Mux_v I__7030 (
            .O(N__40087),
            .I(N__40081));
    LocalMux I__7029 (
            .O(N__40084),
            .I(N__40078));
    Span4Mux_h I__7028 (
            .O(N__40081),
            .I(N__40073));
    Span4Mux_v I__7027 (
            .O(N__40078),
            .I(N__40073));
    Odrv4 I__7026 (
            .O(N__40073),
            .I(\ALU.cZ0Z_5 ));
    CascadeMux I__7025 (
            .O(N__40070),
            .I(N__40066));
    InMux I__7024 (
            .O(N__40069),
            .I(N__40063));
    InMux I__7023 (
            .O(N__40066),
            .I(N__40060));
    LocalMux I__7022 (
            .O(N__40063),
            .I(N__40057));
    LocalMux I__7021 (
            .O(N__40060),
            .I(N__40054));
    Span12Mux_h I__7020 (
            .O(N__40057),
            .I(N__40051));
    Span4Mux_h I__7019 (
            .O(N__40054),
            .I(N__40048));
    Odrv12 I__7018 (
            .O(N__40051),
            .I(\ALU.eZ0Z_5 ));
    Odrv4 I__7017 (
            .O(N__40048),
            .I(\ALU.eZ0Z_5 ));
    InMux I__7016 (
            .O(N__40043),
            .I(N__40040));
    LocalMux I__7015 (
            .O(N__40040),
            .I(N__40037));
    Span4Mux_v I__7014 (
            .O(N__40037),
            .I(N__40033));
    InMux I__7013 (
            .O(N__40036),
            .I(N__40030));
    Span4Mux_v I__7012 (
            .O(N__40033),
            .I(N__40027));
    LocalMux I__7011 (
            .O(N__40030),
            .I(N__40024));
    Span4Mux_h I__7010 (
            .O(N__40027),
            .I(N__40021));
    Span4Mux_v I__7009 (
            .O(N__40024),
            .I(N__40018));
    Odrv4 I__7008 (
            .O(N__40021),
            .I(\ALU.aZ0Z_5 ));
    Odrv4 I__7007 (
            .O(N__40018),
            .I(\ALU.aZ0Z_5 ));
    InMux I__7006 (
            .O(N__40013),
            .I(N__40010));
    LocalMux I__7005 (
            .O(N__40010),
            .I(\ALU.c_RNI8KVQZ0Z_5 ));
    CascadeMux I__7004 (
            .O(N__40007),
            .I(\ALU.e_RNI48JMZ0Z_5_cascade_ ));
    CascadeMux I__7003 (
            .O(N__40004),
            .I(\ALU.operand2_7_ns_1_5_cascade_ ));
    InMux I__7002 (
            .O(N__40001),
            .I(N__39998));
    LocalMux I__7001 (
            .O(N__39998),
            .I(N__39995));
    Span4Mux_v I__7000 (
            .O(N__39995),
            .I(N__39992));
    Span4Mux_h I__6999 (
            .O(N__39992),
            .I(N__39989));
    Odrv4 I__6998 (
            .O(N__39989),
            .I(\ALU.operand2_5 ));
    InMux I__6997 (
            .O(N__39986),
            .I(N__39983));
    LocalMux I__6996 (
            .O(N__39983),
            .I(N__39980));
    Span4Mux_v I__6995 (
            .O(N__39980),
            .I(N__39977));
    Span4Mux_v I__6994 (
            .O(N__39977),
            .I(N__39974));
    Span4Mux_h I__6993 (
            .O(N__39974),
            .I(N__39969));
    InMux I__6992 (
            .O(N__39973),
            .I(N__39966));
    CascadeMux I__6991 (
            .O(N__39972),
            .I(N__39963));
    Span4Mux_v I__6990 (
            .O(N__39969),
            .I(N__39960));
    LocalMux I__6989 (
            .O(N__39966),
            .I(N__39957));
    InMux I__6988 (
            .O(N__39963),
            .I(N__39954));
    Span4Mux_v I__6987 (
            .O(N__39960),
            .I(N__39949));
    Span4Mux_h I__6986 (
            .O(N__39957),
            .I(N__39949));
    LocalMux I__6985 (
            .O(N__39954),
            .I(N__39946));
    Span4Mux_v I__6984 (
            .O(N__39949),
            .I(N__39943));
    Span12Mux_v I__6983 (
            .O(N__39946),
            .I(N__39940));
    Span4Mux_v I__6982 (
            .O(N__39943),
            .I(N__39937));
    Odrv12 I__6981 (
            .O(N__39940),
            .I(f_5));
    Odrv4 I__6980 (
            .O(N__39937),
            .I(f_5));
    InMux I__6979 (
            .O(N__39932),
            .I(N__39929));
    LocalMux I__6978 (
            .O(N__39929),
            .I(N__39926));
    Span4Mux_h I__6977 (
            .O(N__39926),
            .I(N__39923));
    Span4Mux_h I__6976 (
            .O(N__39923),
            .I(N__39919));
    InMux I__6975 (
            .O(N__39922),
            .I(N__39916));
    Sp12to4 I__6974 (
            .O(N__39919),
            .I(N__39913));
    LocalMux I__6973 (
            .O(N__39916),
            .I(N__39910));
    Odrv12 I__6972 (
            .O(N__39913),
            .I(\ALU.bZ0Z_5 ));
    Odrv12 I__6971 (
            .O(N__39910),
            .I(\ALU.bZ0Z_5 ));
    InMux I__6970 (
            .O(N__39905),
            .I(N__39902));
    LocalMux I__6969 (
            .O(N__39902),
            .I(\ALU.b_RNI7HSPZ0Z_5 ));
    InMux I__6968 (
            .O(N__39899),
            .I(N__39896));
    LocalMux I__6967 (
            .O(N__39896),
            .I(N__39892));
    CascadeMux I__6966 (
            .O(N__39895),
            .I(N__39889));
    Span4Mux_v I__6965 (
            .O(N__39892),
            .I(N__39886));
    InMux I__6964 (
            .O(N__39889),
            .I(N__39883));
    Sp12to4 I__6963 (
            .O(N__39886),
            .I(N__39880));
    LocalMux I__6962 (
            .O(N__39883),
            .I(N__39877));
    Span12Mux_h I__6961 (
            .O(N__39880),
            .I(N__39874));
    Span4Mux_h I__6960 (
            .O(N__39877),
            .I(N__39871));
    Odrv12 I__6959 (
            .O(N__39874),
            .I(\ALU.bZ0Z_6 ));
    Odrv4 I__6958 (
            .O(N__39871),
            .I(\ALU.bZ0Z_6 ));
    InMux I__6957 (
            .O(N__39866),
            .I(N__39863));
    LocalMux I__6956 (
            .O(N__39863),
            .I(N__39859));
    InMux I__6955 (
            .O(N__39862),
            .I(N__39856));
    Span4Mux_h I__6954 (
            .O(N__39859),
            .I(N__39851));
    LocalMux I__6953 (
            .O(N__39856),
            .I(N__39851));
    Span4Mux_v I__6952 (
            .O(N__39851),
            .I(N__39848));
    Sp12to4 I__6951 (
            .O(N__39848),
            .I(N__39845));
    Odrv12 I__6950 (
            .O(N__39845),
            .I(\ALU.bZ0Z_3 ));
    InMux I__6949 (
            .O(N__39842),
            .I(N__39836));
    InMux I__6948 (
            .O(N__39841),
            .I(N__39836));
    LocalMux I__6947 (
            .O(N__39836),
            .I(N__39833));
    Span4Mux_h I__6946 (
            .O(N__39833),
            .I(N__39830));
    Span4Mux_h I__6945 (
            .O(N__39830),
            .I(N__39827));
    Sp12to4 I__6944 (
            .O(N__39827),
            .I(N__39824));
    Span12Mux_v I__6943 (
            .O(N__39824),
            .I(N__39821));
    Odrv12 I__6942 (
            .O(N__39821),
            .I(\ALU.bZ0Z_11 ));
    InMux I__6941 (
            .O(N__39818),
            .I(N__39814));
    InMux I__6940 (
            .O(N__39817),
            .I(N__39811));
    LocalMux I__6939 (
            .O(N__39814),
            .I(N__39808));
    LocalMux I__6938 (
            .O(N__39811),
            .I(N__39805));
    Span4Mux_v I__6937 (
            .O(N__39808),
            .I(N__39802));
    Span4Mux_v I__6936 (
            .O(N__39805),
            .I(N__39799));
    Span4Mux_h I__6935 (
            .O(N__39802),
            .I(N__39796));
    Span4Mux_h I__6934 (
            .O(N__39799),
            .I(N__39793));
    Span4Mux_h I__6933 (
            .O(N__39796),
            .I(N__39790));
    Sp12to4 I__6932 (
            .O(N__39793),
            .I(N__39787));
    Sp12to4 I__6931 (
            .O(N__39790),
            .I(N__39782));
    Span12Mux_s7_h I__6930 (
            .O(N__39787),
            .I(N__39782));
    Odrv12 I__6929 (
            .O(N__39782),
            .I(\ALU.bZ0Z_12 ));
    InMux I__6928 (
            .O(N__39779),
            .I(N__39776));
    LocalMux I__6927 (
            .O(N__39776),
            .I(N__39773));
    Span4Mux_v I__6926 (
            .O(N__39773),
            .I(N__39770));
    Span4Mux_v I__6925 (
            .O(N__39770),
            .I(N__39767));
    Odrv4 I__6924 (
            .O(N__39767),
            .I(\CONTROL.gZ0Z3 ));
    InMux I__6923 (
            .O(N__39764),
            .I(N__39761));
    LocalMux I__6922 (
            .O(N__39761),
            .I(N__39758));
    Span4Mux_v I__6921 (
            .O(N__39758),
            .I(N__39755));
    Odrv4 I__6920 (
            .O(N__39755),
            .I(\ALU.lshift_15_0_sx_1 ));
    IoInMux I__6919 (
            .O(N__39752),
            .I(N__39748));
    IoInMux I__6918 (
            .O(N__39751),
            .I(N__39745));
    LocalMux I__6917 (
            .O(N__39748),
            .I(N__39742));
    LocalMux I__6916 (
            .O(N__39745),
            .I(N__39739));
    Span4Mux_s0_h I__6915 (
            .O(N__39742),
            .I(N__39736));
    IoSpan4Mux I__6914 (
            .O(N__39739),
            .I(N__39733));
    Sp12to4 I__6913 (
            .O(N__39736),
            .I(N__39729));
    Sp12to4 I__6912 (
            .O(N__39733),
            .I(N__39726));
    InMux I__6911 (
            .O(N__39732),
            .I(N__39723));
    Span12Mux_v I__6910 (
            .O(N__39729),
            .I(N__39720));
    Span12Mux_s7_h I__6909 (
            .O(N__39726),
            .I(N__39715));
    LocalMux I__6908 (
            .O(N__39723),
            .I(N__39715));
    Span12Mux_h I__6907 (
            .O(N__39720),
            .I(N__39710));
    Span12Mux_h I__6906 (
            .O(N__39715),
            .I(N__39710));
    Odrv12 I__6905 (
            .O(N__39710),
            .I(bus_14));
    CascadeMux I__6904 (
            .O(N__39707),
            .I(\ALU.lshift_15_0_1_cascade_ ));
    InMux I__6903 (
            .O(N__39704),
            .I(N__39701));
    LocalMux I__6902 (
            .O(N__39701),
            .I(\ALU.a_15_m0_sx_14 ));
    InMux I__6901 (
            .O(N__39698),
            .I(N__39695));
    LocalMux I__6900 (
            .O(N__39695),
            .I(\ALU.c_RNI890LZ0Z_13 ));
    CascadeMux I__6899 (
            .O(N__39692),
            .I(\ALU.a_RNI4P741Z0Z_13_cascade_ ));
    InMux I__6898 (
            .O(N__39689),
            .I(N__39686));
    LocalMux I__6897 (
            .O(N__39686),
            .I(\ALU.d_RNIAHCTZ0Z_13 ));
    CascadeMux I__6896 (
            .O(N__39683),
            .I(\ALU.operand2_7_ns_1_13_cascade_ ));
    InMux I__6895 (
            .O(N__39680),
            .I(N__39677));
    LocalMux I__6894 (
            .O(N__39677),
            .I(\ALU.b_RNI61KC1Z0Z_13 ));
    InMux I__6893 (
            .O(N__39674),
            .I(N__39671));
    LocalMux I__6892 (
            .O(N__39671),
            .I(N__39668));
    Span4Mux_h I__6891 (
            .O(N__39668),
            .I(N__39665));
    Span4Mux_h I__6890 (
            .O(N__39665),
            .I(N__39662));
    Span4Mux_v I__6889 (
            .O(N__39662),
            .I(N__39659));
    Odrv4 I__6888 (
            .O(N__39659),
            .I(\ALU.operand2_13 ));
    InMux I__6887 (
            .O(N__39656),
            .I(N__39653));
    LocalMux I__6886 (
            .O(N__39653),
            .I(N__39648));
    InMux I__6885 (
            .O(N__39652),
            .I(N__39645));
    InMux I__6884 (
            .O(N__39651),
            .I(N__39642));
    Span4Mux_v I__6883 (
            .O(N__39648),
            .I(N__39637));
    LocalMux I__6882 (
            .O(N__39645),
            .I(N__39637));
    LocalMux I__6881 (
            .O(N__39642),
            .I(N__39634));
    Span4Mux_v I__6880 (
            .O(N__39637),
            .I(N__39631));
    Span4Mux_v I__6879 (
            .O(N__39634),
            .I(N__39628));
    Span4Mux_v I__6878 (
            .O(N__39631),
            .I(N__39625));
    Span4Mux_v I__6877 (
            .O(N__39628),
            .I(N__39622));
    Span4Mux_h I__6876 (
            .O(N__39625),
            .I(N__39619));
    Odrv4 I__6875 (
            .O(N__39622),
            .I(bus_0_13));
    Odrv4 I__6874 (
            .O(N__39619),
            .I(bus_0_13));
    CascadeMux I__6873 (
            .O(N__39614),
            .I(\ALU.operand2_13_cascade_ ));
    InMux I__6872 (
            .O(N__39611),
            .I(N__39608));
    LocalMux I__6871 (
            .O(N__39608),
            .I(N__39600));
    InMux I__6870 (
            .O(N__39607),
            .I(N__39595));
    InMux I__6869 (
            .O(N__39606),
            .I(N__39592));
    InMux I__6868 (
            .O(N__39605),
            .I(N__39589));
    InMux I__6867 (
            .O(N__39604),
            .I(N__39586));
    InMux I__6866 (
            .O(N__39603),
            .I(N__39583));
    Span4Mux_h I__6865 (
            .O(N__39600),
            .I(N__39580));
    InMux I__6864 (
            .O(N__39599),
            .I(N__39577));
    InMux I__6863 (
            .O(N__39598),
            .I(N__39574));
    LocalMux I__6862 (
            .O(N__39595),
            .I(N__39571));
    LocalMux I__6861 (
            .O(N__39592),
            .I(N__39568));
    LocalMux I__6860 (
            .O(N__39589),
            .I(N__39565));
    LocalMux I__6859 (
            .O(N__39586),
            .I(N__39558));
    LocalMux I__6858 (
            .O(N__39583),
            .I(N__39558));
    Span4Mux_v I__6857 (
            .O(N__39580),
            .I(N__39558));
    LocalMux I__6856 (
            .O(N__39577),
            .I(N__39551));
    LocalMux I__6855 (
            .O(N__39574),
            .I(N__39551));
    Span4Mux_v I__6854 (
            .O(N__39571),
            .I(N__39551));
    Span4Mux_h I__6853 (
            .O(N__39568),
            .I(N__39544));
    Span4Mux_v I__6852 (
            .O(N__39565),
            .I(N__39544));
    Span4Mux_h I__6851 (
            .O(N__39558),
            .I(N__39544));
    Odrv4 I__6850 (
            .O(N__39551),
            .I(\ALU.d_RNI02EVNBZ0Z_4 ));
    Odrv4 I__6849 (
            .O(N__39544),
            .I(\ALU.d_RNI02EVNBZ0Z_4 ));
    InMux I__6848 (
            .O(N__39539),
            .I(N__39536));
    LocalMux I__6847 (
            .O(N__39536),
            .I(N__39532));
    InMux I__6846 (
            .O(N__39535),
            .I(N__39527));
    Span4Mux_h I__6845 (
            .O(N__39532),
            .I(N__39524));
    InMux I__6844 (
            .O(N__39531),
            .I(N__39521));
    InMux I__6843 (
            .O(N__39530),
            .I(N__39518));
    LocalMux I__6842 (
            .O(N__39527),
            .I(N__39511));
    Span4Mux_h I__6841 (
            .O(N__39524),
            .I(N__39504));
    LocalMux I__6840 (
            .O(N__39521),
            .I(N__39504));
    LocalMux I__6839 (
            .O(N__39518),
            .I(N__39504));
    InMux I__6838 (
            .O(N__39517),
            .I(N__39501));
    InMux I__6837 (
            .O(N__39516),
            .I(N__39498));
    InMux I__6836 (
            .O(N__39515),
            .I(N__39495));
    InMux I__6835 (
            .O(N__39514),
            .I(N__39492));
    Odrv4 I__6834 (
            .O(N__39511),
            .I(\ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ));
    Odrv4 I__6833 (
            .O(N__39504),
            .I(\ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ));
    LocalMux I__6832 (
            .O(N__39501),
            .I(\ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ));
    LocalMux I__6831 (
            .O(N__39498),
            .I(\ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ));
    LocalMux I__6830 (
            .O(N__39495),
            .I(\ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ));
    LocalMux I__6829 (
            .O(N__39492),
            .I(\ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ));
    InMux I__6828 (
            .O(N__39479),
            .I(N__39476));
    LocalMux I__6827 (
            .O(N__39476),
            .I(N__39472));
    InMux I__6826 (
            .O(N__39475),
            .I(N__39469));
    Span4Mux_v I__6825 (
            .O(N__39472),
            .I(N__39465));
    LocalMux I__6824 (
            .O(N__39469),
            .I(N__39462));
    InMux I__6823 (
            .O(N__39468),
            .I(N__39459));
    Span4Mux_h I__6822 (
            .O(N__39465),
            .I(N__39450));
    Span4Mux_h I__6821 (
            .O(N__39462),
            .I(N__39450));
    LocalMux I__6820 (
            .O(N__39459),
            .I(N__39447));
    InMux I__6819 (
            .O(N__39458),
            .I(N__39444));
    InMux I__6818 (
            .O(N__39457),
            .I(N__39441));
    InMux I__6817 (
            .O(N__39456),
            .I(N__39438));
    InMux I__6816 (
            .O(N__39455),
            .I(N__39435));
    Odrv4 I__6815 (
            .O(N__39450),
            .I(\ALU.addsub_cry_1_c_RNIICPECZ0Z7 ));
    Odrv4 I__6814 (
            .O(N__39447),
            .I(\ALU.addsub_cry_1_c_RNIICPECZ0Z7 ));
    LocalMux I__6813 (
            .O(N__39444),
            .I(\ALU.addsub_cry_1_c_RNIICPECZ0Z7 ));
    LocalMux I__6812 (
            .O(N__39441),
            .I(\ALU.addsub_cry_1_c_RNIICPECZ0Z7 ));
    LocalMux I__6811 (
            .O(N__39438),
            .I(\ALU.addsub_cry_1_c_RNIICPECZ0Z7 ));
    LocalMux I__6810 (
            .O(N__39435),
            .I(\ALU.addsub_cry_1_c_RNIICPECZ0Z7 ));
    CascadeMux I__6809 (
            .O(N__39422),
            .I(N__39419));
    InMux I__6808 (
            .O(N__39419),
            .I(N__39416));
    LocalMux I__6807 (
            .O(N__39416),
            .I(N__39412));
    InMux I__6806 (
            .O(N__39415),
            .I(N__39409));
    Span4Mux_v I__6805 (
            .O(N__39412),
            .I(N__39404));
    LocalMux I__6804 (
            .O(N__39409),
            .I(N__39404));
    Span4Mux_h I__6803 (
            .O(N__39404),
            .I(N__39401));
    Span4Mux_h I__6802 (
            .O(N__39401),
            .I(N__39398));
    Odrv4 I__6801 (
            .O(N__39398),
            .I(\ALU.bZ0Z_2 ));
    InMux I__6800 (
            .O(N__39395),
            .I(N__39388));
    InMux I__6799 (
            .O(N__39394),
            .I(N__39384));
    InMux I__6798 (
            .O(N__39393),
            .I(N__39381));
    InMux I__6797 (
            .O(N__39392),
            .I(N__39378));
    InMux I__6796 (
            .O(N__39391),
            .I(N__39374));
    LocalMux I__6795 (
            .O(N__39388),
            .I(N__39371));
    InMux I__6794 (
            .O(N__39387),
            .I(N__39368));
    LocalMux I__6793 (
            .O(N__39384),
            .I(N__39365));
    LocalMux I__6792 (
            .O(N__39381),
            .I(N__39360));
    LocalMux I__6791 (
            .O(N__39378),
            .I(N__39360));
    InMux I__6790 (
            .O(N__39377),
            .I(N__39357));
    LocalMux I__6789 (
            .O(N__39374),
            .I(N__39354));
    Span4Mux_v I__6788 (
            .O(N__39371),
            .I(N__39351));
    LocalMux I__6787 (
            .O(N__39368),
            .I(N__39346));
    Span4Mux_v I__6786 (
            .O(N__39365),
            .I(N__39346));
    Span4Mux_v I__6785 (
            .O(N__39360),
            .I(N__39343));
    LocalMux I__6784 (
            .O(N__39357),
            .I(N__39340));
    Span4Mux_v I__6783 (
            .O(N__39354),
            .I(N__39335));
    Span4Mux_h I__6782 (
            .O(N__39351),
            .I(N__39335));
    Span4Mux_h I__6781 (
            .O(N__39346),
            .I(N__39330));
    Span4Mux_h I__6780 (
            .O(N__39343),
            .I(N__39330));
    Odrv4 I__6779 (
            .O(N__39340),
            .I(\ALU.addsub_cry_3_c_RNIM4CUTZ0Z9 ));
    Odrv4 I__6778 (
            .O(N__39335),
            .I(\ALU.addsub_cry_3_c_RNIM4CUTZ0Z9 ));
    Odrv4 I__6777 (
            .O(N__39330),
            .I(\ALU.addsub_cry_3_c_RNIM4CUTZ0Z9 ));
    InMux I__6776 (
            .O(N__39323),
            .I(N__39316));
    InMux I__6775 (
            .O(N__39322),
            .I(N__39311));
    InMux I__6774 (
            .O(N__39321),
            .I(N__39308));
    InMux I__6773 (
            .O(N__39320),
            .I(N__39305));
    InMux I__6772 (
            .O(N__39319),
            .I(N__39302));
    LocalMux I__6771 (
            .O(N__39316),
            .I(N__39298));
    InMux I__6770 (
            .O(N__39315),
            .I(N__39295));
    InMux I__6769 (
            .O(N__39314),
            .I(N__39292));
    LocalMux I__6768 (
            .O(N__39311),
            .I(N__39289));
    LocalMux I__6767 (
            .O(N__39308),
            .I(N__39286));
    LocalMux I__6766 (
            .O(N__39305),
            .I(N__39283));
    LocalMux I__6765 (
            .O(N__39302),
            .I(N__39280));
    InMux I__6764 (
            .O(N__39301),
            .I(N__39277));
    Span4Mux_h I__6763 (
            .O(N__39298),
            .I(N__39274));
    LocalMux I__6762 (
            .O(N__39295),
            .I(N__39265));
    LocalMux I__6761 (
            .O(N__39292),
            .I(N__39265));
    Span4Mux_h I__6760 (
            .O(N__39289),
            .I(N__39265));
    Span4Mux_v I__6759 (
            .O(N__39286),
            .I(N__39265));
    Span4Mux_h I__6758 (
            .O(N__39283),
            .I(N__39260));
    Span4Mux_h I__6757 (
            .O(N__39280),
            .I(N__39260));
    LocalMux I__6756 (
            .O(N__39277),
            .I(\ALU.addsub_cry_4_c_RNI5L6IQAZ0 ));
    Odrv4 I__6755 (
            .O(N__39274),
            .I(\ALU.addsub_cry_4_c_RNI5L6IQAZ0 ));
    Odrv4 I__6754 (
            .O(N__39265),
            .I(\ALU.addsub_cry_4_c_RNI5L6IQAZ0 ));
    Odrv4 I__6753 (
            .O(N__39260),
            .I(\ALU.addsub_cry_4_c_RNI5L6IQAZ0 ));
    InMux I__6752 (
            .O(N__39251),
            .I(N__39248));
    LocalMux I__6751 (
            .O(N__39248),
            .I(N__39245));
    Span4Mux_v I__6750 (
            .O(N__39245),
            .I(N__39241));
    InMux I__6749 (
            .O(N__39244),
            .I(N__39238));
    Odrv4 I__6748 (
            .O(N__39241),
            .I(\ALU.N_1025 ));
    LocalMux I__6747 (
            .O(N__39238),
            .I(\ALU.N_1025 ));
    InMux I__6746 (
            .O(N__39233),
            .I(N__39230));
    LocalMux I__6745 (
            .O(N__39230),
            .I(N__39226));
    InMux I__6744 (
            .O(N__39229),
            .I(N__39223));
    Span4Mux_h I__6743 (
            .O(N__39226),
            .I(N__39218));
    LocalMux I__6742 (
            .O(N__39223),
            .I(N__39218));
    Span4Mux_h I__6741 (
            .O(N__39218),
            .I(N__39215));
    Odrv4 I__6740 (
            .O(N__39215),
            .I(\ALU.N_864 ));
    CascadeMux I__6739 (
            .O(N__39212),
            .I(\ALU.N_965_cascade_ ));
    InMux I__6738 (
            .O(N__39209),
            .I(N__39206));
    LocalMux I__6737 (
            .O(N__39206),
            .I(N__39203));
    Odrv4 I__6736 (
            .O(N__39203),
            .I(\ALU.d_RNIFHCRU4Z0Z_2 ));
    InMux I__6735 (
            .O(N__39200),
            .I(N__39197));
    LocalMux I__6734 (
            .O(N__39197),
            .I(N__39194));
    Span4Mux_v I__6733 (
            .O(N__39194),
            .I(N__39191));
    Odrv4 I__6732 (
            .O(N__39191),
            .I(\ALU.mult_15_15 ));
    InMux I__6731 (
            .O(N__39188),
            .I(N__39185));
    LocalMux I__6730 (
            .O(N__39185),
            .I(\ALU.c_RNINT9PO2Z0Z_10 ));
    InMux I__6729 (
            .O(N__39182),
            .I(N__39179));
    LocalMux I__6728 (
            .O(N__39179),
            .I(\ALU.mult_13 ));
    InMux I__6727 (
            .O(N__39176),
            .I(N__39172));
    InMux I__6726 (
            .O(N__39175),
            .I(N__39169));
    LocalMux I__6725 (
            .O(N__39172),
            .I(N__39166));
    LocalMux I__6724 (
            .O(N__39169),
            .I(N__39163));
    Span4Mux_h I__6723 (
            .O(N__39166),
            .I(N__39160));
    Span4Mux_h I__6722 (
            .O(N__39163),
            .I(N__39155));
    Span4Mux_h I__6721 (
            .O(N__39160),
            .I(N__39155));
    Odrv4 I__6720 (
            .O(N__39155),
            .I(\ALU.N_642 ));
    CascadeMux I__6719 (
            .O(N__39152),
            .I(\ALU.d_RNIULN025Z0Z_2_cascade_ ));
    InMux I__6718 (
            .O(N__39149),
            .I(N__39146));
    LocalMux I__6717 (
            .O(N__39146),
            .I(\ALU.d_RNIULN025_0Z0Z_2 ));
    CascadeMux I__6716 (
            .O(N__39143),
            .I(\ALU.lshift_10_cascade_ ));
    CascadeMux I__6715 (
            .O(N__39140),
            .I(\ALU.c_RNIO0KOKEZ0Z_10_cascade_ ));
    InMux I__6714 (
            .O(N__39137),
            .I(N__39134));
    LocalMux I__6713 (
            .O(N__39134),
            .I(N__39130));
    InMux I__6712 (
            .O(N__39133),
            .I(N__39127));
    Span4Mux_v I__6711 (
            .O(N__39130),
            .I(N__39122));
    LocalMux I__6710 (
            .O(N__39127),
            .I(N__39122));
    Span4Mux_h I__6709 (
            .O(N__39122),
            .I(N__39119));
    Span4Mux_h I__6708 (
            .O(N__39119),
            .I(N__39116));
    Sp12to4 I__6707 (
            .O(N__39116),
            .I(N__39113));
    Span12Mux_v I__6706 (
            .O(N__39113),
            .I(N__39110));
    Span12Mux_h I__6705 (
            .O(N__39110),
            .I(N__39107));
    Odrv12 I__6704 (
            .O(N__39107),
            .I(\ALU.bZ0Z_10 ));
    CascadeMux I__6703 (
            .O(N__39104),
            .I(\ALU.lshift_3_ns_1_15_cascade_ ));
    InMux I__6702 (
            .O(N__39101),
            .I(N__39097));
    InMux I__6701 (
            .O(N__39100),
            .I(N__39092));
    LocalMux I__6700 (
            .O(N__39097),
            .I(N__39083));
    InMux I__6699 (
            .O(N__39096),
            .I(N__39078));
    InMux I__6698 (
            .O(N__39095),
            .I(N__39078));
    LocalMux I__6697 (
            .O(N__39092),
            .I(N__39075));
    InMux I__6696 (
            .O(N__39091),
            .I(N__39068));
    InMux I__6695 (
            .O(N__39090),
            .I(N__39068));
    InMux I__6694 (
            .O(N__39089),
            .I(N__39068));
    InMux I__6693 (
            .O(N__39088),
            .I(N__39061));
    InMux I__6692 (
            .O(N__39087),
            .I(N__39061));
    InMux I__6691 (
            .O(N__39086),
            .I(N__39061));
    Span4Mux_h I__6690 (
            .O(N__39083),
            .I(N__39058));
    LocalMux I__6689 (
            .O(N__39078),
            .I(\ALU.d_RNI64MA6Z0Z_0 ));
    Odrv4 I__6688 (
            .O(N__39075),
            .I(\ALU.d_RNI64MA6Z0Z_0 ));
    LocalMux I__6687 (
            .O(N__39068),
            .I(\ALU.d_RNI64MA6Z0Z_0 ));
    LocalMux I__6686 (
            .O(N__39061),
            .I(\ALU.d_RNI64MA6Z0Z_0 ));
    Odrv4 I__6685 (
            .O(N__39058),
            .I(\ALU.d_RNI64MA6Z0Z_0 ));
    CascadeMux I__6684 (
            .O(N__39047),
            .I(N__39041));
    CascadeMux I__6683 (
            .O(N__39046),
            .I(N__39037));
    CascadeMux I__6682 (
            .O(N__39045),
            .I(N__39034));
    CascadeMux I__6681 (
            .O(N__39044),
            .I(N__39031));
    InMux I__6680 (
            .O(N__39041),
            .I(N__39028));
    InMux I__6679 (
            .O(N__39040),
            .I(N__39020));
    InMux I__6678 (
            .O(N__39037),
            .I(N__39013));
    InMux I__6677 (
            .O(N__39034),
            .I(N__39013));
    InMux I__6676 (
            .O(N__39031),
            .I(N__39013));
    LocalMux I__6675 (
            .O(N__39028),
            .I(N__39010));
    InMux I__6674 (
            .O(N__39027),
            .I(N__39005));
    InMux I__6673 (
            .O(N__39026),
            .I(N__39005));
    InMux I__6672 (
            .O(N__39025),
            .I(N__38998));
    InMux I__6671 (
            .O(N__39024),
            .I(N__38998));
    InMux I__6670 (
            .O(N__39023),
            .I(N__38998));
    LocalMux I__6669 (
            .O(N__39020),
            .I(N__38993));
    LocalMux I__6668 (
            .O(N__39013),
            .I(N__38993));
    Span4Mux_h I__6667 (
            .O(N__39010),
            .I(N__38990));
    LocalMux I__6666 (
            .O(N__39005),
            .I(N_225_0));
    LocalMux I__6665 (
            .O(N__38998),
            .I(N_225_0));
    Odrv4 I__6664 (
            .O(N__38993),
            .I(N_225_0));
    Odrv4 I__6663 (
            .O(N__38990),
            .I(N_225_0));
    InMux I__6662 (
            .O(N__38981),
            .I(N__38978));
    LocalMux I__6661 (
            .O(N__38978),
            .I(N__38974));
    CascadeMux I__6660 (
            .O(N__38977),
            .I(N__38971));
    Span4Mux_v I__6659 (
            .O(N__38974),
            .I(N__38968));
    InMux I__6658 (
            .O(N__38971),
            .I(N__38965));
    Odrv4 I__6657 (
            .O(N__38968),
            .I(\ALU.mult_25_12 ));
    LocalMux I__6656 (
            .O(N__38965),
            .I(\ALU.mult_25_12 ));
    CascadeMux I__6655 (
            .O(N__38960),
            .I(\ALU.mult_13_12_cascade_ ));
    InMux I__6654 (
            .O(N__38957),
            .I(N__38954));
    LocalMux I__6653 (
            .O(N__38954),
            .I(\ALU.mult_467_c_RNICRDK6BZ0 ));
    CascadeMux I__6652 (
            .O(N__38951),
            .I(N__38948));
    InMux I__6651 (
            .O(N__38948),
            .I(N__38945));
    LocalMux I__6650 (
            .O(N__38945),
            .I(\ALU.mult_13_12 ));
    CascadeMux I__6649 (
            .O(N__38942),
            .I(N__38939));
    InMux I__6648 (
            .O(N__38939),
            .I(N__38936));
    LocalMux I__6647 (
            .O(N__38936),
            .I(N__38933));
    Odrv12 I__6646 (
            .O(N__38933),
            .I(\ALU.mult_13_13 ));
    CascadeMux I__6645 (
            .O(N__38930),
            .I(N__38927));
    InMux I__6644 (
            .O(N__38927),
            .I(N__38924));
    LocalMux I__6643 (
            .O(N__38924),
            .I(\ALU.mult_27_13 ));
    InMux I__6642 (
            .O(N__38921),
            .I(\ALU.mult_27_c12 ));
    CascadeMux I__6641 (
            .O(N__38918),
            .I(N__38915));
    InMux I__6640 (
            .O(N__38915),
            .I(N__38912));
    LocalMux I__6639 (
            .O(N__38912),
            .I(\ALU.mult_365_c_RNI8ALOZ0Z96 ));
    CascadeMux I__6638 (
            .O(N__38909),
            .I(N__38906));
    InMux I__6637 (
            .O(N__38906),
            .I(N__38903));
    LocalMux I__6636 (
            .O(N__38903),
            .I(\ALU.mult_27_14 ));
    InMux I__6635 (
            .O(N__38900),
            .I(\ALU.mult_27_c13 ));
    InMux I__6634 (
            .O(N__38897),
            .I(\ALU.mult_27_c14 ));
    CascadeMux I__6633 (
            .O(N__38894),
            .I(N__38891));
    InMux I__6632 (
            .O(N__38891),
            .I(N__38888));
    LocalMux I__6631 (
            .O(N__38888),
            .I(N__38885));
    Odrv4 I__6630 (
            .O(N__38885),
            .I(\ALU.mult_27_c14_THRU_CO ));
    CascadeMux I__6629 (
            .O(N__38882),
            .I(N__38879));
    InMux I__6628 (
            .O(N__38879),
            .I(N__38876));
    LocalMux I__6627 (
            .O(N__38876),
            .I(\ALU.mult_9 ));
    CascadeMux I__6626 (
            .O(N__38873),
            .I(N__38870));
    InMux I__6625 (
            .O(N__38870),
            .I(N__38864));
    InMux I__6624 (
            .O(N__38869),
            .I(N__38864));
    LocalMux I__6623 (
            .O(N__38864),
            .I(N__38861));
    Span4Mux_h I__6622 (
            .O(N__38861),
            .I(N__38858));
    Odrv4 I__6621 (
            .O(N__38858),
            .I(\PROM.ROMDATA.m382_ns ));
    InMux I__6620 (
            .O(N__38855),
            .I(N__38852));
    LocalMux I__6619 (
            .O(N__38852),
            .I(N__38849));
    Span12Mux_v I__6618 (
            .O(N__38849),
            .I(N__38844));
    InMux I__6617 (
            .O(N__38848),
            .I(N__38839));
    InMux I__6616 (
            .O(N__38847),
            .I(N__38839));
    Odrv12 I__6615 (
            .O(N__38844),
            .I(busState_1_RNIAR0U1_2));
    LocalMux I__6614 (
            .O(N__38839),
            .I(busState_1_RNIAR0U1_2));
    CascadeMux I__6613 (
            .O(N__38834),
            .I(N_225_0_cascade_));
    InMux I__6612 (
            .O(N__38831),
            .I(N__38828));
    LocalMux I__6611 (
            .O(N__38828),
            .I(\ALU.mult_13_15 ));
    CascadeMux I__6610 (
            .O(N__38825),
            .I(\ALU.mult_15_14_cascade_ ));
    InMux I__6609 (
            .O(N__38822),
            .I(N__38818));
    InMux I__6608 (
            .O(N__38821),
            .I(N__38815));
    LocalMux I__6607 (
            .O(N__38818),
            .I(\ALU.mult_13_14 ));
    LocalMux I__6606 (
            .O(N__38815),
            .I(\ALU.mult_13_14 ));
    CascadeMux I__6605 (
            .O(N__38810),
            .I(N__38807));
    InMux I__6604 (
            .O(N__38807),
            .I(N__38804));
    LocalMux I__6603 (
            .O(N__38804),
            .I(\CONTROL.N_304_0 ));
    InMux I__6602 (
            .O(N__38801),
            .I(N__38795));
    InMux I__6601 (
            .O(N__38800),
            .I(N__38795));
    LocalMux I__6600 (
            .O(N__38795),
            .I(N__38792));
    Span4Mux_h I__6599 (
            .O(N__38792),
            .I(N__38789));
    Span4Mux_h I__6598 (
            .O(N__38789),
            .I(N__38786));
    Sp12to4 I__6597 (
            .O(N__38786),
            .I(N__38783));
    Odrv12 I__6596 (
            .O(N__38783),
            .I(\PROM.ROMDATA.m433_ns ));
    CascadeMux I__6595 (
            .O(N__38780),
            .I(\PROM.ROMDATA.m294_bm_cascade_ ));
    CascadeMux I__6594 (
            .O(N__38777),
            .I(\PROM.ROMDATA.m31_cascade_ ));
    InMux I__6593 (
            .O(N__38774),
            .I(N__38771));
    LocalMux I__6592 (
            .O(N__38771),
            .I(N__38768));
    Span4Mux_v I__6591 (
            .O(N__38768),
            .I(N__38765));
    Span4Mux_h I__6590 (
            .O(N__38765),
            .I(N__38761));
    InMux I__6589 (
            .O(N__38764),
            .I(N__38758));
    Odrv4 I__6588 (
            .O(N__38761),
            .I(\CONTROL.ctrlOut_12 ));
    LocalMux I__6587 (
            .O(N__38758),
            .I(\CONTROL.ctrlOut_12 ));
    InMux I__6586 (
            .O(N__38753),
            .I(N__38750));
    LocalMux I__6585 (
            .O(N__38750),
            .I(\CONTROL.dout_reto_12 ));
    CascadeMux I__6584 (
            .O(N__38747),
            .I(\PROM.ROMDATA.m391_cascade_ ));
    InMux I__6583 (
            .O(N__38744),
            .I(N__38741));
    LocalMux I__6582 (
            .O(N__38741),
            .I(\PROM.ROMDATA.m433_bm ));
    CascadeMux I__6581 (
            .O(N__38738),
            .I(controlWord_4_cascade_));
    InMux I__6580 (
            .O(N__38735),
            .I(N__38731));
    InMux I__6579 (
            .O(N__38734),
            .I(N__38728));
    LocalMux I__6578 (
            .O(N__38731),
            .I(\CONTROL.N_5_0 ));
    LocalMux I__6577 (
            .O(N__38728),
            .I(\CONTROL.N_5_0 ));
    InMux I__6576 (
            .O(N__38723),
            .I(N__38720));
    LocalMux I__6575 (
            .O(N__38720),
            .I(\CONTROL.g0_12_1 ));
    InMux I__6574 (
            .O(N__38717),
            .I(N__38710));
    InMux I__6573 (
            .O(N__38716),
            .I(N__38707));
    InMux I__6572 (
            .O(N__38715),
            .I(N__38700));
    InMux I__6571 (
            .O(N__38714),
            .I(N__38700));
    InMux I__6570 (
            .O(N__38713),
            .I(N__38700));
    LocalMux I__6569 (
            .O(N__38710),
            .I(N__38696));
    LocalMux I__6568 (
            .O(N__38707),
            .I(N__38693));
    LocalMux I__6567 (
            .O(N__38700),
            .I(N__38690));
    InMux I__6566 (
            .O(N__38699),
            .I(N__38687));
    Span4Mux_h I__6565 (
            .O(N__38696),
            .I(N__38684));
    Span4Mux_v I__6564 (
            .O(N__38693),
            .I(N__38679));
    Span4Mux_v I__6563 (
            .O(N__38690),
            .I(N__38679));
    LocalMux I__6562 (
            .O(N__38687),
            .I(N__38675));
    Span4Mux_v I__6561 (
            .O(N__38684),
            .I(N__38672));
    Span4Mux_h I__6560 (
            .O(N__38679),
            .I(N__38669));
    InMux I__6559 (
            .O(N__38678),
            .I(N__38666));
    Odrv12 I__6558 (
            .O(N__38675),
            .I(\CONTROL.N_360 ));
    Odrv4 I__6557 (
            .O(N__38672),
            .I(\CONTROL.N_360 ));
    Odrv4 I__6556 (
            .O(N__38669),
            .I(\CONTROL.N_360 ));
    LocalMux I__6555 (
            .O(N__38666),
            .I(\CONTROL.N_360 ));
    CascadeMux I__6554 (
            .O(N__38657),
            .I(N__38654));
    InMux I__6553 (
            .O(N__38654),
            .I(N__38651));
    LocalMux I__6552 (
            .O(N__38651),
            .I(N__38648));
    Span4Mux_h I__6551 (
            .O(N__38648),
            .I(N__38645));
    Span4Mux_v I__6550 (
            .O(N__38645),
            .I(N__38641));
    InMux I__6549 (
            .O(N__38644),
            .I(N__38638));
    Odrv4 I__6548 (
            .O(N__38641),
            .I(\CONTROL.N_362 ));
    LocalMux I__6547 (
            .O(N__38638),
            .I(\CONTROL.N_362 ));
    InMux I__6546 (
            .O(N__38633),
            .I(N__38630));
    LocalMux I__6545 (
            .O(N__38630),
            .I(N__38627));
    Odrv4 I__6544 (
            .O(N__38627),
            .I(\CONTROL.m28_0_120_i_i_0 ));
    InMux I__6543 (
            .O(N__38624),
            .I(N__38620));
    InMux I__6542 (
            .O(N__38623),
            .I(N__38617));
    LocalMux I__6541 (
            .O(N__38620),
            .I(N__38614));
    LocalMux I__6540 (
            .O(N__38617),
            .I(N__38611));
    Odrv12 I__6539 (
            .O(N__38614),
            .I(\CONTROL.N_321 ));
    Odrv4 I__6538 (
            .O(N__38611),
            .I(\CONTROL.N_321 ));
    InMux I__6537 (
            .O(N__38606),
            .I(N__38603));
    LocalMux I__6536 (
            .O(N__38603),
            .I(N__38600));
    Odrv12 I__6535 (
            .O(N__38600),
            .I(\CONTROL.N_338 ));
    InMux I__6534 (
            .O(N__38597),
            .I(N__38588));
    InMux I__6533 (
            .O(N__38596),
            .I(N__38588));
    InMux I__6532 (
            .O(N__38595),
            .I(N__38588));
    LocalMux I__6531 (
            .O(N__38588),
            .I(N__38585));
    Span4Mux_v I__6530 (
            .O(N__38585),
            .I(N__38576));
    InMux I__6529 (
            .O(N__38584),
            .I(N__38571));
    InMux I__6528 (
            .O(N__38583),
            .I(N__38571));
    CascadeMux I__6527 (
            .O(N__38582),
            .I(N__38568));
    InMux I__6526 (
            .O(N__38581),
            .I(N__38559));
    InMux I__6525 (
            .O(N__38580),
            .I(N__38559));
    InMux I__6524 (
            .O(N__38579),
            .I(N__38559));
    Span4Mux_h I__6523 (
            .O(N__38576),
            .I(N__38556));
    LocalMux I__6522 (
            .O(N__38571),
            .I(N__38553));
    InMux I__6521 (
            .O(N__38568),
            .I(N__38550));
    InMux I__6520 (
            .O(N__38567),
            .I(N__38545));
    InMux I__6519 (
            .O(N__38566),
            .I(N__38545));
    LocalMux I__6518 (
            .O(N__38559),
            .I(N__38542));
    Odrv4 I__6517 (
            .O(N__38556),
            .I(PROM_ROMDATA_dintern_0ro));
    Odrv4 I__6516 (
            .O(N__38553),
            .I(PROM_ROMDATA_dintern_0ro));
    LocalMux I__6515 (
            .O(N__38550),
            .I(PROM_ROMDATA_dintern_0ro));
    LocalMux I__6514 (
            .O(N__38545),
            .I(PROM_ROMDATA_dintern_0ro));
    Odrv4 I__6513 (
            .O(N__38542),
            .I(PROM_ROMDATA_dintern_0ro));
    CascadeMux I__6512 (
            .O(N__38531),
            .I(PROM_ROMDATA_dintern_0ro_cascade_));
    CascadeMux I__6511 (
            .O(N__38528),
            .I(N__38525));
    InMux I__6510 (
            .O(N__38525),
            .I(N__38522));
    LocalMux I__6509 (
            .O(N__38522),
            .I(N__38519));
    Odrv12 I__6508 (
            .O(N__38519),
            .I(\CONTROL.un1_busState_0_sqmuxa_i_a2_0 ));
    InMux I__6507 (
            .O(N__38516),
            .I(N__38513));
    LocalMux I__6506 (
            .O(N__38513),
            .I(N__38510));
    Span12Mux_s11_v I__6505 (
            .O(N__38510),
            .I(N__38507));
    Odrv12 I__6504 (
            .O(N__38507),
            .I(\CONTROL.N_133_0_1 ));
    CascadeMux I__6503 (
            .O(N__38504),
            .I(PROM_ROMDATA_dintern_3ro_cascade_));
    InMux I__6502 (
            .O(N__38501),
            .I(N__38498));
    LocalMux I__6501 (
            .O(N__38498),
            .I(N__38495));
    Span4Mux_h I__6500 (
            .O(N__38495),
            .I(N__38492));
    Span4Mux_h I__6499 (
            .O(N__38492),
            .I(N__38489));
    Odrv4 I__6498 (
            .O(N__38489),
            .I(\CONTROL.g0_3_i_2_0 ));
    InMux I__6497 (
            .O(N__38486),
            .I(N__38483));
    LocalMux I__6496 (
            .O(N__38483),
            .I(N__38480));
    Odrv12 I__6495 (
            .O(N__38480),
            .I(\CONTROL.g0_2_i_a7Z0Z_3 ));
    InMux I__6494 (
            .O(N__38477),
            .I(N__38474));
    LocalMux I__6493 (
            .O(N__38474),
            .I(\CONTROL.g0_2_i_a7Z0Z_2 ));
    CascadeMux I__6492 (
            .O(N__38471),
            .I(\CONTROL.g0_2_i_2_cascade_ ));
    InMux I__6491 (
            .O(N__38468),
            .I(N__38465));
    LocalMux I__6490 (
            .O(N__38465),
            .I(N__38462));
    Span4Mux_v I__6489 (
            .O(N__38462),
            .I(N__38458));
    CascadeMux I__6488 (
            .O(N__38461),
            .I(N__38455));
    Span4Mux_h I__6487 (
            .O(N__38458),
            .I(N__38452));
    InMux I__6486 (
            .O(N__38455),
            .I(N__38449));
    Odrv4 I__6485 (
            .O(N__38452),
            .I(\CONTROL.addrstack_1_2 ));
    LocalMux I__6484 (
            .O(N__38449),
            .I(\CONTROL.addrstack_1_2 ));
    InMux I__6483 (
            .O(N__38444),
            .I(N__38438));
    InMux I__6482 (
            .O(N__38443),
            .I(N__38432));
    InMux I__6481 (
            .O(N__38442),
            .I(N__38432));
    InMux I__6480 (
            .O(N__38441),
            .I(N__38428));
    LocalMux I__6479 (
            .O(N__38438),
            .I(N__38425));
    InMux I__6478 (
            .O(N__38437),
            .I(N__38422));
    LocalMux I__6477 (
            .O(N__38432),
            .I(N__38419));
    InMux I__6476 (
            .O(N__38431),
            .I(N__38416));
    LocalMux I__6475 (
            .O(N__38428),
            .I(N__38412));
    Span4Mux_v I__6474 (
            .O(N__38425),
            .I(N__38408));
    LocalMux I__6473 (
            .O(N__38422),
            .I(N__38405));
    Span4Mux_v I__6472 (
            .O(N__38419),
            .I(N__38400));
    LocalMux I__6471 (
            .O(N__38416),
            .I(N__38400));
    InMux I__6470 (
            .O(N__38415),
            .I(N__38397));
    Span4Mux_v I__6469 (
            .O(N__38412),
            .I(N__38394));
    InMux I__6468 (
            .O(N__38411),
            .I(N__38391));
    Span4Mux_h I__6467 (
            .O(N__38408),
            .I(N__38384));
    Span4Mux_h I__6466 (
            .O(N__38405),
            .I(N__38384));
    Span4Mux_h I__6465 (
            .O(N__38400),
            .I(N__38384));
    LocalMux I__6464 (
            .O(N__38397),
            .I(\CONTROL.addrstackptrZ0Z_1 ));
    Odrv4 I__6463 (
            .O(N__38394),
            .I(\CONTROL.addrstackptrZ0Z_1 ));
    LocalMux I__6462 (
            .O(N__38391),
            .I(\CONTROL.addrstackptrZ0Z_1 ));
    Odrv4 I__6461 (
            .O(N__38384),
            .I(\CONTROL.addrstackptrZ0Z_1 ));
    CascadeMux I__6460 (
            .O(N__38375),
            .I(\CONTROL.N_5_0_cascade_ ));
    CascadeMux I__6459 (
            .O(N__38372),
            .I(\CONTROL.g0_12_1_cascade_ ));
    CascadeMux I__6458 (
            .O(N__38369),
            .I(N__38366));
    InMux I__6457 (
            .O(N__38366),
            .I(N__38363));
    LocalMux I__6456 (
            .O(N__38363),
            .I(N__38360));
    Span12Mux_h I__6455 (
            .O(N__38360),
            .I(N__38357));
    Odrv12 I__6454 (
            .O(N__38357),
            .I(\CONTROL.addrstackptr_8_2 ));
    CascadeMux I__6453 (
            .O(N__38354),
            .I(controlWord_6_cascade_));
    InMux I__6452 (
            .O(N__38351),
            .I(N__38348));
    LocalMux I__6451 (
            .O(N__38348),
            .I(\CONTROL.N_140_0 ));
    CascadeMux I__6450 (
            .O(N__38345),
            .I(\CONTROL.un1_busState96_1_i_i_a2_1Z0Z_1_cascade_ ));
    InMux I__6449 (
            .O(N__38342),
            .I(N__38339));
    LocalMux I__6448 (
            .O(N__38339),
            .I(\CONTROL.un1_busState96_1_i_i_a2_0Z0Z_1 ));
    CascadeMux I__6447 (
            .O(N__38336),
            .I(\CONTROL.un1_busState96_1_i_iZ0Z_0_cascade_ ));
    CascadeMux I__6446 (
            .O(N__38333),
            .I(controlWord_5_cascade_));
    InMux I__6445 (
            .O(N__38330),
            .I(N__38327));
    LocalMux I__6444 (
            .O(N__38327),
            .I(\CONTROL.N_134_0 ));
    InMux I__6443 (
            .O(N__38324),
            .I(N__38320));
    InMux I__6442 (
            .O(N__38323),
            .I(N__38317));
    LocalMux I__6441 (
            .O(N__38320),
            .I(N__38314));
    LocalMux I__6440 (
            .O(N__38317),
            .I(N__38309));
    Span4Mux_h I__6439 (
            .O(N__38314),
            .I(N__38309));
    Span4Mux_h I__6438 (
            .O(N__38309),
            .I(N__38306));
    Odrv4 I__6437 (
            .O(N__38306),
            .I(\CONTROL.N_327 ));
    InMux I__6436 (
            .O(N__38303),
            .I(N__38300));
    LocalMux I__6435 (
            .O(N__38300),
            .I(N__38297));
    Span4Mux_v I__6434 (
            .O(N__38297),
            .I(N__38294));
    Span4Mux_v I__6433 (
            .O(N__38294),
            .I(N__38291));
    Span4Mux_v I__6432 (
            .O(N__38291),
            .I(N__38288));
    Odrv4 I__6431 (
            .O(N__38288),
            .I(\ALU.status_RNO_2Z0Z_0 ));
    CascadeMux I__6430 (
            .O(N__38285),
            .I(N__38282));
    InMux I__6429 (
            .O(N__38282),
            .I(N__38279));
    LocalMux I__6428 (
            .O(N__38279),
            .I(\ALU.status_e_1_0 ));
    CascadeMux I__6427 (
            .O(N__38276),
            .I(\CONTROL.increment28lto5_1Z0Z_1_cascade_ ));
    InMux I__6426 (
            .O(N__38273),
            .I(N__38269));
    InMux I__6425 (
            .O(N__38272),
            .I(N__38266));
    LocalMux I__6424 (
            .O(N__38269),
            .I(N__38261));
    LocalMux I__6423 (
            .O(N__38266),
            .I(N__38258));
    InMux I__6422 (
            .O(N__38265),
            .I(N__38253));
    InMux I__6421 (
            .O(N__38264),
            .I(N__38253));
    Span4Mux_v I__6420 (
            .O(N__38261),
            .I(N__38250));
    Span4Mux_v I__6419 (
            .O(N__38258),
            .I(N__38244));
    LocalMux I__6418 (
            .O(N__38253),
            .I(N__38241));
    Span4Mux_h I__6417 (
            .O(N__38250),
            .I(N__38238));
    InMux I__6416 (
            .O(N__38249),
            .I(N__38231));
    InMux I__6415 (
            .O(N__38248),
            .I(N__38231));
    InMux I__6414 (
            .O(N__38247),
            .I(N__38231));
    Span4Mux_h I__6413 (
            .O(N__38244),
            .I(N__38226));
    Span4Mux_h I__6412 (
            .O(N__38241),
            .I(N__38226));
    Odrv4 I__6411 (
            .O(N__38238),
            .I(PROM_ROMDATA_dintern_8ro));
    LocalMux I__6410 (
            .O(N__38231),
            .I(PROM_ROMDATA_dintern_8ro));
    Odrv4 I__6409 (
            .O(N__38226),
            .I(PROM_ROMDATA_dintern_8ro));
    CascadeMux I__6408 (
            .O(N__38219),
            .I(\CONTROL.increment28lto5_1_1_2_cascade_ ));
    InMux I__6407 (
            .O(N__38216),
            .I(N__38213));
    LocalMux I__6406 (
            .O(N__38213),
            .I(N__38210));
    Span4Mux_v I__6405 (
            .O(N__38210),
            .I(N__38206));
    InMux I__6404 (
            .O(N__38209),
            .I(N__38201));
    Span4Mux_h I__6403 (
            .O(N__38206),
            .I(N__38198));
    InMux I__6402 (
            .O(N__38205),
            .I(N__38193));
    InMux I__6401 (
            .O(N__38204),
            .I(N__38193));
    LocalMux I__6400 (
            .O(N__38201),
            .I(PROM_ROMDATA_dintern_7ro));
    Odrv4 I__6399 (
            .O(N__38198),
            .I(PROM_ROMDATA_dintern_7ro));
    LocalMux I__6398 (
            .O(N__38193),
            .I(PROM_ROMDATA_dintern_7ro));
    InMux I__6397 (
            .O(N__38186),
            .I(N__38181));
    InMux I__6396 (
            .O(N__38185),
            .I(N__38178));
    InMux I__6395 (
            .O(N__38184),
            .I(N__38175));
    LocalMux I__6394 (
            .O(N__38181),
            .I(N__38172));
    LocalMux I__6393 (
            .O(N__38178),
            .I(N__38167));
    LocalMux I__6392 (
            .O(N__38175),
            .I(N__38167));
    Span4Mux_h I__6391 (
            .O(N__38172),
            .I(N__38164));
    Span4Mux_v I__6390 (
            .O(N__38167),
            .I(N__38161));
    Span4Mux_h I__6389 (
            .O(N__38164),
            .I(N__38157));
    Span4Mux_h I__6388 (
            .O(N__38161),
            .I(N__38154));
    InMux I__6387 (
            .O(N__38160),
            .I(N__38151));
    Odrv4 I__6386 (
            .O(N__38157),
            .I(\CONTROL.increment28lto5_1Z0Z_2 ));
    Odrv4 I__6385 (
            .O(N__38154),
            .I(\CONTROL.increment28lto5_1Z0Z_2 ));
    LocalMux I__6384 (
            .O(N__38151),
            .I(\CONTROL.increment28lto5_1Z0Z_2 ));
    CEMux I__6383 (
            .O(N__38144),
            .I(N__38141));
    LocalMux I__6382 (
            .O(N__38141),
            .I(N__38137));
    CascadeMux I__6381 (
            .O(N__38140),
            .I(N__38134));
    Span4Mux_v I__6380 (
            .O(N__38137),
            .I(N__38131));
    InMux I__6379 (
            .O(N__38134),
            .I(N__38128));
    Span4Mux_h I__6378 (
            .O(N__38131),
            .I(N__38122));
    LocalMux I__6377 (
            .O(N__38128),
            .I(N__38119));
    InMux I__6376 (
            .O(N__38127),
            .I(N__38116));
    CEMux I__6375 (
            .O(N__38126),
            .I(N__38113));
    CEMux I__6374 (
            .O(N__38125),
            .I(N__38110));
    Sp12to4 I__6373 (
            .O(N__38122),
            .I(N__38105));
    Span12Mux_v I__6372 (
            .O(N__38119),
            .I(N__38105));
    LocalMux I__6371 (
            .O(N__38116),
            .I(N__38102));
    LocalMux I__6370 (
            .O(N__38113),
            .I(\CONTROL.N_48_0 ));
    LocalMux I__6369 (
            .O(N__38110),
            .I(\CONTROL.N_48_0 ));
    Odrv12 I__6368 (
            .O(N__38105),
            .I(\CONTROL.N_48_0 ));
    Odrv4 I__6367 (
            .O(N__38102),
            .I(\CONTROL.N_48_0 ));
    CascadeMux I__6366 (
            .O(N__38093),
            .I(\ALU.N_1200_cascade_ ));
    InMux I__6365 (
            .O(N__38090),
            .I(N__38087));
    LocalMux I__6364 (
            .O(N__38087),
            .I(\ALU.N_1248 ));
    CascadeMux I__6363 (
            .O(N__38084),
            .I(\ALU.d_RNIGMEO4Z0Z_3_cascade_ ));
    InMux I__6362 (
            .O(N__38081),
            .I(N__38078));
    LocalMux I__6361 (
            .O(N__38078),
            .I(N__38075));
    Span4Mux_v I__6360 (
            .O(N__38075),
            .I(N__38072));
    Span4Mux_h I__6359 (
            .O(N__38072),
            .I(N__38069));
    Odrv4 I__6358 (
            .O(N__38069),
            .I(\ALU.combOperand2_d_bmZ0Z_3 ));
    InMux I__6357 (
            .O(N__38066),
            .I(N__38062));
    InMux I__6356 (
            .O(N__38065),
            .I(N__38059));
    LocalMux I__6355 (
            .O(N__38062),
            .I(N__38054));
    LocalMux I__6354 (
            .O(N__38059),
            .I(N__38051));
    InMux I__6353 (
            .O(N__38058),
            .I(N__38046));
    InMux I__6352 (
            .O(N__38057),
            .I(N__38046));
    Span4Mux_v I__6351 (
            .O(N__38054),
            .I(N__38043));
    Span4Mux_v I__6350 (
            .O(N__38051),
            .I(N__38040));
    LocalMux I__6349 (
            .O(N__38046),
            .I(N__38037));
    Span4Mux_h I__6348 (
            .O(N__38043),
            .I(N__38032));
    Span4Mux_h I__6347 (
            .O(N__38040),
            .I(N__38032));
    Odrv12 I__6346 (
            .O(N__38037),
            .I(\ALU.d_RNI2CUG6Z0Z_3 ));
    Odrv4 I__6345 (
            .O(N__38032),
            .I(\ALU.d_RNI2CUG6Z0Z_3 ));
    InMux I__6344 (
            .O(N__38027),
            .I(N__38024));
    LocalMux I__6343 (
            .O(N__38024),
            .I(N__38021));
    Span4Mux_v I__6342 (
            .O(N__38021),
            .I(N__38018));
    Span4Mux_v I__6341 (
            .O(N__38018),
            .I(N__38015));
    Span4Mux_v I__6340 (
            .O(N__38015),
            .I(N__38012));
    Span4Mux_v I__6339 (
            .O(N__38012),
            .I(N__38009));
    Span4Mux_h I__6338 (
            .O(N__38009),
            .I(N__38006));
    Span4Mux_h I__6337 (
            .O(N__38006),
            .I(N__38003));
    Span4Mux_h I__6336 (
            .O(N__38003),
            .I(N__38000));
    Span4Mux_h I__6335 (
            .O(N__38000),
            .I(N__37997));
    Odrv4 I__6334 (
            .O(N__37997),
            .I(gpuOut_c_4));
    InMux I__6333 (
            .O(N__37994),
            .I(N__37990));
    InMux I__6332 (
            .O(N__37993),
            .I(N__37987));
    LocalMux I__6331 (
            .O(N__37990),
            .I(N__37984));
    LocalMux I__6330 (
            .O(N__37987),
            .I(N__37981));
    Span4Mux_h I__6329 (
            .O(N__37984),
            .I(N__37978));
    Span4Mux_v I__6328 (
            .O(N__37981),
            .I(N__37973));
    Span4Mux_v I__6327 (
            .O(N__37978),
            .I(N__37973));
    Odrv4 I__6326 (
            .O(N__37973),
            .I(\CONTROL.N_165 ));
    CascadeMux I__6325 (
            .O(N__37970),
            .I(N__37967));
    InMux I__6324 (
            .O(N__37967),
            .I(N__37964));
    LocalMux I__6323 (
            .O(N__37964),
            .I(N__37961));
    Span4Mux_v I__6322 (
            .O(N__37961),
            .I(N__37957));
    InMux I__6321 (
            .O(N__37960),
            .I(N__37954));
    Span4Mux_v I__6320 (
            .O(N__37957),
            .I(N__37951));
    LocalMux I__6319 (
            .O(N__37954),
            .I(N__37948));
    Sp12to4 I__6318 (
            .O(N__37951),
            .I(N__37945));
    Span4Mux_h I__6317 (
            .O(N__37948),
            .I(N__37942));
    Span12Mux_h I__6316 (
            .O(N__37945),
            .I(N__37938));
    Span4Mux_h I__6315 (
            .O(N__37942),
            .I(N__37935));
    InMux I__6314 (
            .O(N__37941),
            .I(N__37932));
    Odrv12 I__6313 (
            .O(N__37938),
            .I(h_9));
    Odrv4 I__6312 (
            .O(N__37935),
            .I(h_9));
    LocalMux I__6311 (
            .O(N__37932),
            .I(h_9));
    InMux I__6310 (
            .O(N__37925),
            .I(N__37922));
    LocalMux I__6309 (
            .O(N__37922),
            .I(N__37919));
    Odrv4 I__6308 (
            .O(N__37919),
            .I(\ALU.e_RNICGJMZ0Z_9 ));
    InMux I__6307 (
            .O(N__37916),
            .I(N__37913));
    LocalMux I__6306 (
            .O(N__37913),
            .I(\ALU.d_RNIKKNJZ0Z_9 ));
    CascadeMux I__6305 (
            .O(N__37910),
            .I(\ALU.operand2_7_ns_1_9_cascade_ ));
    InMux I__6304 (
            .O(N__37907),
            .I(N__37904));
    LocalMux I__6303 (
            .O(N__37904),
            .I(\ALU.b_RNIG8BVZ0Z_9 ));
    CascadeMux I__6302 (
            .O(N__37901),
            .I(\ALU.operand2_9_cascade_ ));
    InMux I__6301 (
            .O(N__37898),
            .I(N__37895));
    LocalMux I__6300 (
            .O(N__37895),
            .I(\ALU.e_RNI933SZ0Z_0 ));
    CascadeMux I__6299 (
            .O(N__37892),
            .I(\ALU.c_RNIDFF01Z0Z_0_cascade_ ));
    InMux I__6298 (
            .O(N__37889),
            .I(N__37886));
    LocalMux I__6297 (
            .O(N__37886),
            .I(\ALU.d_RNI0G5DZ0Z_0 ));
    CascadeMux I__6296 (
            .O(N__37883),
            .I(\ALU.b_RNIS3POZ0Z_0_cascade_ ));
    InMux I__6295 (
            .O(N__37880),
            .I(N__37877));
    LocalMux I__6294 (
            .O(N__37877),
            .I(\ALU.operand2_7_ns_1_0 ));
    InMux I__6293 (
            .O(N__37874),
            .I(N__37871));
    LocalMux I__6292 (
            .O(N__37871),
            .I(N__37867));
    InMux I__6291 (
            .O(N__37870),
            .I(N__37864));
    Span4Mux_v I__6290 (
            .O(N__37867),
            .I(N__37861));
    LocalMux I__6289 (
            .O(N__37864),
            .I(N__37858));
    Span4Mux_v I__6288 (
            .O(N__37861),
            .I(N__37853));
    Span4Mux_h I__6287 (
            .O(N__37858),
            .I(N__37853));
    Odrv4 I__6286 (
            .O(N__37853),
            .I(\ALU.operand2_0 ));
    InMux I__6285 (
            .O(N__37850),
            .I(N__37847));
    LocalMux I__6284 (
            .O(N__37847),
            .I(N__37844));
    Span4Mux_h I__6283 (
            .O(N__37844),
            .I(N__37840));
    InMux I__6282 (
            .O(N__37843),
            .I(N__37837));
    Span4Mux_v I__6281 (
            .O(N__37840),
            .I(N__37832));
    LocalMux I__6280 (
            .O(N__37837),
            .I(N__37832));
    Odrv4 I__6279 (
            .O(N__37832),
            .I(\ALU.dZ0Z_3 ));
    CascadeMux I__6278 (
            .O(N__37829),
            .I(\ALU.operand2_6_ns_1_3_cascade_ ));
    InMux I__6277 (
            .O(N__37826),
            .I(N__37823));
    LocalMux I__6276 (
            .O(N__37823),
            .I(N__37819));
    InMux I__6275 (
            .O(N__37822),
            .I(N__37816));
    Span4Mux_h I__6274 (
            .O(N__37819),
            .I(N__37813));
    LocalMux I__6273 (
            .O(N__37816),
            .I(N__37810));
    Span4Mux_v I__6272 (
            .O(N__37813),
            .I(N__37807));
    Odrv12 I__6271 (
            .O(N__37810),
            .I(\ALU.aZ0Z_3 ));
    Odrv4 I__6270 (
            .O(N__37807),
            .I(\ALU.aZ0Z_3 ));
    CascadeMux I__6269 (
            .O(N__37802),
            .I(N__37798));
    CascadeMux I__6268 (
            .O(N__37801),
            .I(N__37795));
    InMux I__6267 (
            .O(N__37798),
            .I(N__37792));
    InMux I__6266 (
            .O(N__37795),
            .I(N__37789));
    LocalMux I__6265 (
            .O(N__37792),
            .I(N__37786));
    LocalMux I__6264 (
            .O(N__37789),
            .I(N__37783));
    Span4Mux_h I__6263 (
            .O(N__37786),
            .I(N__37780));
    Span4Mux_v I__6262 (
            .O(N__37783),
            .I(N__37777));
    Span4Mux_h I__6261 (
            .O(N__37780),
            .I(N__37774));
    Odrv4 I__6260 (
            .O(N__37777),
            .I(\ALU.eZ0Z_3 ));
    Odrv4 I__6259 (
            .O(N__37774),
            .I(\ALU.eZ0Z_3 ));
    InMux I__6258 (
            .O(N__37769),
            .I(N__37765));
    InMux I__6257 (
            .O(N__37768),
            .I(N__37762));
    LocalMux I__6256 (
            .O(N__37765),
            .I(N__37759));
    LocalMux I__6255 (
            .O(N__37762),
            .I(N__37756));
    Span4Mux_v I__6254 (
            .O(N__37759),
            .I(N__37753));
    Sp12to4 I__6253 (
            .O(N__37756),
            .I(N__37750));
    Odrv4 I__6252 (
            .O(N__37753),
            .I(\ALU.cZ0Z_3 ));
    Odrv12 I__6251 (
            .O(N__37750),
            .I(\ALU.cZ0Z_3 ));
    InMux I__6250 (
            .O(N__37745),
            .I(N__37742));
    LocalMux I__6249 (
            .O(N__37742),
            .I(N__37738));
    InMux I__6248 (
            .O(N__37741),
            .I(N__37734));
    Span4Mux_v I__6247 (
            .O(N__37738),
            .I(N__37731));
    InMux I__6246 (
            .O(N__37737),
            .I(N__37728));
    LocalMux I__6245 (
            .O(N__37734),
            .I(N__37725));
    Span4Mux_v I__6244 (
            .O(N__37731),
            .I(N__37722));
    LocalMux I__6243 (
            .O(N__37728),
            .I(N__37719));
    Span4Mux_v I__6242 (
            .O(N__37725),
            .I(N__37716));
    Span4Mux_v I__6241 (
            .O(N__37722),
            .I(N__37713));
    Span4Mux_v I__6240 (
            .O(N__37719),
            .I(N__37710));
    Span4Mux_h I__6239 (
            .O(N__37716),
            .I(N__37707));
    Span4Mux_h I__6238 (
            .O(N__37713),
            .I(N__37702));
    Span4Mux_v I__6237 (
            .O(N__37710),
            .I(N__37702));
    Span4Mux_v I__6236 (
            .O(N__37707),
            .I(N__37699));
    Odrv4 I__6235 (
            .O(N__37702),
            .I(g_3));
    Odrv4 I__6234 (
            .O(N__37699),
            .I(g_3));
    CascadeMux I__6233 (
            .O(N__37694),
            .I(\ALU.operand2_3_ns_1_3_cascade_ ));
    CascadeMux I__6232 (
            .O(N__37691),
            .I(\ALU.a_15_m2_d_d_ns_1_0_0_cascade_ ));
    IoInMux I__6231 (
            .O(N__37688),
            .I(N__37685));
    LocalMux I__6230 (
            .O(N__37685),
            .I(N__37681));
    IoInMux I__6229 (
            .O(N__37684),
            .I(N__37678));
    IoSpan4Mux I__6228 (
            .O(N__37681),
            .I(N__37675));
    LocalMux I__6227 (
            .O(N__37678),
            .I(N__37672));
    IoSpan4Mux I__6226 (
            .O(N__37675),
            .I(N__37669));
    IoSpan4Mux I__6225 (
            .O(N__37672),
            .I(N__37666));
    Sp12to4 I__6224 (
            .O(N__37669),
            .I(N__37663));
    Span4Mux_s0_h I__6223 (
            .O(N__37666),
            .I(N__37660));
    Span12Mux_s7_h I__6222 (
            .O(N__37663),
            .I(N__37656));
    Sp12to4 I__6221 (
            .O(N__37660),
            .I(N__37653));
    InMux I__6220 (
            .O(N__37659),
            .I(N__37650));
    Span12Mux_h I__6219 (
            .O(N__37656),
            .I(N__37645));
    Span12Mux_h I__6218 (
            .O(N__37653),
            .I(N__37645));
    LocalMux I__6217 (
            .O(N__37650),
            .I(N__37642));
    Odrv12 I__6216 (
            .O(N__37645),
            .I(bus_0));
    Odrv12 I__6215 (
            .O(N__37642),
            .I(bus_0));
    InMux I__6214 (
            .O(N__37637),
            .I(N__37633));
    InMux I__6213 (
            .O(N__37636),
            .I(N__37630));
    LocalMux I__6212 (
            .O(N__37633),
            .I(N__37627));
    LocalMux I__6211 (
            .O(N__37630),
            .I(N__37624));
    Span4Mux_v I__6210 (
            .O(N__37627),
            .I(N__37621));
    Span4Mux_v I__6209 (
            .O(N__37624),
            .I(N__37618));
    Span4Mux_h I__6208 (
            .O(N__37621),
            .I(N__37615));
    Span4Mux_h I__6207 (
            .O(N__37618),
            .I(N__37612));
    Span4Mux_v I__6206 (
            .O(N__37615),
            .I(N__37609));
    Odrv4 I__6205 (
            .O(N__37612),
            .I(\ALU.lshift62 ));
    Odrv4 I__6204 (
            .O(N__37609),
            .I(\ALU.lshift62 ));
    CascadeMux I__6203 (
            .O(N__37604),
            .I(\ALU.d_RNI4D6E01Z0Z_0_cascade_ ));
    CascadeMux I__6202 (
            .O(N__37601),
            .I(\ALU.d_RNIQQ9O83Z0Z_0_cascade_ ));
    InMux I__6201 (
            .O(N__37598),
            .I(N__37595));
    LocalMux I__6200 (
            .O(N__37595),
            .I(\ALU.d_RNI4HL061Z0Z_0 ));
    CascadeMux I__6199 (
            .O(N__37592),
            .I(\ALU.d_RNINUGCF4Z0Z_0_cascade_ ));
    CascadeMux I__6198 (
            .O(N__37589),
            .I(N__37586));
    InMux I__6197 (
            .O(N__37586),
            .I(N__37583));
    LocalMux I__6196 (
            .O(N__37583),
            .I(N__37580));
    Span4Mux_h I__6195 (
            .O(N__37580),
            .I(N__37576));
    InMux I__6194 (
            .O(N__37579),
            .I(N__37573));
    Span4Mux_h I__6193 (
            .O(N__37576),
            .I(N__37570));
    LocalMux I__6192 (
            .O(N__37573),
            .I(\ALU.aZ0Z_0 ));
    Odrv4 I__6191 (
            .O(N__37570),
            .I(\ALU.aZ0Z_0 ));
    InMux I__6190 (
            .O(N__37565),
            .I(N__37562));
    LocalMux I__6189 (
            .O(N__37562),
            .I(N__37558));
    CascadeMux I__6188 (
            .O(N__37561),
            .I(N__37555));
    Span4Mux_v I__6187 (
            .O(N__37558),
            .I(N__37552));
    InMux I__6186 (
            .O(N__37555),
            .I(N__37549));
    Span4Mux_h I__6185 (
            .O(N__37552),
            .I(N__37543));
    LocalMux I__6184 (
            .O(N__37549),
            .I(N__37543));
    InMux I__6183 (
            .O(N__37548),
            .I(N__37540));
    Span4Mux_h I__6182 (
            .O(N__37543),
            .I(N__37537));
    LocalMux I__6181 (
            .O(N__37540),
            .I(h_0));
    Odrv4 I__6180 (
            .O(N__37537),
            .I(h_0));
    InMux I__6179 (
            .O(N__37532),
            .I(N__37528));
    InMux I__6178 (
            .O(N__37531),
            .I(N__37525));
    LocalMux I__6177 (
            .O(N__37528),
            .I(\ALU.a_15_am_snZ0Z_11 ));
    LocalMux I__6176 (
            .O(N__37525),
            .I(\ALU.a_15_am_snZ0Z_11 ));
    InMux I__6175 (
            .O(N__37520),
            .I(N__37517));
    LocalMux I__6174 (
            .O(N__37517),
            .I(N__37513));
    CascadeMux I__6173 (
            .O(N__37516),
            .I(N__37509));
    Span4Mux_v I__6172 (
            .O(N__37513),
            .I(N__37506));
    InMux I__6171 (
            .O(N__37512),
            .I(N__37503));
    InMux I__6170 (
            .O(N__37509),
            .I(N__37500));
    Span4Mux_h I__6169 (
            .O(N__37506),
            .I(N__37495));
    LocalMux I__6168 (
            .O(N__37503),
            .I(N__37495));
    LocalMux I__6167 (
            .O(N__37500),
            .I(N__37492));
    Span4Mux_h I__6166 (
            .O(N__37495),
            .I(N__37487));
    Span4Mux_h I__6165 (
            .O(N__37492),
            .I(N__37487));
    Span4Mux_v I__6164 (
            .O(N__37487),
            .I(N__37484));
    Span4Mux_h I__6163 (
            .O(N__37484),
            .I(N__37481));
    Odrv4 I__6162 (
            .O(N__37481),
            .I(h_1));
    InMux I__6161 (
            .O(N__37478),
            .I(N__37475));
    LocalMux I__6160 (
            .O(N__37475),
            .I(N__37472));
    Span4Mux_v I__6159 (
            .O(N__37472),
            .I(N__37469));
    Odrv4 I__6158 (
            .O(N__37469),
            .I(\ALU.mult_6 ));
    CascadeMux I__6157 (
            .O(N__37466),
            .I(\ALU.mult_489_c_RNIGEUL1AZ0_cascade_ ));
    InMux I__6156 (
            .O(N__37463),
            .I(N__37460));
    LocalMux I__6155 (
            .O(N__37460),
            .I(\ALU.mult_489_c_RNIGEUL1AZ0 ));
    CascadeMux I__6154 (
            .O(N__37457),
            .I(\ALU.mult_489_c_RNIPGBQMCZ0Z_0_cascade_ ));
    InMux I__6153 (
            .O(N__37454),
            .I(N__37451));
    LocalMux I__6152 (
            .O(N__37451),
            .I(\ALU.mult_489_c_RNIPGBQMCZ0 ));
    CascadeMux I__6151 (
            .O(N__37448),
            .I(\ALU.mult_489_c_RNI1J3GCUZ0_cascade_ ));
    CascadeMux I__6150 (
            .O(N__37445),
            .I(N__37442));
    InMux I__6149 (
            .O(N__37442),
            .I(N__37439));
    LocalMux I__6148 (
            .O(N__37439),
            .I(N__37435));
    InMux I__6147 (
            .O(N__37438),
            .I(N__37431));
    Span4Mux_h I__6146 (
            .O(N__37435),
            .I(N__37428));
    InMux I__6145 (
            .O(N__37434),
            .I(N__37425));
    LocalMux I__6144 (
            .O(N__37431),
            .I(N__37422));
    Span4Mux_v I__6143 (
            .O(N__37428),
            .I(N__37417));
    LocalMux I__6142 (
            .O(N__37425),
            .I(N__37417));
    Span4Mux_v I__6141 (
            .O(N__37422),
            .I(N__37414));
    Span4Mux_h I__6140 (
            .O(N__37417),
            .I(N__37411));
    Sp12to4 I__6139 (
            .O(N__37414),
            .I(N__37408));
    Odrv4 I__6138 (
            .O(N__37411),
            .I(h_6));
    Odrv12 I__6137 (
            .O(N__37408),
            .I(h_6));
    InMux I__6136 (
            .O(N__37403),
            .I(N__37400));
    LocalMux I__6135 (
            .O(N__37400),
            .I(N__37397));
    Span4Mux_v I__6134 (
            .O(N__37397),
            .I(N__37394));
    Span4Mux_h I__6133 (
            .O(N__37394),
            .I(N__37391));
    Span4Mux_h I__6132 (
            .O(N__37391),
            .I(N__37388));
    Odrv4 I__6131 (
            .O(N__37388),
            .I(\ALU.status_17_I_39_c_RNOZ0 ));
    CascadeMux I__6130 (
            .O(N__37385),
            .I(N__37382));
    InMux I__6129 (
            .O(N__37382),
            .I(N__37379));
    LocalMux I__6128 (
            .O(N__37379),
            .I(N__37376));
    Odrv12 I__6127 (
            .O(N__37376),
            .I(\ALU.mult_365_c_RNOZ0Z_0 ));
    InMux I__6126 (
            .O(N__37373),
            .I(N__37370));
    LocalMux I__6125 (
            .O(N__37370),
            .I(N__37366));
    InMux I__6124 (
            .O(N__37369),
            .I(N__37363));
    Odrv12 I__6123 (
            .O(N__37366),
            .I(\ALU.N_572 ));
    LocalMux I__6122 (
            .O(N__37363),
            .I(\ALU.N_572 ));
    IoInMux I__6121 (
            .O(N__37358),
            .I(N__37355));
    LocalMux I__6120 (
            .O(N__37355),
            .I(N__37351));
    IoInMux I__6119 (
            .O(N__37354),
            .I(N__37348));
    IoSpan4Mux I__6118 (
            .O(N__37351),
            .I(N__37345));
    LocalMux I__6117 (
            .O(N__37348),
            .I(N__37342));
    Sp12to4 I__6116 (
            .O(N__37345),
            .I(N__37338));
    IoSpan4Mux I__6115 (
            .O(N__37342),
            .I(N__37335));
    InMux I__6114 (
            .O(N__37341),
            .I(N__37332));
    Span12Mux_s7_h I__6113 (
            .O(N__37338),
            .I(N__37329));
    Sp12to4 I__6112 (
            .O(N__37335),
            .I(N__37326));
    LocalMux I__6111 (
            .O(N__37332),
            .I(N__37323));
    Span12Mux_h I__6110 (
            .O(N__37329),
            .I(N__37318));
    Span12Mux_h I__6109 (
            .O(N__37326),
            .I(N__37318));
    Span4Mux_h I__6108 (
            .O(N__37323),
            .I(N__37315));
    Span12Mux_v I__6107 (
            .O(N__37318),
            .I(N__37312));
    Span4Mux_v I__6106 (
            .O(N__37315),
            .I(N__37309));
    Odrv12 I__6105 (
            .O(N__37312),
            .I(bus_11));
    Odrv4 I__6104 (
            .O(N__37309),
            .I(bus_11));
    InMux I__6103 (
            .O(N__37304),
            .I(N__37301));
    LocalMux I__6102 (
            .O(N__37301),
            .I(N__37298));
    Odrv4 I__6101 (
            .O(N__37298),
            .I(\ALU.mult_11 ));
    CascadeMux I__6100 (
            .O(N__37295),
            .I(\ALU.mult_552_c_RNI70R9DAZ0_cascade_ ));
    InMux I__6099 (
            .O(N__37292),
            .I(N__37289));
    LocalMux I__6098 (
            .O(N__37289),
            .I(\ALU.rshift_11 ));
    CascadeMux I__6097 (
            .O(N__37286),
            .I(N__37282));
    InMux I__6096 (
            .O(N__37285),
            .I(N__37277));
    InMux I__6095 (
            .O(N__37282),
            .I(N__37277));
    LocalMux I__6094 (
            .O(N__37277),
            .I(\ALU.a_15_am_rn_0_11 ));
    InMux I__6093 (
            .O(N__37274),
            .I(N__37271));
    LocalMux I__6092 (
            .O(N__37271),
            .I(\ALU.mult_552_c_RNI70R9DAZ0 ));
    CascadeMux I__6091 (
            .O(N__37268),
            .I(\ALU.mult_552_c_RNIOT7VLFZ0_cascade_ ));
    CascadeMux I__6090 (
            .O(N__37265),
            .I(N__37262));
    InMux I__6089 (
            .O(N__37262),
            .I(N__37256));
    InMux I__6088 (
            .O(N__37261),
            .I(N__37256));
    LocalMux I__6087 (
            .O(N__37256),
            .I(N__37253));
    Span4Mux_v I__6086 (
            .O(N__37253),
            .I(N__37250));
    Span4Mux_h I__6085 (
            .O(N__37250),
            .I(N__37247));
    Odrv4 I__6084 (
            .O(N__37247),
            .I(\ALU.aZ0Z_11 ));
    CascadeMux I__6083 (
            .O(N__37244),
            .I(\ALU.a_15_m3_sZ0Z_13_cascade_ ));
    CascadeMux I__6082 (
            .O(N__37241),
            .I(\ALU.a32Z0Z_0_cascade_ ));
    InMux I__6081 (
            .O(N__37238),
            .I(N__37235));
    LocalMux I__6080 (
            .O(N__37235),
            .I(N__37231));
    InMux I__6079 (
            .O(N__37234),
            .I(N__37228));
    Span4Mux_h I__6078 (
            .O(N__37231),
            .I(N__37225));
    LocalMux I__6077 (
            .O(N__37228),
            .I(N__37222));
    Span4Mux_v I__6076 (
            .O(N__37225),
            .I(N__37217));
    Span4Mux_h I__6075 (
            .O(N__37222),
            .I(N__37217));
    Span4Mux_h I__6074 (
            .O(N__37217),
            .I(N__37214));
    Span4Mux_v I__6073 (
            .O(N__37214),
            .I(N__37211));
    Odrv4 I__6072 (
            .O(N__37211),
            .I(\ALU.aZ0Z_1 ));
    CascadeMux I__6071 (
            .O(N__37208),
            .I(\ALU.d_RNICUA7B5Z0Z_0_cascade_ ));
    CascadeMux I__6070 (
            .O(N__37205),
            .I(N__37202));
    InMux I__6069 (
            .O(N__37202),
            .I(N__37199));
    LocalMux I__6068 (
            .O(N__37199),
            .I(N__37196));
    Odrv12 I__6067 (
            .O(N__37196),
            .I(\ALU.d_RNIL3JT71Z0Z_0 ));
    InMux I__6066 (
            .O(N__37193),
            .I(N__37190));
    LocalMux I__6065 (
            .O(N__37190),
            .I(N__37187));
    Span4Mux_h I__6064 (
            .O(N__37187),
            .I(N__37184));
    Odrv4 I__6063 (
            .O(N__37184),
            .I(\ALU.N_556 ));
    CascadeMux I__6062 (
            .O(N__37181),
            .I(\ALU.N_556_cascade_ ));
    InMux I__6061 (
            .O(N__37178),
            .I(N__37175));
    LocalMux I__6060 (
            .O(N__37175),
            .I(\ALU.d_RNI3MGBH1Z0Z_1 ));
    CascadeMux I__6059 (
            .O(N__37172),
            .I(N__37169));
    InMux I__6058 (
            .O(N__37169),
            .I(N__37166));
    LocalMux I__6057 (
            .O(N__37166),
            .I(\ALU.mult_25_11 ));
    InMux I__6056 (
            .O(N__37163),
            .I(\ALU.mult_29_c10 ));
    InMux I__6055 (
            .O(N__37160),
            .I(\ALU.mult_29_c11 ));
    InMux I__6054 (
            .O(N__37157),
            .I(N__37154));
    LocalMux I__6053 (
            .O(N__37154),
            .I(\ALU.mult_25_13 ));
    InMux I__6052 (
            .O(N__37151),
            .I(\ALU.mult_29_c12 ));
    InMux I__6051 (
            .O(N__37148),
            .I(N__37145));
    LocalMux I__6050 (
            .O(N__37145),
            .I(\ALU.mult_25_14 ));
    InMux I__6049 (
            .O(N__37142),
            .I(\ALU.mult_29_c13 ));
    InMux I__6048 (
            .O(N__37139),
            .I(N__37136));
    LocalMux I__6047 (
            .O(N__37136),
            .I(\ALU.mult_516_c_RNI98SKDCZ0 ));
    InMux I__6046 (
            .O(N__37133),
            .I(\ALU.mult_29_c14 ));
    InMux I__6045 (
            .O(N__37130),
            .I(N__37127));
    LocalMux I__6044 (
            .O(N__37127),
            .I(N__37124));
    Span4Mux_v I__6043 (
            .O(N__37124),
            .I(N__37121));
    Span4Mux_h I__6042 (
            .O(N__37121),
            .I(N__37117));
    InMux I__6041 (
            .O(N__37120),
            .I(N__37114));
    Span4Mux_h I__6040 (
            .O(N__37117),
            .I(N__37107));
    LocalMux I__6039 (
            .O(N__37114),
            .I(N__37107));
    InMux I__6038 (
            .O(N__37113),
            .I(N__37104));
    InMux I__6037 (
            .O(N__37112),
            .I(N__37101));
    Odrv4 I__6036 (
            .O(N__37107),
            .I(bus_0_10));
    LocalMux I__6035 (
            .O(N__37104),
            .I(bus_0_10));
    LocalMux I__6034 (
            .O(N__37101),
            .I(bus_0_10));
    InMux I__6033 (
            .O(N__37094),
            .I(N__37091));
    LocalMux I__6032 (
            .O(N__37091),
            .I(\ALU.mult_10 ));
    CascadeMux I__6031 (
            .O(N__37088),
            .I(\ALU.mult_549_c_RNIB6TIDGZ0_cascade_ ));
    InMux I__6030 (
            .O(N__37085),
            .I(N__37082));
    LocalMux I__6029 (
            .O(N__37082),
            .I(\ALU.a_15_am_1_10 ));
    CascadeMux I__6028 (
            .O(N__37079),
            .I(\ALU.mult_549_c_RNIE7260OZ0_cascade_ ));
    InMux I__6027 (
            .O(N__37076),
            .I(N__37072));
    InMux I__6026 (
            .O(N__37075),
            .I(N__37069));
    LocalMux I__6025 (
            .O(N__37072),
            .I(N__37064));
    LocalMux I__6024 (
            .O(N__37069),
            .I(N__37064));
    Span4Mux_v I__6023 (
            .O(N__37064),
            .I(N__37061));
    Span4Mux_v I__6022 (
            .O(N__37061),
            .I(N__37058));
    Sp12to4 I__6021 (
            .O(N__37058),
            .I(N__37055));
    Odrv12 I__6020 (
            .O(N__37055),
            .I(\ALU.aZ0Z_10 ));
    InMux I__6019 (
            .O(N__37052),
            .I(N__37049));
    LocalMux I__6018 (
            .O(N__37049),
            .I(N__37046));
    Span4Mux_h I__6017 (
            .O(N__37046),
            .I(N__37043));
    Odrv4 I__6016 (
            .O(N__37043),
            .I(\ALU.mult_365_c_RNOZ0 ));
    InMux I__6015 (
            .O(N__37040),
            .I(N__37037));
    LocalMux I__6014 (
            .O(N__37037),
            .I(N__37034));
    Span4Mux_h I__6013 (
            .O(N__37034),
            .I(N__37031));
    Odrv4 I__6012 (
            .O(N__37031),
            .I(\ALU.c_RNIF6GEF1Z0Z_12 ));
    CascadeMux I__6011 (
            .O(N__37028),
            .I(N__37025));
    InMux I__6010 (
            .O(N__37025),
            .I(N__37022));
    LocalMux I__6009 (
            .O(N__37022),
            .I(N__37019));
    Odrv4 I__6008 (
            .O(N__37019),
            .I(\ALU.c_RNINUT6PZ0Z_13 ));
    InMux I__6007 (
            .O(N__37016),
            .I(\ALU.mult_13_c13 ));
    InMux I__6006 (
            .O(N__37013),
            .I(N__37010));
    LocalMux I__6005 (
            .O(N__37010),
            .I(N__37007));
    Odrv4 I__6004 (
            .O(N__37007),
            .I(\ALU.c_RNIS83N71Z0Z_12 ));
    InMux I__6003 (
            .O(N__37004),
            .I(\ALU.mult_13_c14 ));
    CascadeMux I__6002 (
            .O(N__37001),
            .I(N__36998));
    InMux I__6001 (
            .O(N__36998),
            .I(N__36995));
    LocalMux I__6000 (
            .O(N__36995),
            .I(N__36992));
    Span4Mux_h I__5999 (
            .O(N__36992),
            .I(N__36989));
    Odrv4 I__5998 (
            .O(N__36989),
            .I(\ALU.d_RNIL4PC21Z0Z_6 ));
    InMux I__5997 (
            .O(N__36986),
            .I(N__36983));
    LocalMux I__5996 (
            .O(N__36983),
            .I(\ALU.mult_5_5 ));
    InMux I__5995 (
            .O(N__36980),
            .I(N__36977));
    LocalMux I__5994 (
            .O(N__36977),
            .I(N__36974));
    Span4Mux_h I__5993 (
            .O(N__36974),
            .I(N__36971));
    Odrv4 I__5992 (
            .O(N__36971),
            .I(\ALU.mult_9_9 ));
    CascadeMux I__5991 (
            .O(N__36968),
            .I(N__36965));
    InMux I__5990 (
            .O(N__36965),
            .I(N__36962));
    LocalMux I__5989 (
            .O(N__36962),
            .I(\ALU.mult_25_9 ));
    InMux I__5988 (
            .O(N__36959),
            .I(\ALU.mult_29_c8 ));
    InMux I__5987 (
            .O(N__36956),
            .I(\ALU.mult_29_c9 ));
    CascadeMux I__5986 (
            .O(N__36953),
            .I(\PROM.ROMDATA.m506_cascade_ ));
    InMux I__5985 (
            .O(N__36950),
            .I(N__36944));
    InMux I__5984 (
            .O(N__36949),
            .I(N__36944));
    LocalMux I__5983 (
            .O(N__36944),
            .I(N__36941));
    Span4Mux_h I__5982 (
            .O(N__36941),
            .I(N__36938));
    Span4Mux_v I__5981 (
            .O(N__36938),
            .I(N__36935));
    Odrv4 I__5980 (
            .O(N__36935),
            .I(\PROM.ROMDATA.N_571_mux ));
    InMux I__5979 (
            .O(N__36932),
            .I(N__36929));
    LocalMux I__5978 (
            .O(N__36929),
            .I(N__36926));
    Span4Mux_v I__5977 (
            .O(N__36926),
            .I(N__36922));
    CascadeMux I__5976 (
            .O(N__36925),
            .I(N__36919));
    Span4Mux_h I__5975 (
            .O(N__36922),
            .I(N__36915));
    InMux I__5974 (
            .O(N__36919),
            .I(N__36910));
    InMux I__5973 (
            .O(N__36918),
            .I(N__36910));
    Span4Mux_v I__5972 (
            .O(N__36915),
            .I(N__36905));
    LocalMux I__5971 (
            .O(N__36910),
            .I(N__36905));
    Span4Mux_v I__5970 (
            .O(N__36905),
            .I(N__36902));
    Odrv4 I__5969 (
            .O(N__36902),
            .I(N_177));
    CascadeMux I__5968 (
            .O(N__36899),
            .I(\ALU.d_RNI64MA6Z0Z_0_cascade_ ));
    CascadeMux I__5967 (
            .O(N__36896),
            .I(\ALU.log_1_3_ns_1_1_0_cascade_ ));
    CascadeMux I__5966 (
            .O(N__36893),
            .I(\ALU.log_1_3_ns_1_0_cascade_ ));
    CascadeMux I__5965 (
            .O(N__36890),
            .I(\ALU.log_1_0_cascade_ ));
    CascadeMux I__5964 (
            .O(N__36887),
            .I(\ALU.status_8_5_0_cascade_ ));
    CascadeMux I__5963 (
            .O(N__36884),
            .I(N__36880));
    CascadeMux I__5962 (
            .O(N__36883),
            .I(N__36875));
    InMux I__5961 (
            .O(N__36880),
            .I(N__36872));
    InMux I__5960 (
            .O(N__36879),
            .I(N__36869));
    InMux I__5959 (
            .O(N__36878),
            .I(N__36866));
    InMux I__5958 (
            .O(N__36875),
            .I(N__36863));
    LocalMux I__5957 (
            .O(N__36872),
            .I(N__36860));
    LocalMux I__5956 (
            .O(N__36869),
            .I(N__36857));
    LocalMux I__5955 (
            .O(N__36866),
            .I(N__36854));
    LocalMux I__5954 (
            .O(N__36863),
            .I(N__36851));
    Span4Mux_h I__5953 (
            .O(N__36860),
            .I(N__36848));
    Span4Mux_h I__5952 (
            .O(N__36857),
            .I(N__36841));
    Span4Mux_h I__5951 (
            .O(N__36854),
            .I(N__36841));
    Span4Mux_h I__5950 (
            .O(N__36851),
            .I(N__36841));
    Odrv4 I__5949 (
            .O(N__36848),
            .I(\CONTROL.N_384_0 ));
    Odrv4 I__5948 (
            .O(N__36841),
            .I(\CONTROL.N_384_0 ));
    CascadeMux I__5947 (
            .O(N__36836),
            .I(\CONTROL.N_209_cascade_ ));
    CascadeMux I__5946 (
            .O(N__36833),
            .I(N__36830));
    InMux I__5945 (
            .O(N__36830),
            .I(N__36827));
    LocalMux I__5944 (
            .O(N__36827),
            .I(\CONTROL.un1_busState114_1_0_0_0 ));
    CascadeMux I__5943 (
            .O(N__36824),
            .I(\CONTROL.N_349_cascade_ ));
    InMux I__5942 (
            .O(N__36821),
            .I(N__36818));
    LocalMux I__5941 (
            .O(N__36818),
            .I(N__36814));
    InMux I__5940 (
            .O(N__36817),
            .I(N__36810));
    Span4Mux_h I__5939 (
            .O(N__36814),
            .I(N__36807));
    InMux I__5938 (
            .O(N__36813),
            .I(N__36804));
    LocalMux I__5937 (
            .O(N__36810),
            .I(\CONTROL.N_246 ));
    Odrv4 I__5936 (
            .O(N__36807),
            .I(\CONTROL.N_246 ));
    LocalMux I__5935 (
            .O(N__36804),
            .I(\CONTROL.N_246 ));
    InMux I__5934 (
            .O(N__36797),
            .I(N__36794));
    LocalMux I__5933 (
            .O(N__36794),
            .I(N__36791));
    Odrv4 I__5932 (
            .O(N__36791),
            .I(\CONTROL.m38_i_1 ));
    InMux I__5931 (
            .O(N__36788),
            .I(N__36785));
    LocalMux I__5930 (
            .O(N__36785),
            .I(\CONTROL.N_348 ));
    InMux I__5929 (
            .O(N__36782),
            .I(N__36779));
    LocalMux I__5928 (
            .O(N__36779),
            .I(N__36775));
    InMux I__5927 (
            .O(N__36778),
            .I(N__36772));
    Span4Mux_h I__5926 (
            .O(N__36775),
            .I(N__36769));
    LocalMux I__5925 (
            .O(N__36772),
            .I(N__36766));
    Span4Mux_h I__5924 (
            .O(N__36769),
            .I(N__36763));
    Span4Mux_h I__5923 (
            .O(N__36766),
            .I(N__36760));
    Odrv4 I__5922 (
            .O(N__36763),
            .I(\CONTROL.programCounter_1_12 ));
    Odrv4 I__5921 (
            .O(N__36760),
            .I(\CONTROL.programCounter_1_12 ));
    InMux I__5920 (
            .O(N__36755),
            .I(N__36752));
    LocalMux I__5919 (
            .O(N__36752),
            .I(\CONTROL.programCounter_1_reto_12 ));
    CascadeMux I__5918 (
            .O(N__36749),
            .I(controlWord_1_cascade_));
    CascadeMux I__5917 (
            .O(N__36746),
            .I(\CONTROL.N_420_cascade_ ));
    InMux I__5916 (
            .O(N__36743),
            .I(N__36740));
    LocalMux I__5915 (
            .O(N__36740),
            .I(N__36737));
    Span4Mux_v I__5914 (
            .O(N__36737),
            .I(N__36734));
    Sp12to4 I__5913 (
            .O(N__36734),
            .I(N__36731));
    Odrv12 I__5912 (
            .O(N__36731),
            .I(\CONTROL.programCounter_1_axb_5 ));
    InMux I__5911 (
            .O(N__36728),
            .I(N__36725));
    LocalMux I__5910 (
            .O(N__36725),
            .I(N__36722));
    Span4Mux_v I__5909 (
            .O(N__36722),
            .I(N__36719));
    Sp12to4 I__5908 (
            .O(N__36719),
            .I(N__36716));
    Odrv12 I__5907 (
            .O(N__36716),
            .I(\CONTROL.programCounter_1_axb_0 ));
    InMux I__5906 (
            .O(N__36713),
            .I(N__36710));
    LocalMux I__5905 (
            .O(N__36710),
            .I(N__36707));
    Span12Mux_h I__5904 (
            .O(N__36707),
            .I(N__36704));
    Odrv12 I__5903 (
            .O(N__36704),
            .I(\CONTROL.N_105_i ));
    InMux I__5902 (
            .O(N__36701),
            .I(N__36698));
    LocalMux I__5901 (
            .O(N__36698),
            .I(N__36695));
    Odrv12 I__5900 (
            .O(N__36695),
            .I(\CONTROL.N_427 ));
    CascadeMux I__5899 (
            .O(N__36692),
            .I(PROM_ROMDATA_dintern_5ro_cascade_));
    InMux I__5898 (
            .O(N__36689),
            .I(N__36685));
    InMux I__5897 (
            .O(N__36688),
            .I(N__36681));
    LocalMux I__5896 (
            .O(N__36685),
            .I(N__36677));
    InMux I__5895 (
            .O(N__36684),
            .I(N__36674));
    LocalMux I__5894 (
            .O(N__36681),
            .I(N__36671));
    InMux I__5893 (
            .O(N__36680),
            .I(N__36668));
    Span4Mux_h I__5892 (
            .O(N__36677),
            .I(N__36663));
    LocalMux I__5891 (
            .O(N__36674),
            .I(N__36663));
    Span4Mux_v I__5890 (
            .O(N__36671),
            .I(N__36658));
    LocalMux I__5889 (
            .O(N__36668),
            .I(N__36658));
    Span4Mux_h I__5888 (
            .O(N__36663),
            .I(N__36655));
    Odrv4 I__5887 (
            .O(N__36658),
            .I(\CONTROL.N_80_0 ));
    Odrv4 I__5886 (
            .O(N__36655),
            .I(\CONTROL.N_80_0 ));
    CascadeMux I__5885 (
            .O(N__36650),
            .I(N__36647));
    InMux I__5884 (
            .O(N__36647),
            .I(N__36644));
    LocalMux I__5883 (
            .O(N__36644),
            .I(N__36641));
    Span4Mux_h I__5882 (
            .O(N__36641),
            .I(N__36638));
    Odrv4 I__5881 (
            .O(N__36638),
            .I(\CONTROL.g0_1_i_3Z0Z_1 ));
    CascadeMux I__5880 (
            .O(N__36635),
            .I(\CONTROL.N_48_0_cascade_ ));
    InMux I__5879 (
            .O(N__36632),
            .I(N__36629));
    LocalMux I__5878 (
            .O(N__36629),
            .I(\CONTROL.un1_controlWord_14_i_0 ));
    CascadeMux I__5877 (
            .O(N__36626),
            .I(N__36622));
    CascadeMux I__5876 (
            .O(N__36625),
            .I(N__36618));
    InMux I__5875 (
            .O(N__36622),
            .I(N__36613));
    InMux I__5874 (
            .O(N__36621),
            .I(N__36613));
    InMux I__5873 (
            .O(N__36618),
            .I(N__36610));
    LocalMux I__5872 (
            .O(N__36613),
            .I(N__36606));
    LocalMux I__5871 (
            .O(N__36610),
            .I(N__36602));
    CascadeMux I__5870 (
            .O(N__36609),
            .I(N__36599));
    Span4Mux_v I__5869 (
            .O(N__36606),
            .I(N__36596));
    InMux I__5868 (
            .O(N__36605),
            .I(N__36593));
    Span4Mux_v I__5867 (
            .O(N__36602),
            .I(N__36590));
    InMux I__5866 (
            .O(N__36599),
            .I(N__36587));
    Odrv4 I__5865 (
            .O(N__36596),
            .I(\CONTROL.N_87_0 ));
    LocalMux I__5864 (
            .O(N__36593),
            .I(\CONTROL.N_87_0 ));
    Odrv4 I__5863 (
            .O(N__36590),
            .I(\CONTROL.N_87_0 ));
    LocalMux I__5862 (
            .O(N__36587),
            .I(\CONTROL.N_87_0 ));
    InMux I__5861 (
            .O(N__36578),
            .I(N__36575));
    LocalMux I__5860 (
            .O(N__36575),
            .I(N__36572));
    Span4Mux_h I__5859 (
            .O(N__36572),
            .I(N__36569));
    Odrv4 I__5858 (
            .O(N__36569),
            .I(\CONTROL.un1_busState97_1_0_1_0 ));
    InMux I__5857 (
            .O(N__36566),
            .I(N__36563));
    LocalMux I__5856 (
            .O(N__36563),
            .I(N__36560));
    Span4Mux_h I__5855 (
            .O(N__36560),
            .I(N__36557));
    Odrv4 I__5854 (
            .O(N__36557),
            .I(\CONTROL.dout_reto_7 ));
    InMux I__5853 (
            .O(N__36554),
            .I(N__36551));
    LocalMux I__5852 (
            .O(N__36551),
            .I(N__36548));
    Span4Mux_h I__5851 (
            .O(N__36548),
            .I(N__36545));
    Span4Mux_h I__5850 (
            .O(N__36545),
            .I(N__36542));
    Odrv4 I__5849 (
            .O(N__36542),
            .I(\CONTROL.addrstack_reto_7 ));
    CascadeMux I__5848 (
            .O(N__36539),
            .I(\CONTROL.N_422_cascade_ ));
    CascadeMux I__5847 (
            .O(N__36536),
            .I(progRomAddress_7_cascade_));
    CascadeMux I__5846 (
            .O(N__36533),
            .I(\CONTROL.N_340_cascade_ ));
    CEMux I__5845 (
            .O(N__36530),
            .I(N__36527));
    LocalMux I__5844 (
            .O(N__36527),
            .I(N__36524));
    Span4Mux_h I__5843 (
            .O(N__36524),
            .I(N__36521));
    Odrv4 I__5842 (
            .O(N__36521),
            .I(\CONTROL.un1_busState103_0_0 ));
    CascadeMux I__5841 (
            .O(N__36518),
            .I(\CONTROL.un1_busState114_2_0_0_xZ0Z0_cascade_ ));
    InMux I__5840 (
            .O(N__36515),
            .I(N__36512));
    LocalMux I__5839 (
            .O(N__36512),
            .I(\CONTROL.un1_busState114_2_0_0_xZ0Z1 ));
    CascadeMux I__5838 (
            .O(N__36509),
            .I(\CONTROL.un1_busState114_2_0_0_0_cascade_ ));
    InMux I__5837 (
            .O(N__36506),
            .I(N__36503));
    LocalMux I__5836 (
            .O(N__36503),
            .I(N__36500));
    Span4Mux_h I__5835 (
            .O(N__36500),
            .I(N__36497));
    Odrv4 I__5834 (
            .O(N__36497),
            .I(\CONTROL.aluReadBus_1_sqmuxa_0_a2_2Z0Z_0 ));
    InMux I__5833 (
            .O(N__36494),
            .I(N__36491));
    LocalMux I__5832 (
            .O(N__36491),
            .I(N__36488));
    Span4Mux_h I__5831 (
            .O(N__36488),
            .I(N__36484));
    CascadeMux I__5830 (
            .O(N__36487),
            .I(N__36481));
    Span4Mux_v I__5829 (
            .O(N__36484),
            .I(N__36478));
    InMux I__5828 (
            .O(N__36481),
            .I(N__36475));
    Odrv4 I__5827 (
            .O(N__36478),
            .I(\CONTROL.N_83_0 ));
    LocalMux I__5826 (
            .O(N__36475),
            .I(\CONTROL.N_83_0 ));
    InMux I__5825 (
            .O(N__36470),
            .I(N__36467));
    LocalMux I__5824 (
            .O(N__36467),
            .I(N__36464));
    Span4Mux_v I__5823 (
            .O(N__36464),
            .I(N__36461));
    Span4Mux_h I__5822 (
            .O(N__36461),
            .I(N__36458));
    Span4Mux_h I__5821 (
            .O(N__36458),
            .I(N__36455));
    Odrv4 I__5820 (
            .O(N__36455),
            .I(\CONTROL.increment28lto5_1_1_0 ));
    InMux I__5819 (
            .O(N__36452),
            .I(N__36449));
    LocalMux I__5818 (
            .O(N__36449),
            .I(N__36444));
    CascadeMux I__5817 (
            .O(N__36448),
            .I(N__36440));
    CascadeMux I__5816 (
            .O(N__36447),
            .I(N__36437));
    Span4Mux_v I__5815 (
            .O(N__36444),
            .I(N__36434));
    InMux I__5814 (
            .O(N__36443),
            .I(N__36426));
    InMux I__5813 (
            .O(N__36440),
            .I(N__36426));
    InMux I__5812 (
            .O(N__36437),
            .I(N__36426));
    Sp12to4 I__5811 (
            .O(N__36434),
            .I(N__36423));
    InMux I__5810 (
            .O(N__36433),
            .I(N__36420));
    LocalMux I__5809 (
            .O(N__36426),
            .I(N__36417));
    Odrv12 I__5808 (
            .O(N__36423),
            .I(\CONTROL.N_101_0 ));
    LocalMux I__5807 (
            .O(N__36420),
            .I(\CONTROL.N_101_0 ));
    Odrv4 I__5806 (
            .O(N__36417),
            .I(\CONTROL.N_101_0 ));
    CascadeMux I__5805 (
            .O(N__36410),
            .I(\CONTROL.N_320_cascade_ ));
    CascadeMux I__5804 (
            .O(N__36407),
            .I(\CONTROL.un1_busState103_0_0_cascade_ ));
    CascadeMux I__5803 (
            .O(N__36404),
            .I(N__36401));
    InMux I__5802 (
            .O(N__36401),
            .I(N__36398));
    LocalMux I__5801 (
            .O(N__36398),
            .I(N__36394));
    CascadeMux I__5800 (
            .O(N__36397),
            .I(N__36391));
    Span4Mux_h I__5799 (
            .O(N__36394),
            .I(N__36388));
    InMux I__5798 (
            .O(N__36391),
            .I(N__36385));
    Span4Mux_h I__5797 (
            .O(N__36388),
            .I(N__36382));
    LocalMux I__5796 (
            .O(N__36385),
            .I(\CONTROL.N_95_0 ));
    Odrv4 I__5795 (
            .O(N__36382),
            .I(\CONTROL.N_95_0 ));
    InMux I__5794 (
            .O(N__36377),
            .I(N__36374));
    LocalMux I__5793 (
            .O(N__36374),
            .I(\CONTROL.N_318 ));
    InMux I__5792 (
            .O(N__36371),
            .I(N__36365));
    InMux I__5791 (
            .O(N__36370),
            .I(N__36365));
    LocalMux I__5790 (
            .O(N__36365),
            .I(N__36358));
    InMux I__5789 (
            .O(N__36364),
            .I(N__36353));
    InMux I__5788 (
            .O(N__36363),
            .I(N__36353));
    InMux I__5787 (
            .O(N__36362),
            .I(N__36348));
    InMux I__5786 (
            .O(N__36361),
            .I(N__36348));
    Odrv4 I__5785 (
            .O(N__36358),
            .I(aluOperand1_fast_2));
    LocalMux I__5784 (
            .O(N__36353),
            .I(aluOperand1_fast_2));
    LocalMux I__5783 (
            .O(N__36348),
            .I(aluOperand1_fast_2));
    InMux I__5782 (
            .O(N__36341),
            .I(N__36333));
    InMux I__5781 (
            .O(N__36340),
            .I(N__36333));
    InMux I__5780 (
            .O(N__36339),
            .I(N__36328));
    InMux I__5779 (
            .O(N__36338),
            .I(N__36328));
    LocalMux I__5778 (
            .O(N__36333),
            .I(N__36319));
    LocalMux I__5777 (
            .O(N__36328),
            .I(N__36319));
    InMux I__5776 (
            .O(N__36327),
            .I(N__36310));
    InMux I__5775 (
            .O(N__36326),
            .I(N__36310));
    InMux I__5774 (
            .O(N__36325),
            .I(N__36305));
    InMux I__5773 (
            .O(N__36324),
            .I(N__36305));
    Span4Mux_h I__5772 (
            .O(N__36319),
            .I(N__36302));
    InMux I__5771 (
            .O(N__36318),
            .I(N__36297));
    InMux I__5770 (
            .O(N__36317),
            .I(N__36297));
    InMux I__5769 (
            .O(N__36316),
            .I(N__36292));
    InMux I__5768 (
            .O(N__36315),
            .I(N__36292));
    LocalMux I__5767 (
            .O(N__36310),
            .I(aluOperand1_fast_1));
    LocalMux I__5766 (
            .O(N__36305),
            .I(aluOperand1_fast_1));
    Odrv4 I__5765 (
            .O(N__36302),
            .I(aluOperand1_fast_1));
    LocalMux I__5764 (
            .O(N__36297),
            .I(aluOperand1_fast_1));
    LocalMux I__5763 (
            .O(N__36292),
            .I(aluOperand1_fast_1));
    InMux I__5762 (
            .O(N__36281),
            .I(N__36278));
    LocalMux I__5761 (
            .O(N__36278),
            .I(N__36275));
    Span4Mux_h I__5760 (
            .O(N__36275),
            .I(N__36272));
    Span4Mux_v I__5759 (
            .O(N__36272),
            .I(N__36269));
    Odrv4 I__5758 (
            .O(N__36269),
            .I(\CONTROL.increment28lto5_1_1_3 ));
    CascadeMux I__5757 (
            .O(N__36266),
            .I(\CONTROL.increment28lto5_1_1_1_cascade_ ));
    CascadeMux I__5756 (
            .O(N__36263),
            .I(N__36260));
    InMux I__5755 (
            .O(N__36260),
            .I(N__36257));
    LocalMux I__5754 (
            .O(N__36257),
            .I(N__36254));
    Odrv4 I__5753 (
            .O(N__36254),
            .I(\CONTROL.g0_3_i_a7Z0Z_3 ));
    CascadeMux I__5752 (
            .O(N__36251),
            .I(\PROM.ROMDATA.m221cf1_cascade_ ));
    InMux I__5751 (
            .O(N__36248),
            .I(N__36245));
    LocalMux I__5750 (
            .O(N__36245),
            .I(\PROM.ROMDATA.m221cf1 ));
    CEMux I__5749 (
            .O(N__36242),
            .I(N__36237));
    CEMux I__5748 (
            .O(N__36241),
            .I(N__36234));
    CEMux I__5747 (
            .O(N__36240),
            .I(N__36231));
    LocalMux I__5746 (
            .O(N__36237),
            .I(N__36228));
    LocalMux I__5745 (
            .O(N__36234),
            .I(N__36225));
    LocalMux I__5744 (
            .O(N__36231),
            .I(N__36222));
    Span4Mux_v I__5743 (
            .O(N__36228),
            .I(N__36219));
    Span4Mux_v I__5742 (
            .O(N__36225),
            .I(N__36216));
    Span4Mux_h I__5741 (
            .O(N__36222),
            .I(N__36213));
    Odrv4 I__5740 (
            .O(N__36219),
            .I(\CONTROL.un1_busState98_1_0_0_0 ));
    Odrv4 I__5739 (
            .O(N__36216),
            .I(\CONTROL.un1_busState98_1_0_0_0 ));
    Odrv4 I__5738 (
            .O(N__36213),
            .I(\CONTROL.un1_busState98_1_0_0_0 ));
    InMux I__5737 (
            .O(N__36206),
            .I(N__36200));
    InMux I__5736 (
            .O(N__36205),
            .I(N__36200));
    LocalMux I__5735 (
            .O(N__36200),
            .I(\PROM.ROMDATA.m217 ));
    InMux I__5734 (
            .O(N__36197),
            .I(N__36191));
    InMux I__5733 (
            .O(N__36196),
            .I(N__36191));
    LocalMux I__5732 (
            .O(N__36191),
            .I(\PROM.ROMDATA.m221cf0 ));
    InMux I__5731 (
            .O(N__36188),
            .I(N__36185));
    LocalMux I__5730 (
            .O(N__36185),
            .I(N__36181));
    InMux I__5729 (
            .O(N__36184),
            .I(N__36178));
    Span4Mux_h I__5728 (
            .O(N__36181),
            .I(N__36175));
    LocalMux I__5727 (
            .O(N__36178),
            .I(\ALU.dZ0Z_11 ));
    Odrv4 I__5726 (
            .O(N__36175),
            .I(\ALU.dZ0Z_11 ));
    InMux I__5725 (
            .O(N__36170),
            .I(N__36167));
    LocalMux I__5724 (
            .O(N__36167),
            .I(N__36164));
    Span4Mux_v I__5723 (
            .O(N__36164),
            .I(N__36161));
    Odrv4 I__5722 (
            .O(N__36161),
            .I(\ALU.d_RNI6DCTZ0Z_11 ));
    InMux I__5721 (
            .O(N__36158),
            .I(N__36155));
    LocalMux I__5720 (
            .O(N__36155),
            .I(N__36152));
    Span4Mux_v I__5719 (
            .O(N__36152),
            .I(N__36149));
    Odrv4 I__5718 (
            .O(N__36149),
            .I(\ALU.N_920 ));
    InMux I__5717 (
            .O(N__36146),
            .I(N__36143));
    LocalMux I__5716 (
            .O(N__36143),
            .I(\ALU.operand2_3_ns_1_15 ));
    CascadeMux I__5715 (
            .O(N__36140),
            .I(\ALU.dout_3_ns_1_15_cascade_ ));
    InMux I__5714 (
            .O(N__36137),
            .I(N__36133));
    InMux I__5713 (
            .O(N__36136),
            .I(N__36130));
    LocalMux I__5712 (
            .O(N__36133),
            .I(N__36127));
    LocalMux I__5711 (
            .O(N__36130),
            .I(N__36124));
    Span4Mux_v I__5710 (
            .O(N__36127),
            .I(N__36121));
    Span4Mux_v I__5709 (
            .O(N__36124),
            .I(N__36118));
    Span4Mux_h I__5708 (
            .O(N__36121),
            .I(N__36115));
    Sp12to4 I__5707 (
            .O(N__36118),
            .I(N__36110));
    Sp12to4 I__5706 (
            .O(N__36115),
            .I(N__36110));
    Span12Mux_h I__5705 (
            .O(N__36110),
            .I(N__36107));
    Odrv12 I__5704 (
            .O(N__36107),
            .I(\ALU.cZ0Z_10 ));
    InMux I__5703 (
            .O(N__36104),
            .I(N__36100));
    InMux I__5702 (
            .O(N__36103),
            .I(N__36097));
    LocalMux I__5701 (
            .O(N__36100),
            .I(N__36092));
    LocalMux I__5700 (
            .O(N__36097),
            .I(N__36092));
    Span4Mux_v I__5699 (
            .O(N__36092),
            .I(N__36089));
    Span4Mux_h I__5698 (
            .O(N__36089),
            .I(N__36086));
    Odrv4 I__5697 (
            .O(N__36086),
            .I(\ALU.cZ0Z_11 ));
    InMux I__5696 (
            .O(N__36083),
            .I(N__36080));
    LocalMux I__5695 (
            .O(N__36080),
            .I(N__36077));
    Span4Mux_h I__5694 (
            .O(N__36077),
            .I(N__36074));
    Span4Mux_v I__5693 (
            .O(N__36074),
            .I(N__36070));
    InMux I__5692 (
            .O(N__36073),
            .I(N__36067));
    Odrv4 I__5691 (
            .O(N__36070),
            .I(\ALU.dZ0Z_2 ));
    LocalMux I__5690 (
            .O(N__36067),
            .I(\ALU.dZ0Z_2 ));
    InMux I__5689 (
            .O(N__36062),
            .I(N__36059));
    LocalMux I__5688 (
            .O(N__36059),
            .I(N__36056));
    Span4Mux_v I__5687 (
            .O(N__36056),
            .I(N__36052));
    InMux I__5686 (
            .O(N__36055),
            .I(N__36049));
    Span4Mux_h I__5685 (
            .O(N__36052),
            .I(N__36046));
    LocalMux I__5684 (
            .O(N__36049),
            .I(N__36043));
    Span4Mux_v I__5683 (
            .O(N__36046),
            .I(N__36040));
    Odrv12 I__5682 (
            .O(N__36043),
            .I(\ALU.dZ0Z_6 ));
    Odrv4 I__5681 (
            .O(N__36040),
            .I(\ALU.dZ0Z_6 ));
    InMux I__5680 (
            .O(N__36035),
            .I(N__36031));
    CascadeMux I__5679 (
            .O(N__36034),
            .I(N__36028));
    LocalMux I__5678 (
            .O(N__36031),
            .I(N__36025));
    InMux I__5677 (
            .O(N__36028),
            .I(N__36022));
    Span4Mux_h I__5676 (
            .O(N__36025),
            .I(N__36019));
    LocalMux I__5675 (
            .O(N__36022),
            .I(N__36016));
    Span4Mux_h I__5674 (
            .O(N__36019),
            .I(N__36013));
    Odrv12 I__5673 (
            .O(N__36016),
            .I(\ALU.dZ0Z_10 ));
    Odrv4 I__5672 (
            .O(N__36013),
            .I(\ALU.dZ0Z_10 ));
    CascadeMux I__5671 (
            .O(N__36008),
            .I(N__36005));
    InMux I__5670 (
            .O(N__36005),
            .I(N__36000));
    CascadeMux I__5669 (
            .O(N__36004),
            .I(N__35997));
    InMux I__5668 (
            .O(N__36003),
            .I(N__35994));
    LocalMux I__5667 (
            .O(N__36000),
            .I(N__35991));
    InMux I__5666 (
            .O(N__35997),
            .I(N__35988));
    LocalMux I__5665 (
            .O(N__35994),
            .I(N__35985));
    Span4Mux_v I__5664 (
            .O(N__35991),
            .I(N__35980));
    LocalMux I__5663 (
            .O(N__35988),
            .I(N__35980));
    Span4Mux_h I__5662 (
            .O(N__35985),
            .I(N__35975));
    Span4Mux_v I__5661 (
            .O(N__35980),
            .I(N__35975));
    Span4Mux_h I__5660 (
            .O(N__35975),
            .I(N__35972));
    Odrv4 I__5659 (
            .O(N__35972),
            .I(f_10));
    CascadeMux I__5658 (
            .O(N__35969),
            .I(N__35964));
    CascadeMux I__5657 (
            .O(N__35968),
            .I(N__35961));
    InMux I__5656 (
            .O(N__35967),
            .I(N__35958));
    InMux I__5655 (
            .O(N__35964),
            .I(N__35953));
    InMux I__5654 (
            .O(N__35961),
            .I(N__35953));
    LocalMux I__5653 (
            .O(N__35958),
            .I(N__35950));
    LocalMux I__5652 (
            .O(N__35953),
            .I(N__35947));
    Sp12to4 I__5651 (
            .O(N__35950),
            .I(N__35944));
    Span4Mux_h I__5650 (
            .O(N__35947),
            .I(N__35941));
    Span12Mux_v I__5649 (
            .O(N__35944),
            .I(N__35938));
    Span4Mux_h I__5648 (
            .O(N__35941),
            .I(N__35935));
    Odrv12 I__5647 (
            .O(N__35938),
            .I(f_11));
    Odrv4 I__5646 (
            .O(N__35935),
            .I(f_11));
    CEMux I__5645 (
            .O(N__35930),
            .I(N__35924));
    CEMux I__5644 (
            .O(N__35929),
            .I(N__35921));
    CEMux I__5643 (
            .O(N__35928),
            .I(N__35918));
    CEMux I__5642 (
            .O(N__35927),
            .I(N__35915));
    LocalMux I__5641 (
            .O(N__35924),
            .I(N__35912));
    LocalMux I__5640 (
            .O(N__35921),
            .I(N__35909));
    LocalMux I__5639 (
            .O(N__35918),
            .I(N__35904));
    LocalMux I__5638 (
            .O(N__35915),
            .I(N__35904));
    Span4Mux_v I__5637 (
            .O(N__35912),
            .I(N__35901));
    Span4Mux_v I__5636 (
            .O(N__35909),
            .I(N__35898));
    Span4Mux_v I__5635 (
            .O(N__35904),
            .I(N__35895));
    Span4Mux_v I__5634 (
            .O(N__35901),
            .I(N__35888));
    Span4Mux_v I__5633 (
            .O(N__35898),
            .I(N__35888));
    Span4Mux_h I__5632 (
            .O(N__35895),
            .I(N__35888));
    Span4Mux_h I__5631 (
            .O(N__35888),
            .I(N__35885));
    Sp12to4 I__5630 (
            .O(N__35885),
            .I(N__35882));
    Span12Mux_v I__5629 (
            .O(N__35882),
            .I(N__35879));
    Odrv12 I__5628 (
            .O(N__35879),
            .I(CONSTANT_ZERO_NET));
    InMux I__5627 (
            .O(N__35876),
            .I(N__35873));
    LocalMux I__5626 (
            .O(N__35873),
            .I(N__35869));
    InMux I__5625 (
            .O(N__35872),
            .I(N__35866));
    Span4Mux_v I__5624 (
            .O(N__35869),
            .I(N__35863));
    LocalMux I__5623 (
            .O(N__35866),
            .I(N__35858));
    Span4Mux_h I__5622 (
            .O(N__35863),
            .I(N__35858));
    Span4Mux_v I__5621 (
            .O(N__35858),
            .I(N__35855));
    Odrv4 I__5620 (
            .O(N__35855),
            .I(\ALU.cZ0Z_2 ));
    InMux I__5619 (
            .O(N__35852),
            .I(N__35848));
    InMux I__5618 (
            .O(N__35851),
            .I(N__35845));
    LocalMux I__5617 (
            .O(N__35848),
            .I(N__35842));
    LocalMux I__5616 (
            .O(N__35845),
            .I(N__35837));
    Span12Mux_v I__5615 (
            .O(N__35842),
            .I(N__35837));
    Odrv12 I__5614 (
            .O(N__35837),
            .I(\ALU.cZ0Z_4 ));
    InMux I__5613 (
            .O(N__35834),
            .I(N__35830));
    InMux I__5612 (
            .O(N__35833),
            .I(N__35827));
    LocalMux I__5611 (
            .O(N__35830),
            .I(N__35824));
    LocalMux I__5610 (
            .O(N__35827),
            .I(N__35821));
    Span4Mux_v I__5609 (
            .O(N__35824),
            .I(N__35818));
    Span4Mux_h I__5608 (
            .O(N__35821),
            .I(N__35815));
    Span4Mux_h I__5607 (
            .O(N__35818),
            .I(N__35812));
    Odrv4 I__5606 (
            .O(N__35815),
            .I(\ALU.cZ0Z_6 ));
    Odrv4 I__5605 (
            .O(N__35812),
            .I(\ALU.cZ0Z_6 ));
    CascadeMux I__5604 (
            .O(N__35807),
            .I(N__35804));
    InMux I__5603 (
            .O(N__35804),
            .I(N__35801));
    LocalMux I__5602 (
            .O(N__35801),
            .I(N__35798));
    Span4Mux_h I__5601 (
            .O(N__35798),
            .I(N__35793));
    InMux I__5600 (
            .O(N__35797),
            .I(N__35790));
    InMux I__5599 (
            .O(N__35796),
            .I(N__35787));
    Span4Mux_h I__5598 (
            .O(N__35793),
            .I(N__35784));
    LocalMux I__5597 (
            .O(N__35790),
            .I(N__35779));
    LocalMux I__5596 (
            .O(N__35787),
            .I(N__35779));
    Sp12to4 I__5595 (
            .O(N__35784),
            .I(N__35776));
    Span12Mux_v I__5594 (
            .O(N__35779),
            .I(N__35773));
    Odrv12 I__5593 (
            .O(N__35776),
            .I(g_4));
    Odrv12 I__5592 (
            .O(N__35773),
            .I(g_4));
    InMux I__5591 (
            .O(N__35768),
            .I(N__35765));
    LocalMux I__5590 (
            .O(N__35765),
            .I(N__35761));
    InMux I__5589 (
            .O(N__35764),
            .I(N__35757));
    Span4Mux_h I__5588 (
            .O(N__35761),
            .I(N__35754));
    InMux I__5587 (
            .O(N__35760),
            .I(N__35751));
    LocalMux I__5586 (
            .O(N__35757),
            .I(N__35748));
    Span4Mux_v I__5585 (
            .O(N__35754),
            .I(N__35745));
    LocalMux I__5584 (
            .O(N__35751),
            .I(N__35742));
    Span4Mux_v I__5583 (
            .O(N__35748),
            .I(N__35739));
    Span4Mux_h I__5582 (
            .O(N__35745),
            .I(N__35736));
    Span12Mux_v I__5581 (
            .O(N__35742),
            .I(N__35731));
    Sp12to4 I__5580 (
            .O(N__35739),
            .I(N__35731));
    Span4Mux_h I__5579 (
            .O(N__35736),
            .I(N__35728));
    Odrv12 I__5578 (
            .O(N__35731),
            .I(g_6));
    Odrv4 I__5577 (
            .O(N__35728),
            .I(g_6));
    CascadeMux I__5576 (
            .O(N__35723),
            .I(N__35719));
    InMux I__5575 (
            .O(N__35722),
            .I(N__35716));
    InMux I__5574 (
            .O(N__35719),
            .I(N__35713));
    LocalMux I__5573 (
            .O(N__35716),
            .I(N__35709));
    LocalMux I__5572 (
            .O(N__35713),
            .I(N__35706));
    InMux I__5571 (
            .O(N__35712),
            .I(N__35703));
    Span4Mux_h I__5570 (
            .O(N__35709),
            .I(N__35700));
    Span4Mux_v I__5569 (
            .O(N__35706),
            .I(N__35695));
    LocalMux I__5568 (
            .O(N__35703),
            .I(N__35695));
    Span4Mux_v I__5567 (
            .O(N__35700),
            .I(N__35692));
    Sp12to4 I__5566 (
            .O(N__35695),
            .I(N__35689));
    Sp12to4 I__5565 (
            .O(N__35692),
            .I(N__35686));
    Span12Mux_h I__5564 (
            .O(N__35689),
            .I(N__35683));
    Odrv12 I__5563 (
            .O(N__35686),
            .I(g_10));
    Odrv12 I__5562 (
            .O(N__35683),
            .I(g_10));
    InMux I__5561 (
            .O(N__35678),
            .I(N__35675));
    LocalMux I__5560 (
            .O(N__35675),
            .I(N__35672));
    Span4Mux_v I__5559 (
            .O(N__35672),
            .I(N__35668));
    CascadeMux I__5558 (
            .O(N__35671),
            .I(N__35665));
    Span4Mux_h I__5557 (
            .O(N__35668),
            .I(N__35661));
    InMux I__5556 (
            .O(N__35665),
            .I(N__35658));
    InMux I__5555 (
            .O(N__35664),
            .I(N__35655));
    Span4Mux_v I__5554 (
            .O(N__35661),
            .I(N__35652));
    LocalMux I__5553 (
            .O(N__35658),
            .I(N__35647));
    LocalMux I__5552 (
            .O(N__35655),
            .I(N__35647));
    Span4Mux_v I__5551 (
            .O(N__35652),
            .I(N__35644));
    Span4Mux_v I__5550 (
            .O(N__35647),
            .I(N__35641));
    Odrv4 I__5549 (
            .O(N__35644),
            .I(g_11));
    Odrv4 I__5548 (
            .O(N__35641),
            .I(g_11));
    InMux I__5547 (
            .O(N__35636),
            .I(N__35633));
    LocalMux I__5546 (
            .O(N__35633),
            .I(N__35628));
    InMux I__5545 (
            .O(N__35632),
            .I(N__35625));
    CascadeMux I__5544 (
            .O(N__35631),
            .I(N__35622));
    Span4Mux_v I__5543 (
            .O(N__35628),
            .I(N__35619));
    LocalMux I__5542 (
            .O(N__35625),
            .I(N__35616));
    InMux I__5541 (
            .O(N__35622),
            .I(N__35613));
    Span4Mux_h I__5540 (
            .O(N__35619),
            .I(N__35610));
    Span4Mux_h I__5539 (
            .O(N__35616),
            .I(N__35605));
    LocalMux I__5538 (
            .O(N__35613),
            .I(N__35605));
    Span4Mux_v I__5537 (
            .O(N__35610),
            .I(N__35602));
    Span4Mux_v I__5536 (
            .O(N__35605),
            .I(N__35599));
    Odrv4 I__5535 (
            .O(N__35602),
            .I(f_2));
    Odrv4 I__5534 (
            .O(N__35599),
            .I(f_2));
    InMux I__5533 (
            .O(N__35594),
            .I(N__35591));
    LocalMux I__5532 (
            .O(N__35591),
            .I(\ALU.d_RNIUT8OG4Z0Z_0 ));
    CascadeMux I__5531 (
            .O(N__35588),
            .I(N__35585));
    InMux I__5530 (
            .O(N__35585),
            .I(N__35582));
    LocalMux I__5529 (
            .O(N__35582),
            .I(N__35579));
    Odrv4 I__5528 (
            .O(N__35579),
            .I(\ALU.lshift_3_ns_1_14 ));
    CascadeMux I__5527 (
            .O(N__35576),
            .I(\ALU.N_646_cascade_ ));
    CascadeMux I__5526 (
            .O(N__35573),
            .I(\ALU.lshift_15_ns_1_14_cascade_ ));
    CascadeMux I__5525 (
            .O(N__35570),
            .I(N__35567));
    InMux I__5524 (
            .O(N__35567),
            .I(N__35563));
    InMux I__5523 (
            .O(N__35566),
            .I(N__35560));
    LocalMux I__5522 (
            .O(N__35563),
            .I(N__35557));
    LocalMux I__5521 (
            .O(N__35560),
            .I(N__35554));
    Span4Mux_h I__5520 (
            .O(N__35557),
            .I(N__35551));
    Span4Mux_v I__5519 (
            .O(N__35554),
            .I(N__35547));
    Span4Mux_h I__5518 (
            .O(N__35551),
            .I(N__35544));
    InMux I__5517 (
            .O(N__35550),
            .I(N__35541));
    Span4Mux_v I__5516 (
            .O(N__35547),
            .I(N__35538));
    Span4Mux_v I__5515 (
            .O(N__35544),
            .I(N__35533));
    LocalMux I__5514 (
            .O(N__35541),
            .I(N__35533));
    Sp12to4 I__5513 (
            .O(N__35538),
            .I(N__35530));
    Span4Mux_v I__5512 (
            .O(N__35533),
            .I(N__35527));
    Span12Mux_h I__5511 (
            .O(N__35530),
            .I(N__35524));
    Span4Mux_h I__5510 (
            .O(N__35527),
            .I(N__35521));
    Odrv12 I__5509 (
            .O(N__35524),
            .I(g_2));
    Odrv4 I__5508 (
            .O(N__35521),
            .I(g_2));
    InMux I__5507 (
            .O(N__35516),
            .I(N__35513));
    LocalMux I__5506 (
            .O(N__35513),
            .I(N__35510));
    Span4Mux_h I__5505 (
            .O(N__35510),
            .I(N__35507));
    Odrv4 I__5504 (
            .O(N__35507),
            .I(\ALU.mult_17_8 ));
    CascadeMux I__5503 (
            .O(N__35504),
            .I(N__35501));
    InMux I__5502 (
            .O(N__35501),
            .I(N__35498));
    LocalMux I__5501 (
            .O(N__35498),
            .I(\ALU.mult_19_8 ));
    InMux I__5500 (
            .O(N__35495),
            .I(\ALU.mult_25_c7 ));
    InMux I__5499 (
            .O(N__35492),
            .I(N__35489));
    LocalMux I__5498 (
            .O(N__35489),
            .I(N__35486));
    Span4Mux_h I__5497 (
            .O(N__35486),
            .I(N__35483));
    Odrv4 I__5496 (
            .O(N__35483),
            .I(\ALU.mult_17_9 ));
    CascadeMux I__5495 (
            .O(N__35480),
            .I(N__35477));
    InMux I__5494 (
            .O(N__35477),
            .I(N__35474));
    LocalMux I__5493 (
            .O(N__35474),
            .I(\ALU.mult_19_9 ));
    InMux I__5492 (
            .O(N__35471),
            .I(\ALU.mult_25_c8 ));
    InMux I__5491 (
            .O(N__35468),
            .I(N__35465));
    LocalMux I__5490 (
            .O(N__35465),
            .I(\ALU.mult_19_10 ));
    CascadeMux I__5489 (
            .O(N__35462),
            .I(N__35459));
    InMux I__5488 (
            .O(N__35459),
            .I(N__35456));
    LocalMux I__5487 (
            .O(N__35456),
            .I(N__35453));
    Span4Mux_h I__5486 (
            .O(N__35453),
            .I(N__35450));
    Odrv4 I__5485 (
            .O(N__35450),
            .I(\ALU.mult_17_10 ));
    InMux I__5484 (
            .O(N__35447),
            .I(\ALU.mult_25_c9 ));
    InMux I__5483 (
            .O(N__35444),
            .I(N__35441));
    LocalMux I__5482 (
            .O(N__35441),
            .I(N__35438));
    Span4Mux_h I__5481 (
            .O(N__35438),
            .I(N__35435));
    Odrv4 I__5480 (
            .O(N__35435),
            .I(\ALU.mult_17_11 ));
    CascadeMux I__5479 (
            .O(N__35432),
            .I(N__35429));
    InMux I__5478 (
            .O(N__35429),
            .I(N__35426));
    LocalMux I__5477 (
            .O(N__35426),
            .I(\ALU.mult_19_11 ));
    InMux I__5476 (
            .O(N__35423),
            .I(\ALU.mult_25_c10 ));
    InMux I__5475 (
            .O(N__35420),
            .I(N__35417));
    LocalMux I__5474 (
            .O(N__35417),
            .I(N__35414));
    Span4Mux_h I__5473 (
            .O(N__35414),
            .I(N__35411));
    Odrv4 I__5472 (
            .O(N__35411),
            .I(\ALU.mult_17_12 ));
    CascadeMux I__5471 (
            .O(N__35408),
            .I(N__35405));
    InMux I__5470 (
            .O(N__35405),
            .I(N__35402));
    LocalMux I__5469 (
            .O(N__35402),
            .I(\ALU.mult_19_12 ));
    InMux I__5468 (
            .O(N__35399),
            .I(bfn_16_10_0_));
    InMux I__5467 (
            .O(N__35396),
            .I(N__35393));
    LocalMux I__5466 (
            .O(N__35393),
            .I(N__35390));
    Span4Mux_h I__5465 (
            .O(N__35390),
            .I(N__35387));
    Odrv4 I__5464 (
            .O(N__35387),
            .I(\ALU.mult_17_13 ));
    CascadeMux I__5463 (
            .O(N__35384),
            .I(N__35381));
    InMux I__5462 (
            .O(N__35381),
            .I(N__35378));
    LocalMux I__5461 (
            .O(N__35378),
            .I(\ALU.mult_19_13 ));
    InMux I__5460 (
            .O(N__35375),
            .I(\ALU.mult_25_c12 ));
    InMux I__5459 (
            .O(N__35372),
            .I(N__35369));
    LocalMux I__5458 (
            .O(N__35369),
            .I(N__35366));
    Span4Mux_h I__5457 (
            .O(N__35366),
            .I(N__35363));
    Odrv4 I__5456 (
            .O(N__35363),
            .I(\ALU.mult_17_14 ));
    CascadeMux I__5455 (
            .O(N__35360),
            .I(N__35357));
    InMux I__5454 (
            .O(N__35357),
            .I(N__35354));
    LocalMux I__5453 (
            .O(N__35354),
            .I(\ALU.mult_19_14 ));
    InMux I__5452 (
            .O(N__35351),
            .I(\ALU.mult_25_c13 ));
    InMux I__5451 (
            .O(N__35348),
            .I(N__35345));
    LocalMux I__5450 (
            .O(N__35345),
            .I(N__35342));
    Span4Mux_h I__5449 (
            .O(N__35342),
            .I(N__35339));
    Odrv4 I__5448 (
            .O(N__35339),
            .I(\ALU.mult_424_c_RNIUVTALZ0Z4 ));
    InMux I__5447 (
            .O(N__35336),
            .I(\ALU.mult_25_c14 ));
    CascadeMux I__5446 (
            .O(N__35333),
            .I(\PROM.ROMDATA.m2_cascade_ ));
    InMux I__5445 (
            .O(N__35330),
            .I(N__35327));
    LocalMux I__5444 (
            .O(N__35327),
            .I(\ALU.mult_7_6 ));
    CascadeMux I__5443 (
            .O(N__35324),
            .I(N__35321));
    InMux I__5442 (
            .O(N__35321),
            .I(N__35318));
    LocalMux I__5441 (
            .O(N__35318),
            .I(N__35315));
    Span4Mux_h I__5440 (
            .O(N__35315),
            .I(N__35312));
    Span4Mux_h I__5439 (
            .O(N__35312),
            .I(N__35309));
    Odrv4 I__5438 (
            .O(N__35309),
            .I(\ALU.status_18_cry_0_c_RNOZ0 ));
    InMux I__5437 (
            .O(N__35306),
            .I(N__35303));
    LocalMux I__5436 (
            .O(N__35303),
            .I(N__35300));
    Odrv4 I__5435 (
            .O(N__35300),
            .I(\ALU.mult_5_4 ));
    CascadeMux I__5434 (
            .O(N__35297),
            .I(N__35294));
    InMux I__5433 (
            .O(N__35294),
            .I(N__35291));
    LocalMux I__5432 (
            .O(N__35291),
            .I(N__35288));
    Span4Mux_h I__5431 (
            .O(N__35288),
            .I(N__35285));
    Odrv4 I__5430 (
            .O(N__35285),
            .I(\ALU.mult_17_4 ));
    InMux I__5429 (
            .O(N__35282),
            .I(N__35279));
    LocalMux I__5428 (
            .O(N__35279),
            .I(N__35276));
    Span4Mux_h I__5427 (
            .O(N__35276),
            .I(N__35273));
    Span4Mux_v I__5426 (
            .O(N__35273),
            .I(N__35270));
    Odrv4 I__5425 (
            .O(N__35270),
            .I(\ALU.mult_391_c_RNIEC73TZ0Z4 ));
    CascadeMux I__5424 (
            .O(N__35267),
            .I(N__35264));
    InMux I__5423 (
            .O(N__35264),
            .I(N__35261));
    LocalMux I__5422 (
            .O(N__35261),
            .I(N__35258));
    Span4Mux_h I__5421 (
            .O(N__35258),
            .I(N__35255));
    Odrv4 I__5420 (
            .O(N__35255),
            .I(\ALU.mult_17_5 ));
    InMux I__5419 (
            .O(N__35252),
            .I(N__35249));
    LocalMux I__5418 (
            .O(N__35249),
            .I(\ALU.mult_5 ));
    InMux I__5417 (
            .O(N__35246),
            .I(\ALU.mult_25_c4 ));
    InMux I__5416 (
            .O(N__35243),
            .I(N__35240));
    LocalMux I__5415 (
            .O(N__35240),
            .I(\ALU.mult_173_c_RNIO8AOZ0Z16 ));
    CascadeMux I__5414 (
            .O(N__35237),
            .I(N__35233));
    InMux I__5413 (
            .O(N__35236),
            .I(N__35230));
    InMux I__5412 (
            .O(N__35233),
            .I(N__35227));
    LocalMux I__5411 (
            .O(N__35230),
            .I(N__35222));
    LocalMux I__5410 (
            .O(N__35227),
            .I(N__35222));
    Span4Mux_h I__5409 (
            .O(N__35222),
            .I(N__35219));
    Odrv4 I__5408 (
            .O(N__35219),
            .I(\ALU.mult_17_6 ));
    InMux I__5407 (
            .O(N__35216),
            .I(\ALU.mult_25_c5 ));
    InMux I__5406 (
            .O(N__35213),
            .I(N__35210));
    LocalMux I__5405 (
            .O(N__35210),
            .I(\ALU.mult_19_7 ));
    CascadeMux I__5404 (
            .O(N__35207),
            .I(N__35204));
    InMux I__5403 (
            .O(N__35204),
            .I(N__35201));
    LocalMux I__5402 (
            .O(N__35201),
            .I(N__35198));
    Span4Mux_h I__5401 (
            .O(N__35198),
            .I(N__35195));
    Odrv4 I__5400 (
            .O(N__35195),
            .I(\ALU.mult_17_7 ));
    InMux I__5399 (
            .O(N__35192),
            .I(\ALU.mult_25_c6 ));
    InMux I__5398 (
            .O(N__35189),
            .I(N__35186));
    LocalMux I__5397 (
            .O(N__35186),
            .I(N__35183));
    Span4Mux_h I__5396 (
            .O(N__35183),
            .I(N__35179));
    InMux I__5395 (
            .O(N__35182),
            .I(N__35176));
    Odrv4 I__5394 (
            .O(N__35179),
            .I(\CONTROL.N_350_1 ));
    LocalMux I__5393 (
            .O(N__35176),
            .I(\CONTROL.N_350_1 ));
    InMux I__5392 (
            .O(N__35171),
            .I(N__35168));
    LocalMux I__5391 (
            .O(N__35168),
            .I(N__35165));
    Span4Mux_h I__5390 (
            .O(N__35165),
            .I(N__35162));
    Span4Mux_v I__5389 (
            .O(N__35162),
            .I(N__35159));
    Odrv4 I__5388 (
            .O(N__35159),
            .I(\CONTROL.N_345 ));
    InMux I__5387 (
            .O(N__35156),
            .I(N__35153));
    LocalMux I__5386 (
            .O(N__35153),
            .I(N__35150));
    Span4Mux_v I__5385 (
            .O(N__35150),
            .I(N__35147));
    Span4Mux_h I__5384 (
            .O(N__35147),
            .I(N__35144));
    Odrv4 I__5383 (
            .O(N__35144),
            .I(\CONTROL.N_346 ));
    InMux I__5382 (
            .O(N__35141),
            .I(N__35138));
    LocalMux I__5381 (
            .O(N__35138),
            .I(N__35135));
    Span4Mux_v I__5380 (
            .O(N__35135),
            .I(N__35131));
    InMux I__5379 (
            .O(N__35134),
            .I(N__35128));
    Span4Mux_h I__5378 (
            .O(N__35131),
            .I(N__35125));
    LocalMux I__5377 (
            .O(N__35128),
            .I(\CONTROL.N_255 ));
    Odrv4 I__5376 (
            .O(N__35125),
            .I(\CONTROL.N_255 ));
    CascadeMux I__5375 (
            .O(N__35120),
            .I(\CONTROL.N_345_cascade_ ));
    IoInMux I__5374 (
            .O(N__35117),
            .I(N__35114));
    LocalMux I__5373 (
            .O(N__35114),
            .I(N__35109));
    IoInMux I__5372 (
            .O(N__35113),
            .I(N__35106));
    IoInMux I__5371 (
            .O(N__35112),
            .I(N__35103));
    IoSpan4Mux I__5370 (
            .O(N__35109),
            .I(N__35090));
    LocalMux I__5369 (
            .O(N__35106),
            .I(N__35090));
    LocalMux I__5368 (
            .O(N__35103),
            .I(N__35090));
    IoInMux I__5367 (
            .O(N__35102),
            .I(N__35087));
    IoInMux I__5366 (
            .O(N__35101),
            .I(N__35084));
    IoInMux I__5365 (
            .O(N__35100),
            .I(N__35081));
    IoInMux I__5364 (
            .O(N__35099),
            .I(N__35078));
    IoInMux I__5363 (
            .O(N__35098),
            .I(N__35075));
    IoInMux I__5362 (
            .O(N__35097),
            .I(N__35072));
    IoSpan4Mux I__5361 (
            .O(N__35090),
            .I(N__35056));
    LocalMux I__5360 (
            .O(N__35087),
            .I(N__35056));
    LocalMux I__5359 (
            .O(N__35084),
            .I(N__35056));
    LocalMux I__5358 (
            .O(N__35081),
            .I(N__35056));
    LocalMux I__5357 (
            .O(N__35078),
            .I(N__35056));
    LocalMux I__5356 (
            .O(N__35075),
            .I(N__35056));
    LocalMux I__5355 (
            .O(N__35072),
            .I(N__35056));
    IoInMux I__5354 (
            .O(N__35071),
            .I(N__35053));
    IoSpan4Mux I__5353 (
            .O(N__35056),
            .I(N__35045));
    LocalMux I__5352 (
            .O(N__35053),
            .I(N__35045));
    IoInMux I__5351 (
            .O(N__35052),
            .I(N__35042));
    IoInMux I__5350 (
            .O(N__35051),
            .I(N__35039));
    IoInMux I__5349 (
            .O(N__35050),
            .I(N__35036));
    IoSpan4Mux I__5348 (
            .O(N__35045),
            .I(N__35027));
    LocalMux I__5347 (
            .O(N__35042),
            .I(N__35027));
    LocalMux I__5346 (
            .O(N__35039),
            .I(N__35027));
    LocalMux I__5345 (
            .O(N__35036),
            .I(N__35027));
    IoSpan4Mux I__5344 (
            .O(N__35027),
            .I(N__35022));
    IoInMux I__5343 (
            .O(N__35026),
            .I(N__35019));
    IoInMux I__5342 (
            .O(N__35025),
            .I(N__35016));
    Span4Mux_s0_h I__5341 (
            .O(N__35022),
            .I(N__35013));
    LocalMux I__5340 (
            .O(N__35019),
            .I(N__35008));
    LocalMux I__5339 (
            .O(N__35016),
            .I(N__35008));
    Span4Mux_h I__5338 (
            .O(N__35013),
            .I(N__35002));
    IoSpan4Mux I__5337 (
            .O(N__35008),
            .I(N__35002));
    IoInMux I__5336 (
            .O(N__35007),
            .I(N__34999));
    Span4Mux_s0_h I__5335 (
            .O(N__35002),
            .I(N__34996));
    LocalMux I__5334 (
            .O(N__34999),
            .I(N__34991));
    Sp12to4 I__5333 (
            .O(N__34996),
            .I(N__34991));
    Span12Mux_s8_h I__5332 (
            .O(N__34991),
            .I(N__34986));
    InMux I__5331 (
            .O(N__34990),
            .I(N__34981));
    InMux I__5330 (
            .O(N__34989),
            .I(N__34981));
    Span12Mux_v I__5329 (
            .O(N__34986),
            .I(N__34978));
    LocalMux I__5328 (
            .O(N__34981),
            .I(N__34975));
    Odrv12 I__5327 (
            .O(N__34978),
            .I(ramWrite));
    Odrv12 I__5326 (
            .O(N__34975),
            .I(ramWrite));
    CEMux I__5325 (
            .O(N__34970),
            .I(N__34967));
    LocalMux I__5324 (
            .O(N__34967),
            .I(N__34961));
    CEMux I__5323 (
            .O(N__34966),
            .I(N__34958));
    CEMux I__5322 (
            .O(N__34965),
            .I(N__34955));
    CEMux I__5321 (
            .O(N__34964),
            .I(N__34951));
    Span4Mux_h I__5320 (
            .O(N__34961),
            .I(N__34946));
    LocalMux I__5319 (
            .O(N__34958),
            .I(N__34946));
    LocalMux I__5318 (
            .O(N__34955),
            .I(N__34943));
    CEMux I__5317 (
            .O(N__34954),
            .I(N__34940));
    LocalMux I__5316 (
            .O(N__34951),
            .I(N__34937));
    Span4Mux_h I__5315 (
            .O(N__34946),
            .I(N__34930));
    Span4Mux_v I__5314 (
            .O(N__34943),
            .I(N__34930));
    LocalMux I__5313 (
            .O(N__34940),
            .I(N__34930));
    Span4Mux_h I__5312 (
            .O(N__34937),
            .I(N__34927));
    Span4Mux_v I__5311 (
            .O(N__34930),
            .I(N__34924));
    Odrv4 I__5310 (
            .O(N__34927),
            .I(\CONTROL.un1_busState114_1_0Z0Z_0 ));
    Odrv4 I__5309 (
            .O(N__34924),
            .I(\CONTROL.un1_busState114_1_0Z0Z_0 ));
    InMux I__5308 (
            .O(N__34919),
            .I(N__34916));
    LocalMux I__5307 (
            .O(N__34916),
            .I(N__34913));
    Span4Mux_v I__5306 (
            .O(N__34913),
            .I(N__34910));
    Span4Mux_h I__5305 (
            .O(N__34910),
            .I(N__34907));
    Span4Mux_v I__5304 (
            .O(N__34907),
            .I(N__34903));
    InMux I__5303 (
            .O(N__34906),
            .I(N__34900));
    Odrv4 I__5302 (
            .O(N__34903),
            .I(\CONTROL.ctrlOut_10 ));
    LocalMux I__5301 (
            .O(N__34900),
            .I(\CONTROL.ctrlOut_10 ));
    InMux I__5300 (
            .O(N__34895),
            .I(N__34892));
    LocalMux I__5299 (
            .O(N__34892),
            .I(N__34889));
    Odrv4 I__5298 (
            .O(N__34889),
            .I(\CONTROL.dout_reto_10 ));
    CascadeMux I__5297 (
            .O(N__34886),
            .I(\PROM.ROMDATA.m1_cascade_ ));
    InMux I__5296 (
            .O(N__34883),
            .I(N__34880));
    LocalMux I__5295 (
            .O(N__34880),
            .I(\CONTROL.N_339 ));
    CascadeMux I__5294 (
            .O(N__34877),
            .I(\CONTROL.N_219_cascade_ ));
    CascadeMux I__5293 (
            .O(N__34874),
            .I(\CONTROL.m28_0_120_i_i_a2_0_0_cascade_ ));
    CascadeMux I__5292 (
            .O(N__34871),
            .I(\CONTROL.busState_1_RNO_1Z0Z_1_cascade_ ));
    InMux I__5291 (
            .O(N__34868),
            .I(N__34865));
    LocalMux I__5290 (
            .O(N__34865),
            .I(N__34862));
    Span4Mux_h I__5289 (
            .O(N__34862),
            .I(N__34859));
    Odrv4 I__5288 (
            .O(N__34859),
            .I(\CONTROL.busState_1_RNO_0Z0Z_1 ));
    InMux I__5287 (
            .O(N__34856),
            .I(N__34853));
    LocalMux I__5286 (
            .O(N__34853),
            .I(N__34850));
    Odrv4 I__5285 (
            .O(N__34850),
            .I(\CONTROL.g0_3_i_1_1 ));
    InMux I__5284 (
            .O(N__34847),
            .I(N__34844));
    LocalMux I__5283 (
            .O(N__34844),
            .I(N__34841));
    Span4Mux_v I__5282 (
            .O(N__34841),
            .I(N__34838));
    Span4Mux_h I__5281 (
            .O(N__34838),
            .I(N__34835));
    Sp12to4 I__5280 (
            .O(N__34835),
            .I(N__34832));
    Odrv12 I__5279 (
            .O(N__34832),
            .I(gpuOut_c_2));
    InMux I__5278 (
            .O(N__34829),
            .I(N__34826));
    LocalMux I__5277 (
            .O(N__34826),
            .I(\CONTROL.N_163 ));
    InMux I__5276 (
            .O(N__34823),
            .I(N__34820));
    LocalMux I__5275 (
            .O(N__34820),
            .I(\CONTROL.g0_3_i_2_1 ));
    InMux I__5274 (
            .O(N__34817),
            .I(N__34811));
    InMux I__5273 (
            .O(N__34816),
            .I(N__34811));
    LocalMux I__5272 (
            .O(N__34811),
            .I(\CONTROL.un1_addrstackptr_c3_0 ));
    InMux I__5271 (
            .O(N__34808),
            .I(N__34802));
    InMux I__5270 (
            .O(N__34807),
            .I(N__34802));
    LocalMux I__5269 (
            .O(N__34802),
            .I(N__34799));
    Span4Mux_h I__5268 (
            .O(N__34799),
            .I(N__34796));
    Span4Mux_v I__5267 (
            .O(N__34796),
            .I(N__34792));
    CascadeMux I__5266 (
            .O(N__34795),
            .I(N__34789));
    Span4Mux_v I__5265 (
            .O(N__34792),
            .I(N__34786));
    InMux I__5264 (
            .O(N__34789),
            .I(N__34783));
    Odrv4 I__5263 (
            .O(N__34786),
            .I(\CONTROL.addrstack_1_3 ));
    LocalMux I__5262 (
            .O(N__34783),
            .I(\CONTROL.addrstack_1_3 ));
    InMux I__5261 (
            .O(N__34778),
            .I(N__34775));
    LocalMux I__5260 (
            .O(N__34775),
            .I(\CONTROL.N_5 ));
    InMux I__5259 (
            .O(N__34772),
            .I(N__34765));
    InMux I__5258 (
            .O(N__34771),
            .I(N__34762));
    InMux I__5257 (
            .O(N__34770),
            .I(N__34757));
    InMux I__5256 (
            .O(N__34769),
            .I(N__34757));
    InMux I__5255 (
            .O(N__34768),
            .I(N__34754));
    LocalMux I__5254 (
            .O(N__34765),
            .I(N__34750));
    LocalMux I__5253 (
            .O(N__34762),
            .I(N__34743));
    LocalMux I__5252 (
            .O(N__34757),
            .I(N__34743));
    LocalMux I__5251 (
            .O(N__34754),
            .I(N__34743));
    CascadeMux I__5250 (
            .O(N__34753),
            .I(N__34740));
    Span4Mux_h I__5249 (
            .O(N__34750),
            .I(N__34736));
    Span4Mux_v I__5248 (
            .O(N__34743),
            .I(N__34733));
    InMux I__5247 (
            .O(N__34740),
            .I(N__34728));
    InMux I__5246 (
            .O(N__34739),
            .I(N__34728));
    Span4Mux_h I__5245 (
            .O(N__34736),
            .I(N__34725));
    Sp12to4 I__5244 (
            .O(N__34733),
            .I(N__34722));
    LocalMux I__5243 (
            .O(N__34728),
            .I(\CONTROL.addrstackptrZ0Z_3 ));
    Odrv4 I__5242 (
            .O(N__34725),
            .I(\CONTROL.addrstackptrZ0Z_3 ));
    Odrv12 I__5241 (
            .O(N__34722),
            .I(\CONTROL.addrstackptrZ0Z_3 ));
    CascadeMux I__5240 (
            .O(N__34715),
            .I(\CONTROL.N_83_0_cascade_ ));
    InMux I__5239 (
            .O(N__34712),
            .I(N__34709));
    LocalMux I__5238 (
            .O(N__34709),
            .I(\CONTROL.m28_0_120_i_i_4 ));
    InMux I__5237 (
            .O(N__34706),
            .I(N__34703));
    LocalMux I__5236 (
            .O(N__34703),
            .I(\CONTROL.N_75_0 ));
    CascadeMux I__5235 (
            .O(N__34700),
            .I(\CONTROL.N_75_0_cascade_ ));
    InMux I__5234 (
            .O(N__34697),
            .I(N__34694));
    LocalMux I__5233 (
            .O(N__34694),
            .I(N__34691));
    Odrv4 I__5232 (
            .O(N__34691),
            .I(\CONTROL.m38_i_2 ));
    CascadeMux I__5231 (
            .O(N__34688),
            .I(\ALU.c_RNIJMOB4_0Z0Z_1_cascade_ ));
    InMux I__5230 (
            .O(N__34685),
            .I(N__34682));
    LocalMux I__5229 (
            .O(N__34682),
            .I(N__34678));
    InMux I__5228 (
            .O(N__34681),
            .I(N__34675));
    Sp12to4 I__5227 (
            .O(N__34678),
            .I(N__34670));
    LocalMux I__5226 (
            .O(N__34675),
            .I(N__34670));
    Odrv12 I__5225 (
            .O(N__34670),
            .I(\ALU.d_RNID42JAZ0Z_1 ));
    InMux I__5224 (
            .O(N__34667),
            .I(N__34664));
    LocalMux I__5223 (
            .O(N__34664),
            .I(\ALU.operand2_6_ns_1_1 ));
    InMux I__5222 (
            .O(N__34661),
            .I(N__34658));
    LocalMux I__5221 (
            .O(N__34658),
            .I(\ALU.N_1246 ));
    CascadeMux I__5220 (
            .O(N__34655),
            .I(\ALU.operand2_3_ns_1_1_cascade_ ));
    InMux I__5219 (
            .O(N__34652),
            .I(N__34649));
    LocalMux I__5218 (
            .O(N__34649),
            .I(\ALU.N_1198 ));
    InMux I__5217 (
            .O(N__34646),
            .I(N__34640));
    InMux I__5216 (
            .O(N__34645),
            .I(N__34640));
    LocalMux I__5215 (
            .O(N__34640),
            .I(\ALU.combOperand2_d_bmZ0Z_1 ));
    CascadeMux I__5214 (
            .O(N__34637),
            .I(\ALU.N_1198_cascade_ ));
    InMux I__5213 (
            .O(N__34634),
            .I(N__34631));
    LocalMux I__5212 (
            .O(N__34631),
            .I(\ALU.c_RNIJMOB4Z0Z_1 ));
    InMux I__5211 (
            .O(N__34628),
            .I(N__34625));
    LocalMux I__5210 (
            .O(N__34625),
            .I(\CONTROL.g0_3_i_a7_2_1 ));
    CascadeMux I__5209 (
            .O(N__34622),
            .I(\CONTROL.N_5_cascade_ ));
    CascadeMux I__5208 (
            .O(N__34619),
            .I(N__34616));
    InMux I__5207 (
            .O(N__34616),
            .I(N__34613));
    LocalMux I__5206 (
            .O(N__34613),
            .I(N__34610));
    Span4Mux_v I__5205 (
            .O(N__34610),
            .I(N__34607));
    Span4Mux_h I__5204 (
            .O(N__34607),
            .I(N__34604));
    Odrv4 I__5203 (
            .O(N__34604),
            .I(\CONTROL.addrstackptr_8_3 ));
    CascadeMux I__5202 (
            .O(N__34601),
            .I(\ALU.dout_3_ns_1_3_cascade_ ));
    InMux I__5201 (
            .O(N__34598),
            .I(N__34595));
    LocalMux I__5200 (
            .O(N__34595),
            .I(\ALU.N_1136 ));
    CascadeMux I__5199 (
            .O(N__34592),
            .I(\ALU.N_1088_cascade_ ));
    CascadeMux I__5198 (
            .O(N__34589),
            .I(aluOut_3_cascade_));
    InMux I__5197 (
            .O(N__34586),
            .I(N__34583));
    LocalMux I__5196 (
            .O(N__34583),
            .I(N__34580));
    Span4Mux_h I__5195 (
            .O(N__34580),
            .I(N__34577));
    Span4Mux_v I__5194 (
            .O(N__34577),
            .I(N__34574));
    Odrv4 I__5193 (
            .O(N__34574),
            .I(busState_1_RNIH16V3_2));
    CascadeMux I__5192 (
            .O(N__34571),
            .I(\ALU.dout_3_ns_1_13_cascade_ ));
    InMux I__5191 (
            .O(N__34568),
            .I(N__34562));
    InMux I__5190 (
            .O(N__34567),
            .I(N__34562));
    LocalMux I__5189 (
            .O(N__34562),
            .I(N__34553));
    InMux I__5188 (
            .O(N__34561),
            .I(N__34548));
    InMux I__5187 (
            .O(N__34560),
            .I(N__34548));
    InMux I__5186 (
            .O(N__34559),
            .I(N__34543));
    InMux I__5185 (
            .O(N__34558),
            .I(N__34543));
    InMux I__5184 (
            .O(N__34557),
            .I(N__34537));
    InMux I__5183 (
            .O(N__34556),
            .I(N__34537));
    Span4Mux_h I__5182 (
            .O(N__34553),
            .I(N__34534));
    LocalMux I__5181 (
            .O(N__34548),
            .I(N__34531));
    LocalMux I__5180 (
            .O(N__34543),
            .I(N__34528));
    InMux I__5179 (
            .O(N__34542),
            .I(N__34525));
    LocalMux I__5178 (
            .O(N__34537),
            .I(N__34518));
    Span4Mux_v I__5177 (
            .O(N__34534),
            .I(N__34518));
    Span4Mux_h I__5176 (
            .O(N__34531),
            .I(N__34518));
    Odrv4 I__5175 (
            .O(N__34528),
            .I(aluOperand1_2_rep2));
    LocalMux I__5174 (
            .O(N__34525),
            .I(aluOperand1_2_rep2));
    Odrv4 I__5173 (
            .O(N__34518),
            .I(aluOperand1_2_rep2));
    CascadeMux I__5172 (
            .O(N__34511),
            .I(\ALU.dout_6_ns_1_13_cascade_ ));
    InMux I__5171 (
            .O(N__34508),
            .I(N__34505));
    LocalMux I__5170 (
            .O(N__34505),
            .I(\ALU.N_1098 ));
    CascadeMux I__5169 (
            .O(N__34502),
            .I(\ALU.N_1146_cascade_ ));
    InMux I__5168 (
            .O(N__34499),
            .I(N__34496));
    LocalMux I__5167 (
            .O(N__34496),
            .I(N__34493));
    Odrv4 I__5166 (
            .O(N__34493),
            .I(\CONTROL.N_190 ));
    InMux I__5165 (
            .O(N__34490),
            .I(N__34487));
    LocalMux I__5164 (
            .O(N__34487),
            .I(N__34484));
    Span4Mux_h I__5163 (
            .O(N__34484),
            .I(N__34478));
    InMux I__5162 (
            .O(N__34483),
            .I(N__34475));
    InMux I__5161 (
            .O(N__34482),
            .I(N__34472));
    InMux I__5160 (
            .O(N__34481),
            .I(N__34469));
    Odrv4 I__5159 (
            .O(N__34478),
            .I(\CONTROL.bus_7_a1_1_8 ));
    LocalMux I__5158 (
            .O(N__34475),
            .I(\CONTROL.bus_7_a1_1_8 ));
    LocalMux I__5157 (
            .O(N__34472),
            .I(\CONTROL.bus_7_a1_1_8 ));
    LocalMux I__5156 (
            .O(N__34469),
            .I(\CONTROL.bus_7_a1_1_8 ));
    CascadeMux I__5155 (
            .O(N__34460),
            .I(aluOut_13_cascade_));
    InMux I__5154 (
            .O(N__34457),
            .I(N__34451));
    InMux I__5153 (
            .O(N__34456),
            .I(N__34451));
    LocalMux I__5152 (
            .O(N__34451),
            .I(N__34448));
    Span4Mux_h I__5151 (
            .O(N__34448),
            .I(N__34445));
    Odrv4 I__5150 (
            .O(N__34445),
            .I(\CONTROL.bus_0_13 ));
    CascadeMux I__5149 (
            .O(N__34442),
            .I(\PROM.ROMDATA.m238_am_1_cascade_ ));
    CascadeMux I__5148 (
            .O(N__34439),
            .I(\PROM.ROMDATA.m238_am_cascade_ ));
    CascadeMux I__5147 (
            .O(N__34436),
            .I(\PROM.ROMDATA.m244_ns_1_cascade_ ));
    CascadeMux I__5146 (
            .O(N__34433),
            .I(N__34429));
    CascadeMux I__5145 (
            .O(N__34432),
            .I(N__34424));
    InMux I__5144 (
            .O(N__34429),
            .I(N__34421));
    InMux I__5143 (
            .O(N__34428),
            .I(N__34414));
    InMux I__5142 (
            .O(N__34427),
            .I(N__34414));
    InMux I__5141 (
            .O(N__34424),
            .I(N__34414));
    LocalMux I__5140 (
            .O(N__34421),
            .I(\PROM.ROMDATA.m244_ns_1 ));
    LocalMux I__5139 (
            .O(N__34414),
            .I(\PROM.ROMDATA.m244_ns_1 ));
    CascadeMux I__5138 (
            .O(N__34409),
            .I(\ALU.dout_6_ns_1_3_cascade_ ));
    CascadeMux I__5137 (
            .O(N__34406),
            .I(aluOut_9_cascade_));
    CascadeMux I__5136 (
            .O(N__34403),
            .I(N__34400));
    InMux I__5135 (
            .O(N__34400),
            .I(N__34396));
    CascadeMux I__5134 (
            .O(N__34399),
            .I(N__34393));
    LocalMux I__5133 (
            .O(N__34396),
            .I(N__34389));
    InMux I__5132 (
            .O(N__34393),
            .I(N__34386));
    InMux I__5131 (
            .O(N__34392),
            .I(N__34383));
    Span4Mux_h I__5130 (
            .O(N__34389),
            .I(N__34380));
    LocalMux I__5129 (
            .O(N__34386),
            .I(N__34377));
    LocalMux I__5128 (
            .O(N__34383),
            .I(N__34374));
    Span4Mux_v I__5127 (
            .O(N__34380),
            .I(N__34371));
    Span4Mux_v I__5126 (
            .O(N__34377),
            .I(N__34366));
    Span4Mux_h I__5125 (
            .O(N__34374),
            .I(N__34366));
    Span4Mux_v I__5124 (
            .O(N__34371),
            .I(N__34363));
    Span4Mux_v I__5123 (
            .O(N__34366),
            .I(N__34360));
    Odrv4 I__5122 (
            .O(N__34363),
            .I(h_2));
    Odrv4 I__5121 (
            .O(N__34360),
            .I(h_2));
    CascadeMux I__5120 (
            .O(N__34355),
            .I(\ALU.dout_6_ns_1_2_cascade_ ));
    InMux I__5119 (
            .O(N__34352),
            .I(N__34349));
    LocalMux I__5118 (
            .O(N__34349),
            .I(N__34345));
    InMux I__5117 (
            .O(N__34348),
            .I(N__34342));
    Span4Mux_v I__5116 (
            .O(N__34345),
            .I(N__34337));
    LocalMux I__5115 (
            .O(N__34342),
            .I(N__34337));
    Odrv4 I__5114 (
            .O(N__34337),
            .I(\ALU.aZ0Z_2 ));
    CascadeMux I__5113 (
            .O(N__34334),
            .I(N__34330));
    CascadeMux I__5112 (
            .O(N__34333),
            .I(N__34327));
    InMux I__5111 (
            .O(N__34330),
            .I(N__34324));
    InMux I__5110 (
            .O(N__34327),
            .I(N__34321));
    LocalMux I__5109 (
            .O(N__34324),
            .I(N__34318));
    LocalMux I__5108 (
            .O(N__34321),
            .I(N__34315));
    Odrv12 I__5107 (
            .O(N__34318),
            .I(\ALU.eZ0Z_2 ));
    Odrv4 I__5106 (
            .O(N__34315),
            .I(\ALU.eZ0Z_2 ));
    CascadeMux I__5105 (
            .O(N__34310),
            .I(\ALU.dout_3_ns_1_2_cascade_ ));
    CascadeMux I__5104 (
            .O(N__34307),
            .I(\ALU.N_1087_cascade_ ));
    InMux I__5103 (
            .O(N__34304),
            .I(N__34301));
    LocalMux I__5102 (
            .O(N__34301),
            .I(\ALU.N_1135 ));
    InMux I__5101 (
            .O(N__34298),
            .I(N__34294));
    InMux I__5100 (
            .O(N__34297),
            .I(N__34291));
    LocalMux I__5099 (
            .O(N__34294),
            .I(ALU_N_1086));
    LocalMux I__5098 (
            .O(N__34291),
            .I(ALU_N_1086));
    InMux I__5097 (
            .O(N__34286),
            .I(N__34283));
    LocalMux I__5096 (
            .O(N__34283),
            .I(\CONTROL.operand1_ne_RNIBQE03_0Z0Z_0 ));
    CascadeMux I__5095 (
            .O(N__34280),
            .I(\ALU.addsub_cry_1_c_RNIJP8KZ0Z37_cascade_ ));
    InMux I__5094 (
            .O(N__34277),
            .I(N__34274));
    LocalMux I__5093 (
            .O(N__34274),
            .I(\ALU.addsub_cry_1_c_RNIJP8KZ0Z37 ));
    CascadeMux I__5092 (
            .O(N__34271),
            .I(\ALU.addsub_cry_1_c_RNIICPECZ0Z7_cascade_ ));
    CascadeMux I__5091 (
            .O(N__34268),
            .I(\ALU.dout_3_ns_1_9_cascade_ ));
    CascadeMux I__5090 (
            .O(N__34265),
            .I(\ALU.dout_6_ns_1_9_cascade_ ));
    InMux I__5089 (
            .O(N__34262),
            .I(N__34259));
    LocalMux I__5088 (
            .O(N__34259),
            .I(\ALU.N_1094 ));
    CascadeMux I__5087 (
            .O(N__34256),
            .I(\ALU.N_1142_cascade_ ));
    InMux I__5086 (
            .O(N__34253),
            .I(N__34250));
    LocalMux I__5085 (
            .O(N__34250),
            .I(\ALU.mult_388_c_RNIBULDPZ0Z3 ));
    CascadeMux I__5084 (
            .O(N__34247),
            .I(\ALU.mult_388_c_RNIEAAJHZ0Z7_cascade_ ));
    IoInMux I__5083 (
            .O(N__34244),
            .I(N__34238));
    IoInMux I__5082 (
            .O(N__34243),
            .I(N__34235));
    InMux I__5081 (
            .O(N__34242),
            .I(N__34230));
    InMux I__5080 (
            .O(N__34241),
            .I(N__34230));
    LocalMux I__5079 (
            .O(N__34238),
            .I(N__34227));
    LocalMux I__5078 (
            .O(N__34235),
            .I(N__34224));
    LocalMux I__5077 (
            .O(N__34230),
            .I(N__34221));
    Span12Mux_s6_h I__5076 (
            .O(N__34227),
            .I(N__34218));
    IoSpan4Mux I__5075 (
            .O(N__34224),
            .I(N__34215));
    Span4Mux_v I__5074 (
            .O(N__34221),
            .I(N__34212));
    Span12Mux_h I__5073 (
            .O(N__34218),
            .I(N__34209));
    Span4Mux_s2_h I__5072 (
            .O(N__34215),
            .I(N__34206));
    Span4Mux_v I__5071 (
            .O(N__34212),
            .I(N__34203));
    Span12Mux_v I__5070 (
            .O(N__34209),
            .I(N__34200));
    Sp12to4 I__5069 (
            .O(N__34206),
            .I(N__34197));
    Span4Mux_h I__5068 (
            .O(N__34203),
            .I(N__34194));
    Odrv12 I__5067 (
            .O(N__34200),
            .I(bus_3));
    Odrv12 I__5066 (
            .O(N__34197),
            .I(bus_3));
    Odrv4 I__5065 (
            .O(N__34194),
            .I(bus_3));
    InMux I__5064 (
            .O(N__34187),
            .I(N__34184));
    LocalMux I__5063 (
            .O(N__34184),
            .I(\ALU.mult_388_c_RNIEAAJHZ0Z7 ));
    CascadeMux I__5062 (
            .O(N__34181),
            .I(\ALU.mult_388_c_RNIPGN6QZ0Z7_cascade_ ));
    InMux I__5061 (
            .O(N__34178),
            .I(N__34174));
    InMux I__5060 (
            .O(N__34177),
            .I(N__34171));
    LocalMux I__5059 (
            .O(N__34174),
            .I(N__34168));
    LocalMux I__5058 (
            .O(N__34171),
            .I(N__34165));
    Span4Mux_h I__5057 (
            .O(N__34168),
            .I(N__34160));
    Span4Mux_v I__5056 (
            .O(N__34165),
            .I(N__34160));
    Odrv4 I__5055 (
            .O(N__34160),
            .I(\ALU.a_15_d_sZ0Z_5 ));
    CascadeMux I__5054 (
            .O(N__34157),
            .I(N__34154));
    InMux I__5053 (
            .O(N__34154),
            .I(N__34151));
    LocalMux I__5052 (
            .O(N__34151),
            .I(N__34148));
    Span4Mux_v I__5051 (
            .O(N__34148),
            .I(N__34145));
    Odrv4 I__5050 (
            .O(N__34145),
            .I(\ALU.mult_2 ));
    InMux I__5049 (
            .O(N__34142),
            .I(N__34139));
    LocalMux I__5048 (
            .O(N__34139),
            .I(N__34136));
    Odrv4 I__5047 (
            .O(N__34136),
            .I(\ALU.log_1_2 ));
    InMux I__5046 (
            .O(N__34133),
            .I(N__34129));
    InMux I__5045 (
            .O(N__34132),
            .I(N__34126));
    LocalMux I__5044 (
            .O(N__34129),
            .I(\ALU.a_15_d_sZ0Z_3 ));
    LocalMux I__5043 (
            .O(N__34126),
            .I(\ALU.a_15_d_sZ0Z_3 ));
    CascadeMux I__5042 (
            .O(N__34121),
            .I(\ALU.addsub_cry_1_c_RNI8FKPLZ0Z3_cascade_ ));
    InMux I__5041 (
            .O(N__34118),
            .I(N__34115));
    LocalMux I__5040 (
            .O(N__34115),
            .I(\ALU.mult_5_c_RNI6ET5DZ0Z3 ));
    InMux I__5039 (
            .O(N__34112),
            .I(N__34109));
    LocalMux I__5038 (
            .O(N__34109),
            .I(N__34106));
    Span4Mux_v I__5037 (
            .O(N__34106),
            .I(N__34103));
    Odrv4 I__5036 (
            .O(N__34103),
            .I(\ALU.mult_3_3 ));
    InMux I__5035 (
            .O(N__34100),
            .I(N__34096));
    InMux I__5034 (
            .O(N__34099),
            .I(N__34092));
    LocalMux I__5033 (
            .O(N__34096),
            .I(N__34089));
    InMux I__5032 (
            .O(N__34095),
            .I(N__34086));
    LocalMux I__5031 (
            .O(N__34092),
            .I(N__34083));
    Sp12to4 I__5030 (
            .O(N__34089),
            .I(N__34078));
    LocalMux I__5029 (
            .O(N__34086),
            .I(N__34078));
    Span4Mux_h I__5028 (
            .O(N__34083),
            .I(N__34075));
    Span12Mux_h I__5027 (
            .O(N__34078),
            .I(N__34072));
    Odrv4 I__5026 (
            .O(N__34075),
            .I(busState_1_RNIBS0U1_2));
    Odrv12 I__5025 (
            .O(N__34072),
            .I(busState_1_RNIBS0U1_2));
    InMux I__5024 (
            .O(N__34067),
            .I(N__34063));
    InMux I__5023 (
            .O(N__34066),
            .I(N__34060));
    LocalMux I__5022 (
            .O(N__34063),
            .I(N__34055));
    LocalMux I__5021 (
            .O(N__34060),
            .I(N__34055));
    Span4Mux_h I__5020 (
            .O(N__34055),
            .I(N__34052));
    Odrv4 I__5019 (
            .O(N__34052),
            .I(operand1_ne_RNIR8FK7_0));
    CascadeMux I__5018 (
            .O(N__34049),
            .I(\ALU.status_19_0_cascade_ ));
    InMux I__5017 (
            .O(N__34046),
            .I(N__34043));
    LocalMux I__5016 (
            .O(N__34043),
            .I(N__34040));
    Span4Mux_h I__5015 (
            .O(N__34040),
            .I(N__34037));
    Odrv4 I__5014 (
            .O(N__34037),
            .I(\ALU.mult_95_c_RNOZ0 ));
    InMux I__5013 (
            .O(N__34034),
            .I(N__34031));
    LocalMux I__5012 (
            .O(N__34031),
            .I(N__34028));
    Span4Mux_v I__5011 (
            .O(N__34028),
            .I(N__34025));
    Odrv4 I__5010 (
            .O(N__34025),
            .I(\ALU.mult_3 ));
    CascadeMux I__5009 (
            .O(N__34022),
            .I(\ALU.addsub_cry_2_c_RNIUFTGNZ0Z3_cascade_ ));
    CascadeMux I__5008 (
            .O(N__34019),
            .I(\ALU.mult_486_c_RNIPJD0IZ0Z5_cascade_ ));
    CascadeMux I__5007 (
            .O(N__34016),
            .I(N__34013));
    InMux I__5006 (
            .O(N__34013),
            .I(N__34008));
    InMux I__5005 (
            .O(N__34012),
            .I(N__34005));
    InMux I__5004 (
            .O(N__34011),
            .I(N__34002));
    LocalMux I__5003 (
            .O(N__34008),
            .I(N__33997));
    LocalMux I__5002 (
            .O(N__34005),
            .I(N__33997));
    LocalMux I__5001 (
            .O(N__34002),
            .I(N__33994));
    Span4Mux_v I__5000 (
            .O(N__33997),
            .I(N__33990));
    Span12Mux_v I__4999 (
            .O(N__33994),
            .I(N__33987));
    InMux I__4998 (
            .O(N__33993),
            .I(N__33984));
    Odrv4 I__4997 (
            .O(N__33990),
            .I(\ALU.combOperand2_0_5 ));
    Odrv12 I__4996 (
            .O(N__33987),
            .I(\ALU.combOperand2_0_5 ));
    LocalMux I__4995 (
            .O(N__33984),
            .I(\ALU.combOperand2_0_5 ));
    CascadeMux I__4994 (
            .O(N__33977),
            .I(N__33974));
    InMux I__4993 (
            .O(N__33974),
            .I(N__33971));
    LocalMux I__4992 (
            .O(N__33971),
            .I(N__33968));
    Odrv4 I__4991 (
            .O(N__33968),
            .I(\ALU.d_RNICGRJGZ0Z_1 ));
    InMux I__4990 (
            .O(N__33965),
            .I(N__33962));
    LocalMux I__4989 (
            .O(N__33962),
            .I(\ALU.addsub_cry_4_c_RNI2RZ0Z6596 ));
    CascadeMux I__4988 (
            .O(N__33959),
            .I(N__33956));
    InMux I__4987 (
            .O(N__33956),
            .I(N__33953));
    LocalMux I__4986 (
            .O(N__33953),
            .I(N__33950));
    Odrv4 I__4985 (
            .O(N__33950),
            .I(\ALU.d_RNIBVMTLZ0Z_5 ));
    InMux I__4984 (
            .O(N__33947),
            .I(N__33944));
    LocalMux I__4983 (
            .O(N__33944),
            .I(N__33941));
    Span4Mux_h I__4982 (
            .O(N__33941),
            .I(N__33938));
    Odrv4 I__4981 (
            .O(N__33938),
            .I(\ALU.d_RNIVMDLOZ0Z_5 ));
    InMux I__4980 (
            .O(N__33935),
            .I(\ALU.mult_19_c8 ));
    InMux I__4979 (
            .O(N__33932),
            .I(N__33929));
    LocalMux I__4978 (
            .O(N__33929),
            .I(N__33926));
    Odrv4 I__4977 (
            .O(N__33926),
            .I(\ALU.mult_7_10 ));
    CascadeMux I__4976 (
            .O(N__33923),
            .I(N__33920));
    InMux I__4975 (
            .O(N__33920),
            .I(N__33917));
    LocalMux I__4974 (
            .O(N__33917),
            .I(\ALU.mult_5_10 ));
    InMux I__4973 (
            .O(N__33914),
            .I(\ALU.mult_19_c9 ));
    InMux I__4972 (
            .O(N__33911),
            .I(N__33908));
    LocalMux I__4971 (
            .O(N__33908),
            .I(N__33905));
    Odrv4 I__4970 (
            .O(N__33905),
            .I(\ALU.mult_7_11 ));
    CascadeMux I__4969 (
            .O(N__33902),
            .I(N__33899));
    InMux I__4968 (
            .O(N__33899),
            .I(N__33896));
    LocalMux I__4967 (
            .O(N__33896),
            .I(N__33893));
    Odrv4 I__4966 (
            .O(N__33893),
            .I(\ALU.mult_5_11 ));
    InMux I__4965 (
            .O(N__33890),
            .I(\ALU.mult_19_c10 ));
    InMux I__4964 (
            .O(N__33887),
            .I(N__33884));
    LocalMux I__4963 (
            .O(N__33884),
            .I(\ALU.mult_5_12 ));
    CascadeMux I__4962 (
            .O(N__33881),
            .I(N__33878));
    InMux I__4961 (
            .O(N__33878),
            .I(N__33875));
    LocalMux I__4960 (
            .O(N__33875),
            .I(N__33872));
    Odrv12 I__4959 (
            .O(N__33872),
            .I(\ALU.mult_7_12 ));
    InMux I__4958 (
            .O(N__33869),
            .I(\ALU.mult_19_c11 ));
    InMux I__4957 (
            .O(N__33866),
            .I(N__33863));
    LocalMux I__4956 (
            .O(N__33863),
            .I(\ALU.mult_5_13 ));
    CascadeMux I__4955 (
            .O(N__33860),
            .I(N__33857));
    InMux I__4954 (
            .O(N__33857),
            .I(N__33854));
    LocalMux I__4953 (
            .O(N__33854),
            .I(N__33851));
    Span4Mux_h I__4952 (
            .O(N__33851),
            .I(N__33848));
    Odrv4 I__4951 (
            .O(N__33848),
            .I(\ALU.mult_7_13 ));
    InMux I__4950 (
            .O(N__33845),
            .I(\ALU.mult_19_c12 ));
    InMux I__4949 (
            .O(N__33842),
            .I(N__33839));
    LocalMux I__4948 (
            .O(N__33839),
            .I(\ALU.mult_5_14 ));
    CascadeMux I__4947 (
            .O(N__33836),
            .I(N__33833));
    InMux I__4946 (
            .O(N__33833),
            .I(N__33830));
    LocalMux I__4945 (
            .O(N__33830),
            .I(N__33827));
    Span4Mux_h I__4944 (
            .O(N__33827),
            .I(N__33824));
    Odrv4 I__4943 (
            .O(N__33824),
            .I(\ALU.mult_7_14 ));
    InMux I__4942 (
            .O(N__33821),
            .I(bfn_15_10_0_));
    InMux I__4941 (
            .O(N__33818),
            .I(\ALU.mult_19_c14 ));
    CascadeMux I__4940 (
            .O(N__33815),
            .I(N__33812));
    InMux I__4939 (
            .O(N__33812),
            .I(N__33809));
    LocalMux I__4938 (
            .O(N__33809),
            .I(\ALU.mult_19_c14_THRU_CO ));
    InMux I__4937 (
            .O(N__33806),
            .I(N__33803));
    LocalMux I__4936 (
            .O(N__33803),
            .I(N__33800));
    Odrv4 I__4935 (
            .O(N__33800),
            .I(\ALU.mult_3_2 ));
    CascadeMux I__4934 (
            .O(N__33797),
            .I(N__33794));
    InMux I__4933 (
            .O(N__33794),
            .I(N__33791));
    LocalMux I__4932 (
            .O(N__33791),
            .I(N__33788));
    Span4Mux_h I__4931 (
            .O(N__33788),
            .I(N__33785));
    Sp12to4 I__4930 (
            .O(N__33785),
            .I(N__33782));
    Span12Mux_v I__4929 (
            .O(N__33782),
            .I(N__33779));
    Span12Mux_v I__4928 (
            .O(N__33779),
            .I(N__33776));
    Odrv12 I__4927 (
            .O(N__33776),
            .I(\CONTROL.addrstack_1_i ));
    CascadeMux I__4926 (
            .O(N__33773),
            .I(N__33770));
    InMux I__4925 (
            .O(N__33770),
            .I(N__33767));
    LocalMux I__4924 (
            .O(N__33767),
            .I(\ALU.d_RNII2KJ41Z0Z_4 ));
    IoInMux I__4923 (
            .O(N__33764),
            .I(N__33760));
    IoInMux I__4922 (
            .O(N__33763),
            .I(N__33757));
    LocalMux I__4921 (
            .O(N__33760),
            .I(N__33754));
    LocalMux I__4920 (
            .O(N__33757),
            .I(N__33751));
    Span4Mux_s3_h I__4919 (
            .O(N__33754),
            .I(N__33748));
    Span4Mux_s3_h I__4918 (
            .O(N__33751),
            .I(N__33745));
    Span4Mux_v I__4917 (
            .O(N__33748),
            .I(N__33741));
    Span4Mux_h I__4916 (
            .O(N__33745),
            .I(N__33738));
    InMux I__4915 (
            .O(N__33744),
            .I(N__33735));
    Sp12to4 I__4914 (
            .O(N__33741),
            .I(N__33732));
    Sp12to4 I__4913 (
            .O(N__33738),
            .I(N__33729));
    LocalMux I__4912 (
            .O(N__33735),
            .I(N__33726));
    Span12Mux_h I__4911 (
            .O(N__33732),
            .I(N__33721));
    Span12Mux_v I__4910 (
            .O(N__33729),
            .I(N__33721));
    Span4Mux_h I__4909 (
            .O(N__33726),
            .I(N__33718));
    Odrv12 I__4908 (
            .O(N__33721),
            .I(bus_4));
    Odrv4 I__4907 (
            .O(N__33718),
            .I(bus_4));
    InMux I__4906 (
            .O(N__33713),
            .I(N__33710));
    LocalMux I__4905 (
            .O(N__33710),
            .I(\ALU.mult_173_c_RNOZ0 ));
    CascadeMux I__4904 (
            .O(N__33707),
            .I(N__33704));
    InMux I__4903 (
            .O(N__33704),
            .I(N__33701));
    LocalMux I__4902 (
            .O(N__33701),
            .I(\ALU.mult_5_6 ));
    InMux I__4901 (
            .O(N__33698),
            .I(N__33695));
    LocalMux I__4900 (
            .O(N__33695),
            .I(N__33692));
    Odrv12 I__4899 (
            .O(N__33692),
            .I(\ALU.mult_7_7 ));
    CascadeMux I__4898 (
            .O(N__33689),
            .I(N__33686));
    InMux I__4897 (
            .O(N__33686),
            .I(N__33683));
    LocalMux I__4896 (
            .O(N__33683),
            .I(\ALU.mult_5_7 ));
    InMux I__4895 (
            .O(N__33680),
            .I(\ALU.mult_19_c6 ));
    InMux I__4894 (
            .O(N__33677),
            .I(N__33674));
    LocalMux I__4893 (
            .O(N__33674),
            .I(N__33671));
    Span4Mux_h I__4892 (
            .O(N__33671),
            .I(N__33668));
    Odrv4 I__4891 (
            .O(N__33668),
            .I(\ALU.mult_7_8 ));
    CascadeMux I__4890 (
            .O(N__33665),
            .I(N__33662));
    InMux I__4889 (
            .O(N__33662),
            .I(N__33659));
    LocalMux I__4888 (
            .O(N__33659),
            .I(\ALU.mult_5_8 ));
    InMux I__4887 (
            .O(N__33656),
            .I(\ALU.mult_19_c7 ));
    InMux I__4886 (
            .O(N__33653),
            .I(N__33650));
    LocalMux I__4885 (
            .O(N__33650),
            .I(N__33647));
    Odrv4 I__4884 (
            .O(N__33647),
            .I(\ALU.mult_7_9 ));
    CascadeMux I__4883 (
            .O(N__33644),
            .I(N__33641));
    InMux I__4882 (
            .O(N__33641),
            .I(N__33638));
    LocalMux I__4881 (
            .O(N__33638),
            .I(\ALU.mult_5_9 ));
    InMux I__4880 (
            .O(N__33635),
            .I(N__33632));
    LocalMux I__4879 (
            .O(N__33632),
            .I(N__33629));
    Span4Mux_h I__4878 (
            .O(N__33629),
            .I(N__33626));
    Span4Mux_h I__4877 (
            .O(N__33626),
            .I(N__33623));
    Odrv4 I__4876 (
            .O(N__33623),
            .I(\CONTROL.tempCounterZ0Z_0 ));
    InMux I__4875 (
            .O(N__33620),
            .I(N__33617));
    LocalMux I__4874 (
            .O(N__33617),
            .I(N__33614));
    Sp12to4 I__4873 (
            .O(N__33614),
            .I(N__33611));
    Span12Mux_h I__4872 (
            .O(N__33611),
            .I(N__33608));
    Odrv12 I__4871 (
            .O(N__33608),
            .I(\CONTROL.tempCounterZ0Z_5 ));
    InMux I__4870 (
            .O(N__33605),
            .I(N__33602));
    LocalMux I__4869 (
            .O(N__33602),
            .I(N__33599));
    Span4Mux_h I__4868 (
            .O(N__33599),
            .I(N__33596));
    Span4Mux_h I__4867 (
            .O(N__33596),
            .I(N__33593));
    Sp12to4 I__4866 (
            .O(N__33593),
            .I(N__33590));
    Odrv12 I__4865 (
            .O(N__33590),
            .I(\CONTROL.tempCounterZ0Z_3 ));
    InMux I__4864 (
            .O(N__33587),
            .I(N__33583));
    InMux I__4863 (
            .O(N__33586),
            .I(N__33580));
    LocalMux I__4862 (
            .O(N__33583),
            .I(N__33577));
    LocalMux I__4861 (
            .O(N__33580),
            .I(N__33572));
    Span4Mux_h I__4860 (
            .O(N__33577),
            .I(N__33572));
    Odrv4 I__4859 (
            .O(N__33572),
            .I(\CONTROL.programCounter_1_8 ));
    InMux I__4858 (
            .O(N__33569),
            .I(N__33566));
    LocalMux I__4857 (
            .O(N__33566),
            .I(N__33563));
    Span4Mux_v I__4856 (
            .O(N__33563),
            .I(N__33560));
    Span4Mux_h I__4855 (
            .O(N__33560),
            .I(N__33557));
    Odrv4 I__4854 (
            .O(N__33557),
            .I(\CONTROL.tempCounterZ0Z_8 ));
    InMux I__4853 (
            .O(N__33554),
            .I(N__33551));
    LocalMux I__4852 (
            .O(N__33551),
            .I(N__33548));
    Span4Mux_h I__4851 (
            .O(N__33548),
            .I(N__33545));
    Span4Mux_h I__4850 (
            .O(N__33545),
            .I(N__33542));
    Odrv4 I__4849 (
            .O(N__33542),
            .I(\CONTROL.tempCounterZ0Z_4 ));
    InMux I__4848 (
            .O(N__33539),
            .I(N__33536));
    LocalMux I__4847 (
            .O(N__33536),
            .I(N__33533));
    Span4Mux_h I__4846 (
            .O(N__33533),
            .I(N__33530));
    Span4Mux_h I__4845 (
            .O(N__33530),
            .I(N__33527));
    Odrv4 I__4844 (
            .O(N__33527),
            .I(\CONTROL.tempCounterZ0Z_1 ));
    InMux I__4843 (
            .O(N__33524),
            .I(N__33521));
    LocalMux I__4842 (
            .O(N__33521),
            .I(N__33518));
    Span4Mux_h I__4841 (
            .O(N__33518),
            .I(N__33515));
    Span4Mux_h I__4840 (
            .O(N__33515),
            .I(N__33512));
    Odrv4 I__4839 (
            .O(N__33512),
            .I(\CONTROL.tempCounterZ0Z_7 ));
    InMux I__4838 (
            .O(N__33509),
            .I(N__33506));
    LocalMux I__4837 (
            .O(N__33506),
            .I(N__33503));
    Span4Mux_h I__4836 (
            .O(N__33503),
            .I(N__33500));
    Odrv4 I__4835 (
            .O(N__33500),
            .I(\CONTROL.tempCounterZ0Z_12 ));
    InMux I__4834 (
            .O(N__33497),
            .I(N__33494));
    LocalMux I__4833 (
            .O(N__33494),
            .I(N__33491));
    Span4Mux_v I__4832 (
            .O(N__33491),
            .I(N__33488));
    Span4Mux_h I__4831 (
            .O(N__33488),
            .I(N__33485));
    Odrv4 I__4830 (
            .O(N__33485),
            .I(\CONTROL.tempCounterZ0Z_2 ));
    InMux I__4829 (
            .O(N__33482),
            .I(N__33479));
    LocalMux I__4828 (
            .O(N__33479),
            .I(N__33476));
    Odrv4 I__4827 (
            .O(N__33476),
            .I(\CONTROL.N_430 ));
    InMux I__4826 (
            .O(N__33473),
            .I(N__33470));
    LocalMux I__4825 (
            .O(N__33470),
            .I(N__33467));
    Span4Mux_h I__4824 (
            .O(N__33467),
            .I(N__33464));
    Odrv4 I__4823 (
            .O(N__33464),
            .I(\CONTROL.un1_busState98_1_1_0Z0Z_0 ));
    InMux I__4822 (
            .O(N__33461),
            .I(N__33458));
    LocalMux I__4821 (
            .O(N__33458),
            .I(N__33454));
    InMux I__4820 (
            .O(N__33457),
            .I(N__33451));
    Span4Mux_h I__4819 (
            .O(N__33454),
            .I(N__33448));
    LocalMux I__4818 (
            .O(N__33451),
            .I(N__33445));
    Odrv4 I__4817 (
            .O(N__33448),
            .I(\CONTROL.programCounter_1_15 ));
    Odrv4 I__4816 (
            .O(N__33445),
            .I(\CONTROL.programCounter_1_15 ));
    InMux I__4815 (
            .O(N__33440),
            .I(N__33437));
    LocalMux I__4814 (
            .O(N__33437),
            .I(\CONTROL.programCounter_1_reto_15 ));
    InMux I__4813 (
            .O(N__33434),
            .I(N__33430));
    InMux I__4812 (
            .O(N__33433),
            .I(N__33427));
    LocalMux I__4811 (
            .O(N__33430),
            .I(\CONTROL.ctrlOut_15 ));
    LocalMux I__4810 (
            .O(N__33427),
            .I(\CONTROL.ctrlOut_15 ));
    InMux I__4809 (
            .O(N__33422),
            .I(N__33419));
    LocalMux I__4808 (
            .O(N__33419),
            .I(\CONTROL.dout_reto_15 ));
    InMux I__4807 (
            .O(N__33416),
            .I(N__33413));
    LocalMux I__4806 (
            .O(N__33413),
            .I(N__33410));
    Span4Mux_v I__4805 (
            .O(N__33410),
            .I(N__33407));
    Span4Mux_h I__4804 (
            .O(N__33407),
            .I(N__33404));
    Odrv4 I__4803 (
            .O(N__33404),
            .I(\PROM.ROMDATA.m465_am ));
    InMux I__4802 (
            .O(N__33401),
            .I(N__33398));
    LocalMux I__4801 (
            .O(N__33398),
            .I(N__33395));
    Span4Mux_h I__4800 (
            .O(N__33395),
            .I(N__33392));
    Span4Mux_v I__4799 (
            .O(N__33392),
            .I(N__33388));
    InMux I__4798 (
            .O(N__33391),
            .I(N__33385));
    Odrv4 I__4797 (
            .O(N__33388),
            .I(\CONTROL.ctrlOut_7 ));
    LocalMux I__4796 (
            .O(N__33385),
            .I(\CONTROL.ctrlOut_7 ));
    InMux I__4795 (
            .O(N__33380),
            .I(N__33377));
    LocalMux I__4794 (
            .O(N__33377),
            .I(\CONTROL.N_180 ));
    InMux I__4793 (
            .O(N__33374),
            .I(N__33371));
    LocalMux I__4792 (
            .O(N__33371),
            .I(N__33368));
    Span4Mux_v I__4791 (
            .O(N__33368),
            .I(N__33365));
    Span4Mux_v I__4790 (
            .O(N__33365),
            .I(N__33362));
    Span4Mux_v I__4789 (
            .O(N__33362),
            .I(N__33359));
    Span4Mux_h I__4788 (
            .O(N__33359),
            .I(N__33356));
    Odrv4 I__4787 (
            .O(N__33356),
            .I(gpuOut_c_3));
    CascadeMux I__4786 (
            .O(N__33353),
            .I(N__33350));
    InMux I__4785 (
            .O(N__33350),
            .I(N__33347));
    LocalMux I__4784 (
            .O(N__33347),
            .I(N_164));
    InMux I__4783 (
            .O(N__33344),
            .I(N__33338));
    InMux I__4782 (
            .O(N__33343),
            .I(N__33338));
    LocalMux I__4781 (
            .O(N__33338),
            .I(N__33335));
    Span4Mux_h I__4780 (
            .O(N__33335),
            .I(N__33332));
    Span4Mux_v I__4779 (
            .O(N__33332),
            .I(N__33329));
    Span4Mux_v I__4778 (
            .O(N__33329),
            .I(N__33326));
    IoSpan4Mux I__4777 (
            .O(N__33326),
            .I(N__33323));
    Odrv4 I__4776 (
            .O(N__33323),
            .I(D3_in_c));
    CascadeMux I__4775 (
            .O(N__33320),
            .I(N_164_cascade_));
    InMux I__4774 (
            .O(N__33317),
            .I(N__33314));
    LocalMux I__4773 (
            .O(N__33314),
            .I(N__33310));
    InMux I__4772 (
            .O(N__33313),
            .I(N__33307));
    Span4Mux_h I__4771 (
            .O(N__33310),
            .I(N__33301));
    LocalMux I__4770 (
            .O(N__33307),
            .I(N__33301));
    InMux I__4769 (
            .O(N__33306),
            .I(N__33298));
    Odrv4 I__4768 (
            .O(N__33301),
            .I(controlWord_16));
    LocalMux I__4767 (
            .O(N__33298),
            .I(controlWord_16));
    CascadeMux I__4766 (
            .O(N__33293),
            .I(N__33290));
    CascadeBuf I__4765 (
            .O(N__33290),
            .I(N__33287));
    CascadeMux I__4764 (
            .O(N__33287),
            .I(N__33284));
    CascadeBuf I__4763 (
            .O(N__33284),
            .I(N__33281));
    CascadeMux I__4762 (
            .O(N__33281),
            .I(N__33278));
    CascadeBuf I__4761 (
            .O(N__33278),
            .I(N__33275));
    CascadeMux I__4760 (
            .O(N__33275),
            .I(N__33272));
    InMux I__4759 (
            .O(N__33272),
            .I(N__33269));
    LocalMux I__4758 (
            .O(N__33269),
            .I(N__33266));
    Span4Mux_h I__4757 (
            .O(N__33266),
            .I(N__33263));
    Span4Mux_h I__4756 (
            .O(N__33263),
            .I(N__33260));
    Odrv4 I__4755 (
            .O(N__33260),
            .I(CONTROL_romAddReg_7_0));
    InMux I__4754 (
            .O(N__33257),
            .I(N__33254));
    LocalMux I__4753 (
            .O(N__33254),
            .I(N__33251));
    Span4Mux_h I__4752 (
            .O(N__33251),
            .I(N__33248));
    Span4Mux_h I__4751 (
            .O(N__33248),
            .I(N__33244));
    InMux I__4750 (
            .O(N__33247),
            .I(N__33241));
    Odrv4 I__4749 (
            .O(N__33244),
            .I(controlWord_17));
    LocalMux I__4748 (
            .O(N__33241),
            .I(controlWord_17));
    CascadeMux I__4747 (
            .O(N__33236),
            .I(controlWord_17_cascade_));
    CascadeMux I__4746 (
            .O(N__33233),
            .I(N__33230));
    CascadeBuf I__4745 (
            .O(N__33230),
            .I(N__33227));
    CascadeMux I__4744 (
            .O(N__33227),
            .I(N__33224));
    CascadeBuf I__4743 (
            .O(N__33224),
            .I(N__33221));
    CascadeMux I__4742 (
            .O(N__33221),
            .I(N__33218));
    CascadeBuf I__4741 (
            .O(N__33218),
            .I(N__33215));
    CascadeMux I__4740 (
            .O(N__33215),
            .I(N__33212));
    InMux I__4739 (
            .O(N__33212),
            .I(N__33209));
    LocalMux I__4738 (
            .O(N__33209),
            .I(N__33206));
    Span12Mux_s10_v I__4737 (
            .O(N__33206),
            .I(N__33203));
    Odrv12 I__4736 (
            .O(N__33203),
            .I(CONTROL_romAddReg_7_1));
    InMux I__4735 (
            .O(N__33200),
            .I(N__33197));
    LocalMux I__4734 (
            .O(N__33197),
            .I(N__33194));
    Odrv4 I__4733 (
            .O(N__33194),
            .I(\CONTROL.N_169 ));
    CascadeMux I__4732 (
            .O(N__33191),
            .I(N__33188));
    InMux I__4731 (
            .O(N__33188),
            .I(N__33185));
    LocalMux I__4730 (
            .O(N__33185),
            .I(N__33182));
    Span4Mux_v I__4729 (
            .O(N__33182),
            .I(N__33179));
    Span4Mux_v I__4728 (
            .O(N__33179),
            .I(N__33176));
    Sp12to4 I__4727 (
            .O(N__33176),
            .I(N__33173));
    Span12Mux_h I__4726 (
            .O(N__33173),
            .I(N__33170));
    Odrv12 I__4725 (
            .O(N__33170),
            .I(D8_in_c));
    InMux I__4724 (
            .O(N__33167),
            .I(N__33163));
    InMux I__4723 (
            .O(N__33166),
            .I(N__33160));
    LocalMux I__4722 (
            .O(N__33163),
            .I(N__33157));
    LocalMux I__4721 (
            .O(N__33160),
            .I(N__33154));
    Span4Mux_v I__4720 (
            .O(N__33157),
            .I(N__33151));
    Span4Mux_h I__4719 (
            .O(N__33154),
            .I(N__33148));
    Odrv4 I__4718 (
            .O(N__33151),
            .I(\CONTROL.N_185 ));
    Odrv4 I__4717 (
            .O(N__33148),
            .I(\CONTROL.N_185 ));
    CascadeMux I__4716 (
            .O(N__33143),
            .I(N__33140));
    InMux I__4715 (
            .O(N__33140),
            .I(N__33136));
    CascadeMux I__4714 (
            .O(N__33139),
            .I(N__33133));
    LocalMux I__4713 (
            .O(N__33136),
            .I(N__33130));
    InMux I__4712 (
            .O(N__33133),
            .I(N__33127));
    Span4Mux_v I__4711 (
            .O(N__33130),
            .I(N__33124));
    LocalMux I__4710 (
            .O(N__33127),
            .I(N__33121));
    Span4Mux_v I__4709 (
            .O(N__33124),
            .I(N__33116));
    Span4Mux_v I__4708 (
            .O(N__33121),
            .I(N__33116));
    Span4Mux_h I__4707 (
            .O(N__33116),
            .I(N__33113));
    Span4Mux_h I__4706 (
            .O(N__33113),
            .I(N__33110));
    Sp12to4 I__4705 (
            .O(N__33110),
            .I(N__33107));
    Span12Mux_v I__4704 (
            .O(N__33107),
            .I(N__33104));
    Odrv12 I__4703 (
            .O(N__33104),
            .I(D4_in_c));
    InMux I__4702 (
            .O(N__33101),
            .I(N__33098));
    LocalMux I__4701 (
            .O(N__33098),
            .I(N__33095));
    Span12Mux_h I__4700 (
            .O(N__33095),
            .I(N__33092));
    Span12Mux_v I__4699 (
            .O(N__33092),
            .I(N__33089));
    Odrv12 I__4698 (
            .O(N__33089),
            .I(\CONTROL.busState_1_RNIU83C1_0Z0Z_2 ));
    CascadeMux I__4697 (
            .O(N__33086),
            .I(N__33083));
    InMux I__4696 (
            .O(N__33083),
            .I(N__33080));
    LocalMux I__4695 (
            .O(N__33080),
            .I(N__33077));
    Span4Mux_v I__4694 (
            .O(N__33077),
            .I(N__33074));
    Sp12to4 I__4693 (
            .O(N__33074),
            .I(N__33071));
    Span12Mux_h I__4692 (
            .O(N__33071),
            .I(N__33068));
    Odrv12 I__4691 (
            .O(N__33068),
            .I(D2_in_c));
    InMux I__4690 (
            .O(N__33065),
            .I(N__33062));
    LocalMux I__4689 (
            .O(N__33062),
            .I(N__33059));
    Span4Mux_v I__4688 (
            .O(N__33059),
            .I(N__33054));
    InMux I__4687 (
            .O(N__33058),
            .I(N__33051));
    CascadeMux I__4686 (
            .O(N__33057),
            .I(N__33048));
    Span4Mux_v I__4685 (
            .O(N__33054),
            .I(N__33043));
    LocalMux I__4684 (
            .O(N__33051),
            .I(N__33043));
    InMux I__4683 (
            .O(N__33048),
            .I(N__33040));
    Span4Mux_h I__4682 (
            .O(N__33043),
            .I(N__33037));
    LocalMux I__4681 (
            .O(N__33040),
            .I(N_228_0));
    Odrv4 I__4680 (
            .O(N__33037),
            .I(N_228_0));
    InMux I__4679 (
            .O(N__33032),
            .I(N__33029));
    LocalMux I__4678 (
            .O(N__33029),
            .I(N__33026));
    Span4Mux_v I__4677 (
            .O(N__33026),
            .I(N__33023));
    Sp12to4 I__4676 (
            .O(N__33023),
            .I(N__33020));
    Odrv12 I__4675 (
            .O(N__33020),
            .I(\CONTROL.busState_1_RNILAEH1Z0Z_2 ));
    InMux I__4674 (
            .O(N__33017),
            .I(N__33014));
    LocalMux I__4673 (
            .O(N__33014),
            .I(N__33011));
    Span4Mux_v I__4672 (
            .O(N__33011),
            .I(N__33008));
    Span4Mux_v I__4671 (
            .O(N__33008),
            .I(N__33005));
    Span4Mux_v I__4670 (
            .O(N__33005),
            .I(N__33002));
    Span4Mux_h I__4669 (
            .O(N__33002),
            .I(N__32999));
    IoSpan4Mux I__4668 (
            .O(N__32999),
            .I(N__32996));
    Odrv4 I__4667 (
            .O(N__32996),
            .I(gpuOut_c_1));
    CascadeMux I__4666 (
            .O(N__32993),
            .I(N__32990));
    InMux I__4665 (
            .O(N__32990),
            .I(N__32987));
    LocalMux I__4664 (
            .O(N__32987),
            .I(N_162));
    InMux I__4663 (
            .O(N__32984),
            .I(N__32978));
    InMux I__4662 (
            .O(N__32983),
            .I(N__32978));
    LocalMux I__4661 (
            .O(N__32978),
            .I(N__32975));
    Span4Mux_v I__4660 (
            .O(N__32975),
            .I(N__32972));
    Span4Mux_h I__4659 (
            .O(N__32972),
            .I(N__32969));
    Sp12to4 I__4658 (
            .O(N__32969),
            .I(N__32966));
    Odrv12 I__4657 (
            .O(N__32966),
            .I(D1_in_c));
    CascadeMux I__4656 (
            .O(N__32963),
            .I(N_162_cascade_));
    CascadeMux I__4655 (
            .O(N__32960),
            .I(\ALU.operand2_3_ns_1_2_cascade_ ));
    CascadeMux I__4654 (
            .O(N__32957),
            .I(\ALU.N_1199_cascade_ ));
    InMux I__4653 (
            .O(N__32954),
            .I(N__32951));
    LocalMux I__4652 (
            .O(N__32951),
            .I(\ALU.N_1199 ));
    CascadeMux I__4651 (
            .O(N__32948),
            .I(\ALU.c_RNIJ1JO4_0Z0Z_2_cascade_ ));
    InMux I__4650 (
            .O(N__32945),
            .I(N__32942));
    LocalMux I__4649 (
            .O(N__32942),
            .I(\ALU.c_RNIJ1JO4Z0Z_2 ));
    InMux I__4648 (
            .O(N__32939),
            .I(N__32930));
    InMux I__4647 (
            .O(N__32938),
            .I(N__32930));
    InMux I__4646 (
            .O(N__32937),
            .I(N__32930));
    LocalMux I__4645 (
            .O(N__32930),
            .I(N__32927));
    Odrv12 I__4644 (
            .O(N__32927),
            .I(\ALU.d_RNIARKGBZ0Z_2 ));
    InMux I__4643 (
            .O(N__32924),
            .I(N__32921));
    LocalMux I__4642 (
            .O(N__32921),
            .I(\ALU.operand2_6_ns_1_2 ));
    InMux I__4641 (
            .O(N__32918),
            .I(N__32915));
    LocalMux I__4640 (
            .O(N__32915),
            .I(\ALU.N_1247 ));
    InMux I__4639 (
            .O(N__32912),
            .I(N__32909));
    LocalMux I__4638 (
            .O(N__32909),
            .I(N__32906));
    Span4Mux_v I__4637 (
            .O(N__32906),
            .I(N__32903));
    Span4Mux_v I__4636 (
            .O(N__32903),
            .I(N__32900));
    Sp12to4 I__4635 (
            .O(N__32900),
            .I(N__32897));
    Span12Mux_h I__4634 (
            .O(N__32897),
            .I(N__32894));
    Odrv12 I__4633 (
            .O(N__32894),
            .I(gpuOut_c_13));
    InMux I__4632 (
            .O(N__32891),
            .I(N__32888));
    LocalMux I__4631 (
            .O(N__32888),
            .I(N__32885));
    Span4Mux_h I__4630 (
            .O(N__32885),
            .I(N__32882));
    Span4Mux_v I__4629 (
            .O(N__32882),
            .I(N__32879));
    Span4Mux_v I__4628 (
            .O(N__32879),
            .I(N__32876));
    Span4Mux_v I__4627 (
            .O(N__32876),
            .I(N__32873));
    Span4Mux_h I__4626 (
            .O(N__32873),
            .I(N__32870));
    Odrv4 I__4625 (
            .O(N__32870),
            .I(D13_in_c));
    CascadeMux I__4624 (
            .O(N__32867),
            .I(\CONTROL.N_174_cascade_ ));
    InMux I__4623 (
            .O(N__32864),
            .I(N__32861));
    LocalMux I__4622 (
            .O(N__32861),
            .I(N__32858));
    Span4Mux_v I__4621 (
            .O(N__32858),
            .I(N__32855));
    Span4Mux_v I__4620 (
            .O(N__32855),
            .I(N__32852));
    Odrv4 I__4619 (
            .O(N__32852),
            .I(\ALU.d_RNIHD7AOZ0Z_7 ));
    CascadeMux I__4618 (
            .O(N__32849),
            .I(\CONTROL.operand1_ne_RNIHKCU2Z0Z_0_cascade_ ));
    CascadeMux I__4617 (
            .O(N__32846),
            .I(N__32842));
    InMux I__4616 (
            .O(N__32845),
            .I(N__32837));
    InMux I__4615 (
            .O(N__32842),
            .I(N__32837));
    LocalMux I__4614 (
            .O(N__32837),
            .I(N__32834));
    Odrv4 I__4613 (
            .O(N__32834),
            .I(operand1_ne_RNIDN8E7_0));
    InMux I__4612 (
            .O(N__32831),
            .I(N__32828));
    LocalMux I__4611 (
            .O(N__32828),
            .I(\ALU.dout_6_ns_1_0 ));
    InMux I__4610 (
            .O(N__32825),
            .I(N__32816));
    InMux I__4609 (
            .O(N__32824),
            .I(N__32816));
    InMux I__4608 (
            .O(N__32823),
            .I(N__32811));
    InMux I__4607 (
            .O(N__32822),
            .I(N__32811));
    InMux I__4606 (
            .O(N__32821),
            .I(N__32806));
    LocalMux I__4605 (
            .O(N__32816),
            .I(N__32801));
    LocalMux I__4604 (
            .O(N__32811),
            .I(N__32801));
    InMux I__4603 (
            .O(N__32810),
            .I(N__32796));
    InMux I__4602 (
            .O(N__32809),
            .I(N__32796));
    LocalMux I__4601 (
            .O(N__32806),
            .I(aluOperand1_2_rep1));
    Odrv4 I__4600 (
            .O(N__32801),
            .I(aluOperand1_2_rep1));
    LocalMux I__4599 (
            .O(N__32796),
            .I(aluOperand1_2_rep1));
    CascadeMux I__4598 (
            .O(N__32789),
            .I(\ALU.dout_3_ns_1_0_cascade_ ));
    CascadeMux I__4597 (
            .O(N__32786),
            .I(ALU_N_1085_cascade_));
    InMux I__4596 (
            .O(N__32783),
            .I(N__32780));
    LocalMux I__4595 (
            .O(N__32780),
            .I(\CONTROL.operand1_ne_RNIHKCU2_0Z0Z_0 ));
    InMux I__4594 (
            .O(N__32777),
            .I(N__32771));
    InMux I__4593 (
            .O(N__32776),
            .I(N__32771));
    LocalMux I__4592 (
            .O(N__32771),
            .I(ALU_N_1133));
    InMux I__4591 (
            .O(N__32768),
            .I(N__32762));
    InMux I__4590 (
            .O(N__32767),
            .I(N__32762));
    LocalMux I__4589 (
            .O(N__32762),
            .I(ALU_N_1085));
    InMux I__4588 (
            .O(N__32759),
            .I(N__32753));
    InMux I__4587 (
            .O(N__32758),
            .I(N__32753));
    LocalMux I__4586 (
            .O(N__32753),
            .I(N__32750));
    Odrv4 I__4585 (
            .O(N__32750),
            .I(busState_1_RNI9P5V3_2));
    CascadeMux I__4584 (
            .O(N__32747),
            .I(\ALU.dout_3_ns_1_1_cascade_ ));
    CascadeMux I__4583 (
            .O(N__32744),
            .I(ALU_N_1086_cascade_));
    InMux I__4582 (
            .O(N__32741),
            .I(N__32738));
    LocalMux I__4581 (
            .O(N__32738),
            .I(ALU_N_1134));
    CascadeMux I__4580 (
            .O(N__32735),
            .I(\ALU.dout_6_ns_1_6_cascade_ ));
    InMux I__4579 (
            .O(N__32732),
            .I(N__32729));
    LocalMux I__4578 (
            .O(N__32729),
            .I(N__32725));
    CascadeMux I__4577 (
            .O(N__32728),
            .I(N__32722));
    Span4Mux_h I__4576 (
            .O(N__32725),
            .I(N__32719));
    InMux I__4575 (
            .O(N__32722),
            .I(N__32716));
    Sp12to4 I__4574 (
            .O(N__32719),
            .I(N__32713));
    LocalMux I__4573 (
            .O(N__32716),
            .I(\ALU.eZ0Z_6 ));
    Odrv12 I__4572 (
            .O(N__32713),
            .I(\ALU.eZ0Z_6 ));
    CascadeMux I__4571 (
            .O(N__32708),
            .I(\ALU.dout_3_ns_1_6_cascade_ ));
    CascadeMux I__4570 (
            .O(N__32705),
            .I(\ALU.N_1091_cascade_ ));
    InMux I__4569 (
            .O(N__32702),
            .I(N__32699));
    LocalMux I__4568 (
            .O(N__32699),
            .I(\ALU.N_1139 ));
    CascadeMux I__4567 (
            .O(N__32696),
            .I(aluOut_6_cascade_));
    CascadeMux I__4566 (
            .O(N__32693),
            .I(N__32690));
    InMux I__4565 (
            .O(N__32690),
            .I(N__32684));
    InMux I__4564 (
            .O(N__32689),
            .I(N__32684));
    LocalMux I__4563 (
            .O(N__32684),
            .I(N__32681));
    Span4Mux_v I__4562 (
            .O(N__32681),
            .I(N__32678));
    Odrv4 I__4561 (
            .O(N__32678),
            .I(\ALU.d_RNIR3N75Z0Z_6 ));
    CascadeMux I__4560 (
            .O(N__32675),
            .I(\ALU.dout_6_ns_1_1_cascade_ ));
    CascadeMux I__4559 (
            .O(N__32672),
            .I(ALU_N_1134_cascade_));
    InMux I__4558 (
            .O(N__32669),
            .I(N__32666));
    LocalMux I__4557 (
            .O(N__32666),
            .I(\CONTROL.operand1_ne_RNIBQE03Z0Z_0 ));
    CascadeMux I__4556 (
            .O(N__32663),
            .I(N__32659));
    CascadeMux I__4555 (
            .O(N__32662),
            .I(N__32656));
    InMux I__4554 (
            .O(N__32659),
            .I(N__32653));
    InMux I__4553 (
            .O(N__32656),
            .I(N__32650));
    LocalMux I__4552 (
            .O(N__32653),
            .I(N__32645));
    LocalMux I__4551 (
            .O(N__32650),
            .I(N__32645));
    Span4Mux_v I__4550 (
            .O(N__32645),
            .I(N__32642));
    Span4Mux_h I__4549 (
            .O(N__32642),
            .I(N__32639));
    Odrv4 I__4548 (
            .O(N__32639),
            .I(\ALU.eZ0Z_4 ));
    CascadeMux I__4547 (
            .O(N__32636),
            .I(N__32632));
    InMux I__4546 (
            .O(N__32635),
            .I(N__32629));
    InMux I__4545 (
            .O(N__32632),
            .I(N__32626));
    LocalMux I__4544 (
            .O(N__32629),
            .I(N__32623));
    LocalMux I__4543 (
            .O(N__32626),
            .I(N__32620));
    Span4Mux_v I__4542 (
            .O(N__32623),
            .I(N__32617));
    Span4Mux_v I__4541 (
            .O(N__32620),
            .I(N__32614));
    Sp12to4 I__4540 (
            .O(N__32617),
            .I(N__32609));
    Sp12to4 I__4539 (
            .O(N__32614),
            .I(N__32609));
    Odrv12 I__4538 (
            .O(N__32609),
            .I(\ALU.eZ0Z_10 ));
    CascadeMux I__4537 (
            .O(N__32606),
            .I(N__32603));
    InMux I__4536 (
            .O(N__32603),
            .I(N__32600));
    LocalMux I__4535 (
            .O(N__32600),
            .I(N__32596));
    InMux I__4534 (
            .O(N__32599),
            .I(N__32593));
    Span4Mux_v I__4533 (
            .O(N__32596),
            .I(N__32590));
    LocalMux I__4532 (
            .O(N__32593),
            .I(N__32587));
    Span4Mux_h I__4531 (
            .O(N__32590),
            .I(N__32584));
    Span12Mux_v I__4530 (
            .O(N__32587),
            .I(N__32581));
    Span4Mux_v I__4529 (
            .O(N__32584),
            .I(N__32578));
    Odrv12 I__4528 (
            .O(N__32581),
            .I(\ALU.eZ0Z_11 ));
    Odrv4 I__4527 (
            .O(N__32578),
            .I(\ALU.eZ0Z_11 ));
    IoInMux I__4526 (
            .O(N__32573),
            .I(N__32570));
    LocalMux I__4525 (
            .O(N__32570),
            .I(N__32564));
    CascadeMux I__4524 (
            .O(N__32569),
            .I(N__32559));
    CascadeMux I__4523 (
            .O(N__32568),
            .I(N__32555));
    CascadeMux I__4522 (
            .O(N__32567),
            .I(N__32551));
    IoSpan4Mux I__4521 (
            .O(N__32564),
            .I(N__32548));
    SRMux I__4520 (
            .O(N__32563),
            .I(N__32545));
    InMux I__4519 (
            .O(N__32562),
            .I(N__32531));
    InMux I__4518 (
            .O(N__32559),
            .I(N__32531));
    InMux I__4517 (
            .O(N__32558),
            .I(N__32531));
    InMux I__4516 (
            .O(N__32555),
            .I(N__32531));
    InMux I__4515 (
            .O(N__32554),
            .I(N__32531));
    InMux I__4514 (
            .O(N__32551),
            .I(N__32531));
    Span4Mux_s3_v I__4513 (
            .O(N__32548),
            .I(N__32527));
    LocalMux I__4512 (
            .O(N__32545),
            .I(N__32524));
    SRMux I__4511 (
            .O(N__32544),
            .I(N__32521));
    LocalMux I__4510 (
            .O(N__32531),
            .I(N__32518));
    SRMux I__4509 (
            .O(N__32530),
            .I(N__32515));
    Span4Mux_v I__4508 (
            .O(N__32527),
            .I(N__32502));
    Span4Mux_v I__4507 (
            .O(N__32524),
            .I(N__32502));
    LocalMux I__4506 (
            .O(N__32521),
            .I(N__32502));
    Span4Mux_h I__4505 (
            .O(N__32518),
            .I(N__32502));
    LocalMux I__4504 (
            .O(N__32515),
            .I(N__32502));
    SRMux I__4503 (
            .O(N__32514),
            .I(N__32499));
    SRMux I__4502 (
            .O(N__32513),
            .I(N__32496));
    Span4Mux_v I__4501 (
            .O(N__32502),
            .I(N__32486));
    LocalMux I__4500 (
            .O(N__32499),
            .I(N__32486));
    LocalMux I__4499 (
            .O(N__32496),
            .I(N__32486));
    SRMux I__4498 (
            .O(N__32495),
            .I(N__32483));
    IoInMux I__4497 (
            .O(N__32494),
            .I(N__32476));
    IoInMux I__4496 (
            .O(N__32493),
            .I(N__32473));
    Span4Mux_v I__4495 (
            .O(N__32486),
            .I(N__32468));
    LocalMux I__4494 (
            .O(N__32483),
            .I(N__32468));
    CascadeMux I__4493 (
            .O(N__32482),
            .I(N__32465));
    CascadeMux I__4492 (
            .O(N__32481),
            .I(N__32461));
    CascadeMux I__4491 (
            .O(N__32480),
            .I(N__32458));
    CascadeMux I__4490 (
            .O(N__32479),
            .I(N__32453));
    LocalMux I__4489 (
            .O(N__32476),
            .I(N__32448));
    LocalMux I__4488 (
            .O(N__32473),
            .I(N__32448));
    Span4Mux_v I__4487 (
            .O(N__32468),
            .I(N__32445));
    InMux I__4486 (
            .O(N__32465),
            .I(N__32442));
    InMux I__4485 (
            .O(N__32464),
            .I(N__32429));
    InMux I__4484 (
            .O(N__32461),
            .I(N__32429));
    InMux I__4483 (
            .O(N__32458),
            .I(N__32429));
    InMux I__4482 (
            .O(N__32457),
            .I(N__32429));
    InMux I__4481 (
            .O(N__32456),
            .I(N__32429));
    InMux I__4480 (
            .O(N__32453),
            .I(N__32429));
    Span4Mux_s3_h I__4479 (
            .O(N__32448),
            .I(N__32424));
    Span4Mux_v I__4478 (
            .O(N__32445),
            .I(N__32424));
    LocalMux I__4477 (
            .O(N__32442),
            .I(N__32417));
    LocalMux I__4476 (
            .O(N__32429),
            .I(N__32417));
    Sp12to4 I__4475 (
            .O(N__32424),
            .I(N__32417));
    Span12Mux_h I__4474 (
            .O(N__32417),
            .I(N__32414));
    Odrv12 I__4473 (
            .O(N__32414),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4472 (
            .O(N__32411),
            .I(N__32408));
    InMux I__4471 (
            .O(N__32408),
            .I(N__32405));
    LocalMux I__4470 (
            .O(N__32405),
            .I(\ALU.d_RNI290AE1Z0Z_0 ));
    InMux I__4469 (
            .O(N__32402),
            .I(N__32399));
    LocalMux I__4468 (
            .O(N__32399),
            .I(\ALU.d_RNI5MTIOZ0Z_1 ));
    CascadeMux I__4467 (
            .O(N__32396),
            .I(busState_1_RNICT0U1_2_cascade_));
    CascadeMux I__4466 (
            .O(N__32393),
            .I(N__32389));
    InMux I__4465 (
            .O(N__32392),
            .I(N__32384));
    InMux I__4464 (
            .O(N__32389),
            .I(N__32384));
    LocalMux I__4463 (
            .O(N__32384),
            .I(busState_1_RNICT0U1_2));
    CascadeMux I__4462 (
            .O(N__32381),
            .I(N_227_0_cascade_));
    CascadeMux I__4461 (
            .O(N__32378),
            .I(N__32375));
    InMux I__4460 (
            .O(N__32375),
            .I(N__32372));
    LocalMux I__4459 (
            .O(N__32372),
            .I(N__32369));
    Span4Mux_h I__4458 (
            .O(N__32369),
            .I(N__32366));
    Span4Mux_h I__4457 (
            .O(N__32366),
            .I(N__32363));
    Span4Mux_h I__4456 (
            .O(N__32363),
            .I(N__32360));
    Odrv4 I__4455 (
            .O(N__32360),
            .I(\ALU.status_18_cry_2_c_RNOZ0 ));
    CascadeMux I__4454 (
            .O(N__32357),
            .I(N__32354));
    InMux I__4453 (
            .O(N__32354),
            .I(N__32351));
    LocalMux I__4452 (
            .O(N__32351),
            .I(DROM_ROMDATA_dintern_2ro));
    InMux I__4451 (
            .O(N__32348),
            .I(N__32342));
    InMux I__4450 (
            .O(N__32347),
            .I(N__32342));
    LocalMux I__4449 (
            .O(N__32342),
            .I(N__32339));
    Span4Mux_h I__4448 (
            .O(N__32339),
            .I(N__32336));
    Span4Mux_v I__4447 (
            .O(N__32336),
            .I(N__32333));
    Odrv4 I__4446 (
            .O(N__32333),
            .I(\DROM.ROMDATA.dintern_0_0_NEW_2 ));
    InMux I__4445 (
            .O(N__32330),
            .I(N__32327));
    LocalMux I__4444 (
            .O(N__32327),
            .I(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_2 ));
    CEMux I__4443 (
            .O(N__32324),
            .I(N__32315));
    CEMux I__4442 (
            .O(N__32323),
            .I(N__32312));
    InMux I__4441 (
            .O(N__32322),
            .I(N__32309));
    CEMux I__4440 (
            .O(N__32321),
            .I(N__32304));
    CEMux I__4439 (
            .O(N__32320),
            .I(N__32296));
    CEMux I__4438 (
            .O(N__32319),
            .I(N__32290));
    InMux I__4437 (
            .O(N__32318),
            .I(N__32290));
    LocalMux I__4436 (
            .O(N__32315),
            .I(N__32287));
    LocalMux I__4435 (
            .O(N__32312),
            .I(N__32282));
    LocalMux I__4434 (
            .O(N__32309),
            .I(N__32282));
    InMux I__4433 (
            .O(N__32308),
            .I(N__32277));
    InMux I__4432 (
            .O(N__32307),
            .I(N__32277));
    LocalMux I__4431 (
            .O(N__32304),
            .I(N__32274));
    InMux I__4430 (
            .O(N__32303),
            .I(N__32265));
    InMux I__4429 (
            .O(N__32302),
            .I(N__32265));
    InMux I__4428 (
            .O(N__32301),
            .I(N__32265));
    InMux I__4427 (
            .O(N__32300),
            .I(N__32265));
    CEMux I__4426 (
            .O(N__32299),
            .I(N__32257));
    LocalMux I__4425 (
            .O(N__32296),
            .I(N__32254));
    InMux I__4424 (
            .O(N__32295),
            .I(N__32251));
    LocalMux I__4423 (
            .O(N__32290),
            .I(N__32248));
    Span4Mux_h I__4422 (
            .O(N__32287),
            .I(N__32243));
    Span4Mux_h I__4421 (
            .O(N__32282),
            .I(N__32240));
    LocalMux I__4420 (
            .O(N__32277),
            .I(N__32237));
    Span4Mux_v I__4419 (
            .O(N__32274),
            .I(N__32232));
    LocalMux I__4418 (
            .O(N__32265),
            .I(N__32232));
    InMux I__4417 (
            .O(N__32264),
            .I(N__32221));
    InMux I__4416 (
            .O(N__32263),
            .I(N__32221));
    InMux I__4415 (
            .O(N__32262),
            .I(N__32221));
    InMux I__4414 (
            .O(N__32261),
            .I(N__32221));
    InMux I__4413 (
            .O(N__32260),
            .I(N__32221));
    LocalMux I__4412 (
            .O(N__32257),
            .I(N__32212));
    Span4Mux_v I__4411 (
            .O(N__32254),
            .I(N__32212));
    LocalMux I__4410 (
            .O(N__32251),
            .I(N__32212));
    Span4Mux_h I__4409 (
            .O(N__32248),
            .I(N__32212));
    InMux I__4408 (
            .O(N__32247),
            .I(N__32207));
    InMux I__4407 (
            .O(N__32246),
            .I(N__32207));
    Span4Mux_v I__4406 (
            .O(N__32243),
            .I(N__32200));
    Span4Mux_v I__4405 (
            .O(N__32240),
            .I(N__32200));
    Span4Mux_h I__4404 (
            .O(N__32237),
            .I(N__32200));
    Odrv4 I__4403 (
            .O(N__32232),
            .I(\DROM.ROMDATA.dintern_0_0_sr_enZ0 ));
    LocalMux I__4402 (
            .O(N__32221),
            .I(\DROM.ROMDATA.dintern_0_0_sr_enZ0 ));
    Odrv4 I__4401 (
            .O(N__32212),
            .I(\DROM.ROMDATA.dintern_0_0_sr_enZ0 ));
    LocalMux I__4400 (
            .O(N__32207),
            .I(\DROM.ROMDATA.dintern_0_0_sr_enZ0 ));
    Odrv4 I__4399 (
            .O(N__32200),
            .I(\DROM.ROMDATA.dintern_0_0_sr_enZ0 ));
    InMux I__4398 (
            .O(N__32189),
            .I(N__32186));
    LocalMux I__4397 (
            .O(N__32186),
            .I(\ALU.mult_1_12 ));
    CascadeMux I__4396 (
            .O(N__32183),
            .I(N__32180));
    InMux I__4395 (
            .O(N__32180),
            .I(N__32177));
    LocalMux I__4394 (
            .O(N__32177),
            .I(N__32174));
    Span4Mux_v I__4393 (
            .O(N__32174),
            .I(N__32171));
    Odrv4 I__4392 (
            .O(N__32171),
            .I(\ALU.mult_3_12 ));
    InMux I__4391 (
            .O(N__32168),
            .I(\ALU.mult_17_c11 ));
    InMux I__4390 (
            .O(N__32165),
            .I(N__32162));
    LocalMux I__4389 (
            .O(N__32162),
            .I(\ALU.mult_1_13 ));
    CascadeMux I__4388 (
            .O(N__32159),
            .I(N__32156));
    InMux I__4387 (
            .O(N__32156),
            .I(N__32153));
    LocalMux I__4386 (
            .O(N__32153),
            .I(N__32150));
    Span4Mux_h I__4385 (
            .O(N__32150),
            .I(N__32147));
    Odrv4 I__4384 (
            .O(N__32147),
            .I(\ALU.mult_3_13 ));
    InMux I__4383 (
            .O(N__32144),
            .I(\ALU.mult_17_c12 ));
    InMux I__4382 (
            .O(N__32141),
            .I(N__32138));
    LocalMux I__4381 (
            .O(N__32138),
            .I(\ALU.mult_1_14 ));
    CascadeMux I__4380 (
            .O(N__32135),
            .I(N__32132));
    InMux I__4379 (
            .O(N__32132),
            .I(N__32129));
    LocalMux I__4378 (
            .O(N__32129),
            .I(N__32126));
    Span4Mux_h I__4377 (
            .O(N__32126),
            .I(N__32123));
    Odrv4 I__4376 (
            .O(N__32123),
            .I(\ALU.mult_3_14 ));
    InMux I__4375 (
            .O(N__32120),
            .I(\ALU.mult_17_c13 ));
    InMux I__4374 (
            .O(N__32117),
            .I(N__32114));
    LocalMux I__4373 (
            .O(N__32114),
            .I(N__32111));
    Odrv4 I__4372 (
            .O(N__32111),
            .I(\ALU.mult_227_c_RNIBPRVZ0Z92 ));
    InMux I__4371 (
            .O(N__32108),
            .I(N__32105));
    LocalMux I__4370 (
            .O(N__32105),
            .I(\ALU.mult_83_c_RNIKEU6BZ0Z2 ));
    InMux I__4369 (
            .O(N__32102),
            .I(\ALU.mult_17_c14 ));
    InMux I__4368 (
            .O(N__32099),
            .I(N__32096));
    LocalMux I__4367 (
            .O(N__32096),
            .I(\ALU.d_RNIHU6RLZ0Z_1 ));
    CascadeMux I__4366 (
            .O(N__32093),
            .I(N__32090));
    InMux I__4365 (
            .O(N__32090),
            .I(N__32087));
    LocalMux I__4364 (
            .O(N__32087),
            .I(N__32084));
    Span4Mux_h I__4363 (
            .O(N__32084),
            .I(N__32081));
    Odrv4 I__4362 (
            .O(N__32081),
            .I(\ALU.d_RNI2E4JE1Z0Z_4 ));
    InMux I__4361 (
            .O(N__32078),
            .I(N__32075));
    LocalMux I__4360 (
            .O(N__32075),
            .I(N__32072));
    Span4Mux_h I__4359 (
            .O(N__32072),
            .I(N__32069));
    Span4Mux_v I__4358 (
            .O(N__32069),
            .I(N__32066));
    Odrv4 I__4357 (
            .O(N__32066),
            .I(\ALU.N_860 ));
    InMux I__4356 (
            .O(N__32063),
            .I(N__32060));
    LocalMux I__4355 (
            .O(N__32060),
            .I(\ALU.mult_5_c_RNOZ0 ));
    InMux I__4354 (
            .O(N__32057),
            .I(N__32054));
    LocalMux I__4353 (
            .O(N__32054),
            .I(N__32051));
    Span4Mux_v I__4352 (
            .O(N__32051),
            .I(N__32048));
    Odrv4 I__4351 (
            .O(N__32048),
            .I(\ALU.mult_3_4 ));
    CascadeMux I__4350 (
            .O(N__32045),
            .I(N__32042));
    InMux I__4349 (
            .O(N__32042),
            .I(N__32039));
    LocalMux I__4348 (
            .O(N__32039),
            .I(\ALU.mult_1_4 ));
    InMux I__4347 (
            .O(N__32036),
            .I(\ALU.mult_17_c3 ));
    InMux I__4346 (
            .O(N__32033),
            .I(N__32030));
    LocalMux I__4345 (
            .O(N__32030),
            .I(\ALU.mult_1_5 ));
    CascadeMux I__4344 (
            .O(N__32027),
            .I(N__32024));
    InMux I__4343 (
            .O(N__32024),
            .I(N__32021));
    LocalMux I__4342 (
            .O(N__32021),
            .I(N__32018));
    Span4Mux_h I__4341 (
            .O(N__32018),
            .I(N__32015));
    Odrv4 I__4340 (
            .O(N__32015),
            .I(\ALU.mult_3_5 ));
    InMux I__4339 (
            .O(N__32012),
            .I(\ALU.mult_17_c4 ));
    InMux I__4338 (
            .O(N__32009),
            .I(N__32006));
    LocalMux I__4337 (
            .O(N__32006),
            .I(N__32003));
    Odrv4 I__4336 (
            .O(N__32003),
            .I(\ALU.mult_1_6 ));
    CascadeMux I__4335 (
            .O(N__32000),
            .I(N__31997));
    InMux I__4334 (
            .O(N__31997),
            .I(N__31994));
    LocalMux I__4333 (
            .O(N__31994),
            .I(N__31991));
    Span4Mux_h I__4332 (
            .O(N__31991),
            .I(N__31988));
    Odrv4 I__4331 (
            .O(N__31988),
            .I(\ALU.mult_3_6 ));
    InMux I__4330 (
            .O(N__31985),
            .I(\ALU.mult_17_c5 ));
    InMux I__4329 (
            .O(N__31982),
            .I(N__31979));
    LocalMux I__4328 (
            .O(N__31979),
            .I(\ALU.mult_1_7 ));
    CascadeMux I__4327 (
            .O(N__31976),
            .I(N__31973));
    InMux I__4326 (
            .O(N__31973),
            .I(N__31970));
    LocalMux I__4325 (
            .O(N__31970),
            .I(N__31967));
    Span4Mux_h I__4324 (
            .O(N__31967),
            .I(N__31964));
    Odrv4 I__4323 (
            .O(N__31964),
            .I(\ALU.mult_3_7 ));
    InMux I__4322 (
            .O(N__31961),
            .I(\ALU.mult_17_c6 ));
    InMux I__4321 (
            .O(N__31958),
            .I(N__31955));
    LocalMux I__4320 (
            .O(N__31955),
            .I(\ALU.mult_1_8 ));
    CascadeMux I__4319 (
            .O(N__31952),
            .I(N__31949));
    InMux I__4318 (
            .O(N__31949),
            .I(N__31946));
    LocalMux I__4317 (
            .O(N__31946),
            .I(N__31943));
    Span4Mux_h I__4316 (
            .O(N__31943),
            .I(N__31940));
    Odrv4 I__4315 (
            .O(N__31940),
            .I(\ALU.mult_3_8 ));
    InMux I__4314 (
            .O(N__31937),
            .I(\ALU.mult_17_c7 ));
    InMux I__4313 (
            .O(N__31934),
            .I(N__31931));
    LocalMux I__4312 (
            .O(N__31931),
            .I(N__31928));
    Odrv4 I__4311 (
            .O(N__31928),
            .I(\ALU.mult_1_9 ));
    CascadeMux I__4310 (
            .O(N__31925),
            .I(N__31922));
    InMux I__4309 (
            .O(N__31922),
            .I(N__31919));
    LocalMux I__4308 (
            .O(N__31919),
            .I(N__31916));
    Span4Mux_h I__4307 (
            .O(N__31916),
            .I(N__31913));
    Odrv4 I__4306 (
            .O(N__31913),
            .I(\ALU.mult_3_9 ));
    InMux I__4305 (
            .O(N__31910),
            .I(\ALU.mult_17_c8 ));
    InMux I__4304 (
            .O(N__31907),
            .I(N__31904));
    LocalMux I__4303 (
            .O(N__31904),
            .I(N__31901));
    Odrv12 I__4302 (
            .O(N__31901),
            .I(\ALU.mult_3_10 ));
    CascadeMux I__4301 (
            .O(N__31898),
            .I(N__31895));
    InMux I__4300 (
            .O(N__31895),
            .I(N__31892));
    LocalMux I__4299 (
            .O(N__31892),
            .I(\ALU.mult_1_10 ));
    InMux I__4298 (
            .O(N__31889),
            .I(bfn_14_11_0_));
    InMux I__4297 (
            .O(N__31886),
            .I(N__31883));
    LocalMux I__4296 (
            .O(N__31883),
            .I(\ALU.mult_1_11 ));
    CascadeMux I__4295 (
            .O(N__31880),
            .I(N__31877));
    InMux I__4294 (
            .O(N__31877),
            .I(N__31874));
    LocalMux I__4293 (
            .O(N__31874),
            .I(N__31871));
    Span4Mux_v I__4292 (
            .O(N__31871),
            .I(N__31868));
    Odrv4 I__4291 (
            .O(N__31868),
            .I(\ALU.mult_3_11 ));
    InMux I__4290 (
            .O(N__31865),
            .I(\ALU.mult_17_c10 ));
    InMux I__4289 (
            .O(N__31862),
            .I(N__31859));
    LocalMux I__4288 (
            .O(N__31859),
            .I(N__31856));
    Span4Mux_h I__4287 (
            .O(N__31856),
            .I(N__31853));
    Odrv4 I__4286 (
            .O(N__31853),
            .I(\ALU.d_RNIB5POHZ0Z_5 ));
    CascadeMux I__4285 (
            .O(N__31850),
            .I(N__31847));
    InMux I__4284 (
            .O(N__31847),
            .I(N__31844));
    LocalMux I__4283 (
            .O(N__31844),
            .I(N__31841));
    Odrv12 I__4282 (
            .O(N__31841),
            .I(\ALU.d_RNIPNF141Z0Z_4 ));
    InMux I__4281 (
            .O(N__31838),
            .I(bfn_14_9_0_));
    InMux I__4280 (
            .O(N__31835),
            .I(N__31832));
    LocalMux I__4279 (
            .O(N__31832),
            .I(N__31829));
    Odrv12 I__4278 (
            .O(N__31829),
            .I(\ALU.d_RNI88K161Z0Z_4 ));
    CascadeMux I__4277 (
            .O(N__31826),
            .I(N__31823));
    InMux I__4276 (
            .O(N__31823),
            .I(N__31820));
    LocalMux I__4275 (
            .O(N__31820),
            .I(N__31817));
    Span4Mux_v I__4274 (
            .O(N__31817),
            .I(N__31814));
    Odrv4 I__4273 (
            .O(N__31814),
            .I(\ALU.d_RNIMQM8IZ0Z_5 ));
    InMux I__4272 (
            .O(N__31811),
            .I(\ALU.mult_5_c13 ));
    InMux I__4271 (
            .O(N__31808),
            .I(N__31805));
    LocalMux I__4270 (
            .O(N__31805),
            .I(\ALU.mult_7_c14_THRU_CO ));
    InMux I__4269 (
            .O(N__31802),
            .I(N__31799));
    LocalMux I__4268 (
            .O(N__31799),
            .I(N__31796));
    Span4Mux_h I__4267 (
            .O(N__31796),
            .I(N__31793));
    Span4Mux_v I__4266 (
            .O(N__31793),
            .I(N__31790));
    Odrv4 I__4265 (
            .O(N__31790),
            .I(\ALU.d_RNIKDVI51Z0Z_4 ));
    CascadeMux I__4264 (
            .O(N__31787),
            .I(N__31784));
    InMux I__4263 (
            .O(N__31784),
            .I(N__31781));
    LocalMux I__4262 (
            .O(N__31781),
            .I(N__31778));
    Span4Mux_v I__4261 (
            .O(N__31778),
            .I(N__31775));
    Span4Mux_h I__4260 (
            .O(N__31775),
            .I(N__31772));
    Odrv4 I__4259 (
            .O(N__31772),
            .I(\ALU.d_RNIRU9M31Z0Z_6 ));
    InMux I__4258 (
            .O(N__31769),
            .I(\ALU.mult_5_c14 ));
    InMux I__4257 (
            .O(N__31766),
            .I(N__31763));
    LocalMux I__4256 (
            .O(N__31763),
            .I(N__31760));
    Span4Mux_h I__4255 (
            .O(N__31760),
            .I(N__31757));
    Span4Mux_h I__4254 (
            .O(N__31757),
            .I(N__31752));
    InMux I__4253 (
            .O(N__31756),
            .I(N__31747));
    InMux I__4252 (
            .O(N__31755),
            .I(N__31747));
    Sp12to4 I__4251 (
            .O(N__31752),
            .I(N__31744));
    LocalMux I__4250 (
            .O(N__31747),
            .I(N__31741));
    Span12Mux_v I__4249 (
            .O(N__31744),
            .I(N__31738));
    Span4Mux_v I__4248 (
            .O(N__31741),
            .I(N__31735));
    Odrv12 I__4247 (
            .O(N__31738),
            .I(bus_0_12));
    Odrv4 I__4246 (
            .O(N__31735),
            .I(bus_0_12));
    CascadeMux I__4245 (
            .O(N__31730),
            .I(N__31727));
    InMux I__4244 (
            .O(N__31727),
            .I(N__31724));
    LocalMux I__4243 (
            .O(N__31724),
            .I(\ALU.mult_239_c_RNOZ0Z_0 ));
    InMux I__4242 (
            .O(N__31721),
            .I(N__31718));
    LocalMux I__4241 (
            .O(N__31718),
            .I(\ALU.mult_239_c_RNOZ0 ));
    CascadeMux I__4240 (
            .O(N__31715),
            .I(N__31711));
    InMux I__4239 (
            .O(N__31714),
            .I(N__31706));
    InMux I__4238 (
            .O(N__31711),
            .I(N__31706));
    LocalMux I__4237 (
            .O(N__31706),
            .I(N__31703));
    Odrv4 I__4236 (
            .O(N__31703),
            .I(\ALU.mult_1_2 ));
    CascadeMux I__4235 (
            .O(N__31700),
            .I(N__31697));
    InMux I__4234 (
            .O(N__31697),
            .I(N__31694));
    LocalMux I__4233 (
            .O(N__31694),
            .I(\ALU.mult_1_3 ));
    InMux I__4232 (
            .O(N__31691),
            .I(\ALU.mult_17_c2 ));
    CascadeMux I__4231 (
            .O(N__31688),
            .I(N__31685));
    InMux I__4230 (
            .O(N__31685),
            .I(N__31682));
    LocalMux I__4229 (
            .O(N__31682),
            .I(\ALU.mult_173_c_RNOZ0Z_0 ));
    InMux I__4228 (
            .O(N__31679),
            .I(\ALU.mult_5_c5 ));
    InMux I__4227 (
            .O(N__31676),
            .I(N__31673));
    LocalMux I__4226 (
            .O(N__31673),
            .I(N__31670));
    Odrv4 I__4225 (
            .O(N__31670),
            .I(\ALU.d_RNIFGNR61Z0Z_4 ));
    InMux I__4224 (
            .O(N__31667),
            .I(\ALU.mult_5_c6 ));
    InMux I__4223 (
            .O(N__31664),
            .I(N__31661));
    LocalMux I__4222 (
            .O(N__31661),
            .I(\ALU.d_RNICP0UGZ0Z_5 ));
    CascadeMux I__4221 (
            .O(N__31658),
            .I(N__31655));
    InMux I__4220 (
            .O(N__31655),
            .I(N__31652));
    LocalMux I__4219 (
            .O(N__31652),
            .I(\ALU.d_RNI6CL331Z0Z_4 ));
    InMux I__4218 (
            .O(N__31649),
            .I(\ALU.mult_5_c7 ));
    InMux I__4217 (
            .O(N__31646),
            .I(N__31643));
    LocalMux I__4216 (
            .O(N__31643),
            .I(N__31640));
    Span4Mux_h I__4215 (
            .O(N__31640),
            .I(N__31637));
    Odrv4 I__4214 (
            .O(N__31637),
            .I(\ALU.d_RNI2RK5IZ0Z_5 ));
    InMux I__4213 (
            .O(N__31634),
            .I(\ALU.mult_5_c8 ));
    InMux I__4212 (
            .O(N__31631),
            .I(N__31628));
    LocalMux I__4211 (
            .O(N__31628),
            .I(N__31625));
    Span4Mux_h I__4210 (
            .O(N__31625),
            .I(N__31622));
    Odrv4 I__4209 (
            .O(N__31622),
            .I(\ALU.d_RNIOFVDIZ0Z_5 ));
    CascadeMux I__4208 (
            .O(N__31619),
            .I(N__31616));
    InMux I__4207 (
            .O(N__31616),
            .I(N__31613));
    LocalMux I__4206 (
            .O(N__31613),
            .I(N__31610));
    Odrv4 I__4205 (
            .O(N__31610),
            .I(\ALU.d_RNI5SIF41Z0Z_4 ));
    InMux I__4204 (
            .O(N__31607),
            .I(\ALU.mult_5_c9 ));
    InMux I__4203 (
            .O(N__31604),
            .I(N__31601));
    LocalMux I__4202 (
            .O(N__31601),
            .I(N__31598));
    Span4Mux_h I__4201 (
            .O(N__31598),
            .I(N__31595));
    Span4Mux_h I__4200 (
            .O(N__31595),
            .I(N__31592));
    Odrv4 I__4199 (
            .O(N__31592),
            .I(\ALU.d_RNILKJ1IZ0Z_5 ));
    CascadeMux I__4198 (
            .O(N__31589),
            .I(N__31586));
    InMux I__4197 (
            .O(N__31586),
            .I(N__31583));
    LocalMux I__4196 (
            .O(N__31583),
            .I(N__31580));
    Span4Mux_h I__4195 (
            .O(N__31580),
            .I(N__31577));
    Odrv4 I__4194 (
            .O(N__31577),
            .I(\ALU.d_RNIJTUN21Z0Z_4 ));
    InMux I__4193 (
            .O(N__31574),
            .I(\ALU.mult_5_c10 ));
    InMux I__4192 (
            .O(N__31571),
            .I(N__31568));
    LocalMux I__4191 (
            .O(N__31568),
            .I(N__31565));
    Span4Mux_v I__4190 (
            .O(N__31565),
            .I(N__31562));
    Odrv4 I__4189 (
            .O(N__31562),
            .I(\ALU.d_RNI6HBMGZ0Z_5 ));
    CascadeMux I__4188 (
            .O(N__31559),
            .I(N__31556));
    InMux I__4187 (
            .O(N__31556),
            .I(N__31553));
    LocalMux I__4186 (
            .O(N__31553),
            .I(N__31550));
    Span4Mux_h I__4185 (
            .O(N__31550),
            .I(N__31547));
    Odrv4 I__4184 (
            .O(N__31547),
            .I(\ALU.d_RNI9E4F21Z0Z_4 ));
    InMux I__4183 (
            .O(N__31544),
            .I(\ALU.mult_5_c11 ));
    InMux I__4182 (
            .O(N__31541),
            .I(N__31538));
    LocalMux I__4181 (
            .O(N__31538),
            .I(\CONTROL.g1_0 ));
    InMux I__4180 (
            .O(N__31535),
            .I(N__31532));
    LocalMux I__4179 (
            .O(N__31532),
            .I(N__31528));
    CascadeMux I__4178 (
            .O(N__31531),
            .I(N__31525));
    Span4Mux_v I__4177 (
            .O(N__31528),
            .I(N__31521));
    InMux I__4176 (
            .O(N__31525),
            .I(N__31518));
    CascadeMux I__4175 (
            .O(N__31524),
            .I(N__31515));
    Span4Mux_h I__4174 (
            .O(N__31521),
            .I(N__31512));
    LocalMux I__4173 (
            .O(N__31518),
            .I(N__31509));
    InMux I__4172 (
            .O(N__31515),
            .I(N__31506));
    Odrv4 I__4171 (
            .O(N__31512),
            .I(\CONTROL.addrstack_1_1 ));
    Odrv4 I__4170 (
            .O(N__31509),
            .I(\CONTROL.addrstack_1_1 ));
    LocalMux I__4169 (
            .O(N__31506),
            .I(\CONTROL.addrstack_1_1 ));
    CascadeMux I__4168 (
            .O(N__31499),
            .I(\CONTROL.g1_0_cascade_ ));
    CascadeMux I__4167 (
            .O(N__31496),
            .I(\CONTROL.g0_1_i_a6Z0Z_4_cascade_ ));
    InMux I__4166 (
            .O(N__31493),
            .I(N__31489));
    InMux I__4165 (
            .O(N__31492),
            .I(N__31486));
    LocalMux I__4164 (
            .O(N__31489),
            .I(\CONTROL.N_9 ));
    LocalMux I__4163 (
            .O(N__31486),
            .I(\CONTROL.N_9 ));
    CascadeMux I__4162 (
            .O(N__31481),
            .I(N__31478));
    InMux I__4161 (
            .O(N__31478),
            .I(N__31475));
    LocalMux I__4160 (
            .O(N__31475),
            .I(N__31472));
    Span4Mux_h I__4159 (
            .O(N__31472),
            .I(N__31469));
    Odrv4 I__4158 (
            .O(N__31469),
            .I(\CONTROL.g0_0_1 ));
    InMux I__4157 (
            .O(N__31466),
            .I(N__31463));
    LocalMux I__4156 (
            .O(N__31463),
            .I(N__31459));
    InMux I__4155 (
            .O(N__31462),
            .I(N__31456));
    Span4Mux_h I__4154 (
            .O(N__31459),
            .I(N__31451));
    LocalMux I__4153 (
            .O(N__31456),
            .I(N__31451));
    Span4Mux_v I__4152 (
            .O(N__31451),
            .I(N__31448));
    Odrv4 I__4151 (
            .O(N__31448),
            .I(\CONTROL.N_366 ));
    InMux I__4150 (
            .O(N__31445),
            .I(N__31441));
    InMux I__4149 (
            .O(N__31444),
            .I(N__31438));
    LocalMux I__4148 (
            .O(N__31441),
            .I(\CONTROL.g0_1_i_3 ));
    LocalMux I__4147 (
            .O(N__31438),
            .I(\CONTROL.g0_1_i_3 ));
    InMux I__4146 (
            .O(N__31433),
            .I(N__31430));
    LocalMux I__4145 (
            .O(N__31430),
            .I(N__31427));
    Odrv12 I__4144 (
            .O(N__31427),
            .I(\CONTROL.addrstack_15 ));
    CascadeMux I__4143 (
            .O(N__31424),
            .I(N__31421));
    InMux I__4142 (
            .O(N__31421),
            .I(N__31418));
    LocalMux I__4141 (
            .O(N__31418),
            .I(N__31415));
    Odrv4 I__4140 (
            .O(N__31415),
            .I(\CONTROL.addrstack_reto_15 ));
    CascadeMux I__4139 (
            .O(N__31412),
            .I(N__31408));
    InMux I__4138 (
            .O(N__31411),
            .I(N__31405));
    InMux I__4137 (
            .O(N__31408),
            .I(N__31401));
    LocalMux I__4136 (
            .O(N__31405),
            .I(N__31398));
    InMux I__4135 (
            .O(N__31404),
            .I(N__31395));
    LocalMux I__4134 (
            .O(N__31401),
            .I(N__31390));
    Span4Mux_h I__4133 (
            .O(N__31398),
            .I(N__31390));
    LocalMux I__4132 (
            .O(N__31395),
            .I(N__31387));
    Span4Mux_h I__4131 (
            .O(N__31390),
            .I(N__31384));
    Span12Mux_v I__4130 (
            .O(N__31387),
            .I(N__31381));
    Odrv4 I__4129 (
            .O(N__31384),
            .I(controlWord_30));
    Odrv12 I__4128 (
            .O(N__31381),
            .I(controlWord_30));
    InMux I__4127 (
            .O(N__31376),
            .I(N__31373));
    LocalMux I__4126 (
            .O(N__31373),
            .I(N__31370));
    Odrv12 I__4125 (
            .O(N__31370),
            .I(\PROM.ROMDATA.m471_ns ));
    InMux I__4124 (
            .O(N__31367),
            .I(N__31364));
    LocalMux I__4123 (
            .O(N__31364),
            .I(N__31361));
    Span4Mux_v I__4122 (
            .O(N__31361),
            .I(N__31358));
    Span4Mux_v I__4121 (
            .O(N__31358),
            .I(N__31355));
    Sp12to4 I__4120 (
            .O(N__31355),
            .I(N__31352));
    Span12Mux_h I__4119 (
            .O(N__31352),
            .I(N__31349));
    Odrv12 I__4118 (
            .O(N__31349),
            .I(gpuOut_c_8));
    InMux I__4117 (
            .O(N__31346),
            .I(N__31342));
    InMux I__4116 (
            .O(N__31345),
            .I(N__31339));
    LocalMux I__4115 (
            .O(N__31342),
            .I(\CONTROL.ctrlOut_8 ));
    LocalMux I__4114 (
            .O(N__31339),
            .I(\CONTROL.ctrlOut_8 ));
    IoInMux I__4113 (
            .O(N__31334),
            .I(N__31331));
    LocalMux I__4112 (
            .O(N__31331),
            .I(N__31328));
    IoSpan4Mux I__4111 (
            .O(N__31328),
            .I(N__31325));
    Sp12to4 I__4110 (
            .O(N__31325),
            .I(N__31322));
    Span12Mux_s7_h I__4109 (
            .O(N__31322),
            .I(N__31319));
    Span12Mux_v I__4108 (
            .O(N__31319),
            .I(N__31316));
    Span12Mux_h I__4107 (
            .O(N__31316),
            .I(N__31313));
    Odrv12 I__4106 (
            .O(N__31313),
            .I(A0_c));
    IoInMux I__4105 (
            .O(N__31310),
            .I(N__31307));
    LocalMux I__4104 (
            .O(N__31307),
            .I(N__31304));
    IoSpan4Mux I__4103 (
            .O(N__31304),
            .I(N__31301));
    Span4Mux_s2_h I__4102 (
            .O(N__31301),
            .I(N__31298));
    Span4Mux_h I__4101 (
            .O(N__31298),
            .I(N__31295));
    Sp12to4 I__4100 (
            .O(N__31295),
            .I(N__31291));
    InMux I__4099 (
            .O(N__31294),
            .I(N__31288));
    Span12Mux_h I__4098 (
            .O(N__31291),
            .I(N__31285));
    LocalMux I__4097 (
            .O(N__31288),
            .I(N__31282));
    Odrv12 I__4096 (
            .O(N__31285),
            .I(A1_c));
    Odrv4 I__4095 (
            .O(N__31282),
            .I(A1_c));
    InMux I__4094 (
            .O(N__31277),
            .I(N__31272));
    InMux I__4093 (
            .O(N__31276),
            .I(N__31269));
    InMux I__4092 (
            .O(N__31275),
            .I(N__31266));
    LocalMux I__4091 (
            .O(N__31272),
            .I(N__31263));
    LocalMux I__4090 (
            .O(N__31269),
            .I(N__31260));
    LocalMux I__4089 (
            .O(N__31266),
            .I(N__31257));
    Span4Mux_h I__4088 (
            .O(N__31263),
            .I(N__31254));
    Span4Mux_h I__4087 (
            .O(N__31260),
            .I(N__31251));
    Span4Mux_v I__4086 (
            .O(N__31257),
            .I(N__31246));
    Span4Mux_h I__4085 (
            .O(N__31254),
            .I(N__31246));
    Span4Mux_h I__4084 (
            .O(N__31251),
            .I(N__31243));
    Odrv4 I__4083 (
            .O(N__31246),
            .I(controlWord_26));
    Odrv4 I__4082 (
            .O(N__31243),
            .I(controlWord_26));
    CascadeMux I__4081 (
            .O(N__31238),
            .I(N__31235));
    InMux I__4080 (
            .O(N__31235),
            .I(N__31230));
    InMux I__4079 (
            .O(N__31234),
            .I(N__31227));
    CascadeMux I__4078 (
            .O(N__31233),
            .I(N__31224));
    LocalMux I__4077 (
            .O(N__31230),
            .I(N__31221));
    LocalMux I__4076 (
            .O(N__31227),
            .I(N__31218));
    InMux I__4075 (
            .O(N__31224),
            .I(N__31215));
    Span4Mux_v I__4074 (
            .O(N__31221),
            .I(N__31212));
    Span12Mux_v I__4073 (
            .O(N__31218),
            .I(N__31207));
    LocalMux I__4072 (
            .O(N__31215),
            .I(N__31207));
    Odrv4 I__4071 (
            .O(N__31212),
            .I(controlWord_27));
    Odrv12 I__4070 (
            .O(N__31207),
            .I(controlWord_27));
    IoInMux I__4069 (
            .O(N__31202),
            .I(N__31199));
    LocalMux I__4068 (
            .O(N__31199),
            .I(N__31196));
    Span12Mux_s9_v I__4067 (
            .O(N__31196),
            .I(N__31193));
    Span12Mux_h I__4066 (
            .O(N__31193),
            .I(N__31189));
    InMux I__4065 (
            .O(N__31192),
            .I(N__31186));
    Odrv12 I__4064 (
            .O(N__31189),
            .I(A10_c));
    LocalMux I__4063 (
            .O(N__31186),
            .I(A10_c));
    IoInMux I__4062 (
            .O(N__31181),
            .I(N__31178));
    LocalMux I__4061 (
            .O(N__31178),
            .I(N__31175));
    IoSpan4Mux I__4060 (
            .O(N__31175),
            .I(N__31172));
    Sp12to4 I__4059 (
            .O(N__31172),
            .I(N__31169));
    Span12Mux_s7_h I__4058 (
            .O(N__31169),
            .I(N__31165));
    CascadeMux I__4057 (
            .O(N__31168),
            .I(N__31162));
    Span12Mux_h I__4056 (
            .O(N__31165),
            .I(N__31159));
    InMux I__4055 (
            .O(N__31162),
            .I(N__31156));
    Odrv12 I__4054 (
            .O(N__31159),
            .I(A11_c));
    LocalMux I__4053 (
            .O(N__31156),
            .I(A11_c));
    InMux I__4052 (
            .O(N__31151),
            .I(N__31148));
    LocalMux I__4051 (
            .O(N__31148),
            .I(N__31145));
    Span4Mux_h I__4050 (
            .O(N__31145),
            .I(N__31142));
    Sp12to4 I__4049 (
            .O(N__31142),
            .I(N__31139));
    Odrv12 I__4048 (
            .O(N__31139),
            .I(\RAM.un1_WR_105_0Z0Z_9 ));
    CascadeMux I__4047 (
            .O(N__31136),
            .I(N__31133));
    InMux I__4046 (
            .O(N__31133),
            .I(N__31130));
    LocalMux I__4045 (
            .O(N__31130),
            .I(N__31127));
    Span4Mux_h I__4044 (
            .O(N__31127),
            .I(N__31124));
    Span4Mux_v I__4043 (
            .O(N__31124),
            .I(N__31120));
    InMux I__4042 (
            .O(N__31123),
            .I(N__31117));
    Odrv4 I__4041 (
            .O(N__31120),
            .I(controlWord_25));
    LocalMux I__4040 (
            .O(N__31117),
            .I(controlWord_25));
    IoInMux I__4039 (
            .O(N__31112),
            .I(N__31109));
    LocalMux I__4038 (
            .O(N__31109),
            .I(N__31106));
    Span4Mux_s3_v I__4037 (
            .O(N__31106),
            .I(N__31103));
    Span4Mux_h I__4036 (
            .O(N__31103),
            .I(N__31100));
    Sp12to4 I__4035 (
            .O(N__31100),
            .I(N__31097));
    Span12Mux_h I__4034 (
            .O(N__31097),
            .I(N__31093));
    InMux I__4033 (
            .O(N__31096),
            .I(N__31090));
    Odrv12 I__4032 (
            .O(N__31093),
            .I(A9_c));
    LocalMux I__4031 (
            .O(N__31090),
            .I(A9_c));
    CascadeMux I__4030 (
            .O(N__31085),
            .I(N__31081));
    InMux I__4029 (
            .O(N__31084),
            .I(N__31078));
    InMux I__4028 (
            .O(N__31081),
            .I(N__31075));
    LocalMux I__4027 (
            .O(N__31078),
            .I(N__31072));
    LocalMux I__4026 (
            .O(N__31075),
            .I(N__31069));
    Span4Mux_v I__4025 (
            .O(N__31072),
            .I(N__31066));
    Span4Mux_v I__4024 (
            .O(N__31069),
            .I(N__31063));
    Odrv4 I__4023 (
            .O(N__31066),
            .I(controlWord_24));
    Odrv4 I__4022 (
            .O(N__31063),
            .I(controlWord_24));
    IoInMux I__4021 (
            .O(N__31058),
            .I(N__31055));
    LocalMux I__4020 (
            .O(N__31055),
            .I(N__31052));
    Span4Mux_s3_h I__4019 (
            .O(N__31052),
            .I(N__31049));
    Span4Mux_h I__4018 (
            .O(N__31049),
            .I(N__31046));
    Span4Mux_h I__4017 (
            .O(N__31046),
            .I(N__31043));
    Span4Mux_h I__4016 (
            .O(N__31043),
            .I(N__31040));
    Span4Mux_h I__4015 (
            .O(N__31040),
            .I(N__31036));
    InMux I__4014 (
            .O(N__31039),
            .I(N__31033));
    Odrv4 I__4013 (
            .O(N__31036),
            .I(A8_c));
    LocalMux I__4012 (
            .O(N__31033),
            .I(A8_c));
    InMux I__4011 (
            .O(N__31028),
            .I(N__31025));
    LocalMux I__4010 (
            .O(N__31025),
            .I(N__31022));
    Span4Mux_h I__4009 (
            .O(N__31022),
            .I(N__31019));
    Span4Mux_v I__4008 (
            .O(N__31019),
            .I(N__31016));
    Span4Mux_v I__4007 (
            .O(N__31016),
            .I(N__31013));
    Odrv4 I__4006 (
            .O(N__31013),
            .I(gpuOut_c_0));
    InMux I__4005 (
            .O(N__31010),
            .I(N__31007));
    LocalMux I__4004 (
            .O(N__31007),
            .I(N__31004));
    Span12Mux_v I__4003 (
            .O(N__31004),
            .I(N__31001));
    Odrv12 I__4002 (
            .O(N__31001),
            .I(D0_in_c));
    CascadeMux I__4001 (
            .O(N__30998),
            .I(\CONTROL.N_161_cascade_ ));
    CascadeMux I__4000 (
            .O(N__30995),
            .I(N__30989));
    InMux I__3999 (
            .O(N__30994),
            .I(N__30984));
    InMux I__3998 (
            .O(N__30993),
            .I(N__30984));
    InMux I__3997 (
            .O(N__30992),
            .I(N__30979));
    InMux I__3996 (
            .O(N__30989),
            .I(N__30979));
    LocalMux I__3995 (
            .O(N__30984),
            .I(N__30976));
    LocalMux I__3994 (
            .O(N__30979),
            .I(N__30973));
    Span4Mux_h I__3993 (
            .O(N__30976),
            .I(N__30970));
    Span4Mux_h I__3992 (
            .O(N__30973),
            .I(N__30967));
    Odrv4 I__3991 (
            .O(N__30970),
            .I(\PROM.ROMDATA.m520 ));
    Odrv4 I__3990 (
            .O(N__30967),
            .I(\PROM.ROMDATA.m520 ));
    InMux I__3989 (
            .O(N__30962),
            .I(N__30959));
    LocalMux I__3988 (
            .O(N__30959),
            .I(N__30956));
    Span4Mux_v I__3987 (
            .O(N__30956),
            .I(N__30953));
    Span4Mux_v I__3986 (
            .O(N__30953),
            .I(N__30950));
    Sp12to4 I__3985 (
            .O(N__30950),
            .I(N__30947));
    Span12Mux_h I__3984 (
            .O(N__30947),
            .I(N__30944));
    Odrv12 I__3983 (
            .O(N__30944),
            .I(gpuOut_c_15));
    InMux I__3982 (
            .O(N__30941),
            .I(N__30938));
    LocalMux I__3981 (
            .O(N__30938),
            .I(N_176));
    CascadeMux I__3980 (
            .O(N__30935),
            .I(N__30931));
    InMux I__3979 (
            .O(N__30934),
            .I(N__30928));
    InMux I__3978 (
            .O(N__30931),
            .I(N__30925));
    LocalMux I__3977 (
            .O(N__30928),
            .I(N__30922));
    LocalMux I__3976 (
            .O(N__30925),
            .I(N__30919));
    Span4Mux_h I__3975 (
            .O(N__30922),
            .I(N__30916));
    Span4Mux_v I__3974 (
            .O(N__30919),
            .I(N__30913));
    Span4Mux_v I__3973 (
            .O(N__30916),
            .I(N__30910));
    Span4Mux_v I__3972 (
            .O(N__30913),
            .I(N__30907));
    Span4Mux_v I__3971 (
            .O(N__30910),
            .I(N__30904));
    Span4Mux_h I__3970 (
            .O(N__30907),
            .I(N__30901));
    Span4Mux_h I__3969 (
            .O(N__30904),
            .I(N__30898));
    IoSpan4Mux I__3968 (
            .O(N__30901),
            .I(N__30895));
    Odrv4 I__3967 (
            .O(N__30898),
            .I(D15_in_c));
    Odrv4 I__3966 (
            .O(N__30895),
            .I(D15_in_c));
    CascadeMux I__3965 (
            .O(N__30890),
            .I(N_176_cascade_));
    CascadeMux I__3964 (
            .O(N__30887),
            .I(\CONTROL.N_89_cascade_ ));
    CascadeMux I__3963 (
            .O(N__30884),
            .I(\CONTROL.aluReadBus_1_sqmuxa_0_a2_0Z0Z_0_cascade_ ));
    InMux I__3962 (
            .O(N__30881),
            .I(N__30872));
    InMux I__3961 (
            .O(N__30880),
            .I(N__30872));
    InMux I__3960 (
            .O(N__30879),
            .I(N__30872));
    LocalMux I__3959 (
            .O(N__30872),
            .I(\CONTROL.aluReadBus_1_sqmuxa_0_o2_0_0 ));
    InMux I__3958 (
            .O(N__30869),
            .I(N__30866));
    LocalMux I__3957 (
            .O(N__30866),
            .I(N__30863));
    Span4Mux_h I__3956 (
            .O(N__30863),
            .I(N__30860));
    Sp12to4 I__3955 (
            .O(N__30860),
            .I(N__30857));
    Odrv12 I__3954 (
            .O(N__30857),
            .I(gpuOut_c_10));
    InMux I__3953 (
            .O(N__30854),
            .I(N__30851));
    LocalMux I__3952 (
            .O(N__30851),
            .I(N__30848));
    Span4Mux_v I__3951 (
            .O(N__30848),
            .I(N__30845));
    Span4Mux_v I__3950 (
            .O(N__30845),
            .I(N__30842));
    Span4Mux_v I__3949 (
            .O(N__30842),
            .I(N__30839));
    Odrv4 I__3948 (
            .O(N__30839),
            .I(D10_in_c));
    CascadeMux I__3947 (
            .O(N__30836),
            .I(\CONTROL.N_171_cascade_ ));
    InMux I__3946 (
            .O(N__30833),
            .I(N__30830));
    LocalMux I__3945 (
            .O(N__30830),
            .I(N__30827));
    Span4Mux_v I__3944 (
            .O(N__30827),
            .I(N__30824));
    Odrv4 I__3943 (
            .O(N__30824),
            .I(\CONTROL.N_187 ));
    CascadeMux I__3942 (
            .O(N__30821),
            .I(\CONTROL.un1_busState12_2_i_a2_0_1_tz_0_cascade_ ));
    CascadeMux I__3941 (
            .O(N__30818),
            .I(\CONTROL.N_244_cascade_ ));
    InMux I__3940 (
            .O(N__30815),
            .I(N__30812));
    LocalMux I__3939 (
            .O(N__30812),
            .I(\CONTROL.un1_busState14_1_i_o2_0 ));
    InMux I__3938 (
            .O(N__30809),
            .I(N__30806));
    LocalMux I__3937 (
            .O(N__30806),
            .I(N__30803));
    Odrv4 I__3936 (
            .O(N__30803),
            .I(\CONTROL.aluReadBus_r_1 ));
    InMux I__3935 (
            .O(N__30800),
            .I(N__30797));
    LocalMux I__3934 (
            .O(N__30797),
            .I(\CONTROL.un1_busState14_1_i_a2_1_iZ0Z_1 ));
    InMux I__3933 (
            .O(N__30794),
            .I(N__30784));
    InMux I__3932 (
            .O(N__30793),
            .I(N__30784));
    InMux I__3931 (
            .O(N__30792),
            .I(N__30781));
    InMux I__3930 (
            .O(N__30791),
            .I(N__30778));
    InMux I__3929 (
            .O(N__30790),
            .I(N__30773));
    InMux I__3928 (
            .O(N__30789),
            .I(N__30773));
    LocalMux I__3927 (
            .O(N__30784),
            .I(N__30770));
    LocalMux I__3926 (
            .O(N__30781),
            .I(\CONTROL.N_244 ));
    LocalMux I__3925 (
            .O(N__30778),
            .I(\CONTROL.N_244 ));
    LocalMux I__3924 (
            .O(N__30773),
            .I(\CONTROL.N_244 ));
    Odrv4 I__3923 (
            .O(N__30770),
            .I(\CONTROL.N_244 ));
    CEMux I__3922 (
            .O(N__30761),
            .I(N__30756));
    CEMux I__3921 (
            .O(N__30760),
            .I(N__30753));
    CEMux I__3920 (
            .O(N__30759),
            .I(N__30749));
    LocalMux I__3919 (
            .O(N__30756),
            .I(N__30746));
    LocalMux I__3918 (
            .O(N__30753),
            .I(N__30743));
    CEMux I__3917 (
            .O(N__30752),
            .I(N__30740));
    LocalMux I__3916 (
            .O(N__30749),
            .I(N__30736));
    Span4Mux_v I__3915 (
            .O(N__30746),
            .I(N__30729));
    Span4Mux_h I__3914 (
            .O(N__30743),
            .I(N__30729));
    LocalMux I__3913 (
            .O(N__30740),
            .I(N__30729));
    CEMux I__3912 (
            .O(N__30739),
            .I(N__30726));
    Span4Mux_v I__3911 (
            .O(N__30736),
            .I(N__30723));
    Span4Mux_h I__3910 (
            .O(N__30729),
            .I(N__30720));
    LocalMux I__3909 (
            .O(N__30726),
            .I(N__30717));
    Span4Mux_v I__3908 (
            .O(N__30723),
            .I(N__30714));
    Odrv4 I__3907 (
            .O(N__30720),
            .I(\CONTROL.N_58 ));
    Odrv12 I__3906 (
            .O(N__30717),
            .I(\CONTROL.N_58 ));
    Odrv4 I__3905 (
            .O(N__30714),
            .I(\CONTROL.N_58 ));
    InMux I__3904 (
            .O(N__30707),
            .I(N__30704));
    LocalMux I__3903 (
            .O(N__30704),
            .I(\CONTROL.N_89 ));
    InMux I__3902 (
            .O(N__30701),
            .I(N__30698));
    LocalMux I__3901 (
            .O(N__30698),
            .I(N__30695));
    Span4Mux_v I__3900 (
            .O(N__30695),
            .I(N__30692));
    Span4Mux_v I__3899 (
            .O(N__30692),
            .I(N__30689));
    Span4Mux_v I__3898 (
            .O(N__30689),
            .I(N__30686));
    IoSpan4Mux I__3897 (
            .O(N__30686),
            .I(N__30683));
    Odrv4 I__3896 (
            .O(N__30683),
            .I(D11_in_c));
    CascadeMux I__3895 (
            .O(N__30680),
            .I(\CONTROL.N_172_cascade_ ));
    InMux I__3894 (
            .O(N__30677),
            .I(N__30674));
    LocalMux I__3893 (
            .O(N__30674),
            .I(N__30671));
    Odrv4 I__3892 (
            .O(N__30671),
            .I(N_188));
    InMux I__3891 (
            .O(N__30668),
            .I(N__30665));
    LocalMux I__3890 (
            .O(N__30665),
            .I(N__30661));
    InMux I__3889 (
            .O(N__30664),
            .I(N__30658));
    Odrv4 I__3888 (
            .O(N__30661),
            .I(N_204));
    LocalMux I__3887 (
            .O(N__30658),
            .I(N_204));
    CascadeMux I__3886 (
            .O(N__30653),
            .I(N_188_cascade_));
    InMux I__3885 (
            .O(N__30650),
            .I(N__30647));
    LocalMux I__3884 (
            .O(N__30647),
            .I(N__30644));
    Span4Mux_v I__3883 (
            .O(N__30644),
            .I(N__30640));
    InMux I__3882 (
            .O(N__30643),
            .I(N__30637));
    Odrv4 I__3881 (
            .O(N__30640),
            .I(\CONTROL.ctrlOut_11 ));
    LocalMux I__3880 (
            .O(N__30637),
            .I(\CONTROL.ctrlOut_11 ));
    InMux I__3879 (
            .O(N__30632),
            .I(N__30629));
    LocalMux I__3878 (
            .O(N__30629),
            .I(N__30626));
    Span4Mux_h I__3877 (
            .O(N__30626),
            .I(N__30623));
    Span4Mux_v I__3876 (
            .O(N__30623),
            .I(N__30620));
    Span4Mux_v I__3875 (
            .O(N__30620),
            .I(N__30617));
    Span4Mux_v I__3874 (
            .O(N__30617),
            .I(N__30614));
    Odrv4 I__3873 (
            .O(N__30614),
            .I(gpuOut_c_12));
    InMux I__3872 (
            .O(N__30611),
            .I(N__30608));
    LocalMux I__3871 (
            .O(N__30608),
            .I(N__30605));
    Span4Mux_v I__3870 (
            .O(N__30605),
            .I(N__30602));
    Span4Mux_v I__3869 (
            .O(N__30602),
            .I(N__30599));
    Span4Mux_v I__3868 (
            .O(N__30599),
            .I(N__30596));
    Span4Mux_h I__3867 (
            .O(N__30596),
            .I(N__30593));
    Odrv4 I__3866 (
            .O(N__30593),
            .I(D12_in_c));
    CascadeMux I__3865 (
            .O(N__30590),
            .I(\CONTROL.N_173_cascade_ ));
    InMux I__3864 (
            .O(N__30587),
            .I(N__30584));
    LocalMux I__3863 (
            .O(N__30584),
            .I(\CONTROL.N_189 ));
    CascadeMux I__3862 (
            .O(N__30581),
            .I(\CONTROL.un1_busState14_1_i_o2_0_cascade_ ));
    CascadeMux I__3861 (
            .O(N__30578),
            .I(\CONTROL.busState_1_RNIRA1I6Z0Z_2_cascade_ ));
    CascadeMux I__3860 (
            .O(N__30575),
            .I(N__30572));
    InMux I__3859 (
            .O(N__30572),
            .I(N__30569));
    LocalMux I__3858 (
            .O(N__30569),
            .I(N__30566));
    Span4Mux_v I__3857 (
            .O(N__30566),
            .I(N__30563));
    Odrv4 I__3856 (
            .O(N__30563),
            .I(\ALU.d_RNI8VHNHZ0Z_1 ));
    CascadeMux I__3855 (
            .O(N__30560),
            .I(\ALU.dout_3_ns_1_12_cascade_ ));
    CascadeMux I__3854 (
            .O(N__30557),
            .I(\ALU.dout_6_ns_1_12_cascade_ ));
    InMux I__3853 (
            .O(N__30554),
            .I(N__30551));
    LocalMux I__3852 (
            .O(N__30551),
            .I(\ALU.N_1097 ));
    CascadeMux I__3851 (
            .O(N__30548),
            .I(\ALU.N_1145_cascade_ ));
    CascadeMux I__3850 (
            .O(N__30545),
            .I(aluOut_12_cascade_));
    InMux I__3849 (
            .O(N__30542),
            .I(N__30536));
    InMux I__3848 (
            .O(N__30541),
            .I(N__30536));
    LocalMux I__3847 (
            .O(N__30536),
            .I(N__30533));
    Span4Mux_h I__3846 (
            .O(N__30533),
            .I(N__30530));
    Odrv4 I__3845 (
            .O(N__30530),
            .I(\CONTROL.bus_0_12 ));
    InMux I__3844 (
            .O(N__30527),
            .I(N__30524));
    LocalMux I__3843 (
            .O(N__30524),
            .I(N__30521));
    Span4Mux_h I__3842 (
            .O(N__30521),
            .I(N__30518));
    Span4Mux_v I__3841 (
            .O(N__30518),
            .I(N__30515));
    Span4Mux_v I__3840 (
            .O(N__30515),
            .I(N__30512));
    Span4Mux_v I__3839 (
            .O(N__30512),
            .I(N__30509));
    Span4Mux_h I__3838 (
            .O(N__30509),
            .I(N__30506));
    Odrv4 I__3837 (
            .O(N__30506),
            .I(gpuOut_c_11));
    CascadeMux I__3836 (
            .O(N__30503),
            .I(N__30500));
    InMux I__3835 (
            .O(N__30500),
            .I(N__30497));
    LocalMux I__3834 (
            .O(N__30497),
            .I(N__30494));
    Odrv12 I__3833 (
            .O(N__30494),
            .I(\ALU.mult_5_c_RNOZ0Z_0 ));
    InMux I__3832 (
            .O(N__30491),
            .I(N__30485));
    InMux I__3831 (
            .O(N__30490),
            .I(N__30485));
    LocalMux I__3830 (
            .O(N__30485),
            .I(N__30482));
    Span4Mux_h I__3829 (
            .O(N__30482),
            .I(N__30479));
    Span4Mux_h I__3828 (
            .O(N__30479),
            .I(N__30476));
    Odrv4 I__3827 (
            .O(N__30476),
            .I(\DROM.ROMDATA.dintern_0_0_NEW_0 ));
    InMux I__3826 (
            .O(N__30473),
            .I(N__30470));
    LocalMux I__3825 (
            .O(N__30470),
            .I(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_0 ));
    InMux I__3824 (
            .O(N__30467),
            .I(N__30464));
    LocalMux I__3823 (
            .O(N__30464),
            .I(N__30461));
    Span12Mux_v I__3822 (
            .O(N__30461),
            .I(N__30458));
    Span12Mux_h I__3821 (
            .O(N__30458),
            .I(N__30455));
    Odrv12 I__3820 (
            .O(N__30455),
            .I(gpuOut_c_14));
    InMux I__3819 (
            .O(N__30452),
            .I(N__30449));
    LocalMux I__3818 (
            .O(N__30449),
            .I(N__30446));
    Span12Mux_h I__3817 (
            .O(N__30446),
            .I(N__30442));
    InMux I__3816 (
            .O(N__30445),
            .I(N__30439));
    Odrv12 I__3815 (
            .O(N__30442),
            .I(\CONTROL.ctrlOut_14 ));
    LocalMux I__3814 (
            .O(N__30439),
            .I(\CONTROL.ctrlOut_14 ));
    InMux I__3813 (
            .O(N__30434),
            .I(N__30431));
    LocalMux I__3812 (
            .O(N__30431),
            .I(N__30428));
    Span4Mux_h I__3811 (
            .O(N__30428),
            .I(N__30425));
    Span4Mux_h I__3810 (
            .O(N__30425),
            .I(N__30422));
    Sp12to4 I__3809 (
            .O(N__30422),
            .I(N__30419));
    Span12Mux_v I__3808 (
            .O(N__30419),
            .I(N__30416));
    Odrv12 I__3807 (
            .O(N__30416),
            .I(D14_in_c));
    CascadeMux I__3806 (
            .O(N__30413),
            .I(\CONTROL.N_175_cascade_ ));
    CascadeMux I__3805 (
            .O(N__30410),
            .I(N_191_cascade_));
    CascadeMux I__3804 (
            .O(N__30407),
            .I(N__30403));
    InMux I__3803 (
            .O(N__30406),
            .I(N__30400));
    InMux I__3802 (
            .O(N__30403),
            .I(N__30397));
    LocalMux I__3801 (
            .O(N__30400),
            .I(N__30394));
    LocalMux I__3800 (
            .O(N__30397),
            .I(N__30391));
    Span4Mux_h I__3799 (
            .O(N__30394),
            .I(N__30388));
    Span4Mux_h I__3798 (
            .O(N__30391),
            .I(N__30383));
    Span4Mux_v I__3797 (
            .O(N__30388),
            .I(N__30383));
    Span4Mux_v I__3796 (
            .O(N__30383),
            .I(N__30380));
    Odrv4 I__3795 (
            .O(N__30380),
            .I(CONTROL_addrstack_reto_11));
    InMux I__3794 (
            .O(N__30377),
            .I(N__30374));
    LocalMux I__3793 (
            .O(N__30374),
            .I(N__30370));
    InMux I__3792 (
            .O(N__30373),
            .I(N__30367));
    Span4Mux_v I__3791 (
            .O(N__30370),
            .I(N__30364));
    LocalMux I__3790 (
            .O(N__30367),
            .I(N__30361));
    Span4Mux_v I__3789 (
            .O(N__30364),
            .I(N__30358));
    Span4Mux_v I__3788 (
            .O(N__30361),
            .I(N__30355));
    Odrv4 I__3787 (
            .O(N__30358),
            .I(N_426));
    Odrv4 I__3786 (
            .O(N__30355),
            .I(N_426));
    InMux I__3785 (
            .O(N__30350),
            .I(N__30347));
    LocalMux I__3784 (
            .O(N__30347),
            .I(N__30343));
    InMux I__3783 (
            .O(N__30346),
            .I(N__30340));
    Span4Mux_v I__3782 (
            .O(N__30343),
            .I(N__30335));
    LocalMux I__3781 (
            .O(N__30340),
            .I(N__30335));
    Span4Mux_v I__3780 (
            .O(N__30335),
            .I(N__30332));
    Span4Mux_h I__3779 (
            .O(N__30332),
            .I(N__30329));
    Odrv4 I__3778 (
            .O(N__30329),
            .I(progRomAddress_11));
    InMux I__3777 (
            .O(N__30326),
            .I(N__30323));
    LocalMux I__3776 (
            .O(N__30323),
            .I(N__30320));
    Span4Mux_v I__3775 (
            .O(N__30320),
            .I(N__30317));
    Odrv4 I__3774 (
            .O(N__30317),
            .I(\ALU.d_RNILJMRC1_0Z0Z_8 ));
    CascadeMux I__3773 (
            .O(N__30314),
            .I(\ALU.combOperand2_1Z0Z_0_cascade_ ));
    InMux I__3772 (
            .O(N__30311),
            .I(N__30308));
    LocalMux I__3771 (
            .O(N__30308),
            .I(N__30305));
    Span4Mux_v I__3770 (
            .O(N__30305),
            .I(N__30302));
    Odrv4 I__3769 (
            .O(N__30302),
            .I(dintern_adflt_3_x));
    CascadeMux I__3768 (
            .O(N__30299),
            .I(DROM_ROMDATA_dintern_0ro_cascade_));
    InMux I__3767 (
            .O(N__30296),
            .I(N__30293));
    LocalMux I__3766 (
            .O(N__30293),
            .I(N__30290));
    Span4Mux_h I__3765 (
            .O(N__30290),
            .I(N__30287));
    Odrv4 I__3764 (
            .O(N__30287),
            .I(\CONTROL.bus_6_a0_sx_0 ));
    InMux I__3763 (
            .O(N__30284),
            .I(N__30281));
    LocalMux I__3762 (
            .O(N__30281),
            .I(\ALU.mult_3_c14_THRU_CO ));
    CascadeMux I__3761 (
            .O(N__30278),
            .I(N__30275));
    InMux I__3760 (
            .O(N__30275),
            .I(N__30272));
    LocalMux I__3759 (
            .O(N__30272),
            .I(N__30269));
    Span4Mux_h I__3758 (
            .O(N__30269),
            .I(N__30266));
    Odrv4 I__3757 (
            .O(N__30266),
            .I(\ALU.d_RNI3D2O61Z0Z_2 ));
    InMux I__3756 (
            .O(N__30263),
            .I(\ALU.mult_1_c14 ));
    InMux I__3755 (
            .O(N__30260),
            .I(N__30257));
    LocalMux I__3754 (
            .O(N__30257),
            .I(\ALU.d_RNI83GO51Z0Z_0 ));
    CascadeMux I__3753 (
            .O(N__30254),
            .I(N__30251));
    InMux I__3752 (
            .O(N__30251),
            .I(N__30248));
    LocalMux I__3751 (
            .O(N__30248),
            .I(\ALU.d_RNIPIBO31Z0Z_0 ));
    InMux I__3750 (
            .O(N__30245),
            .I(N__30242));
    LocalMux I__3749 (
            .O(N__30242),
            .I(N__30239));
    Odrv4 I__3748 (
            .O(N__30239),
            .I(\ALU.d_RNIIHC6LZ0Z_3 ));
    InMux I__3747 (
            .O(N__30236),
            .I(N__30233));
    LocalMux I__3746 (
            .O(N__30233),
            .I(\ALU.d_RNITH0K51Z0Z_0 ));
    InMux I__3745 (
            .O(N__30230),
            .I(N__30227));
    LocalMux I__3744 (
            .O(N__30227),
            .I(N__30224));
    Odrv4 I__3743 (
            .O(N__30224),
            .I(\ALU.d_RNI0H41KZ0Z_1 ));
    CascadeMux I__3742 (
            .O(N__30221),
            .I(N__30218));
    InMux I__3741 (
            .O(N__30218),
            .I(N__30215));
    LocalMux I__3740 (
            .O(N__30215),
            .I(\ALU.d_RNIETL861Z0Z_0 ));
    InMux I__3739 (
            .O(N__30212),
            .I(N__30209));
    LocalMux I__3738 (
            .O(N__30209),
            .I(\ALU.d_RNI8FM541Z0Z_0 ));
    InMux I__3737 (
            .O(N__30206),
            .I(N__30203));
    LocalMux I__3736 (
            .O(N__30203),
            .I(N__30200));
    Odrv4 I__3735 (
            .O(N__30200),
            .I(\ALU.d_RNIGIF4D1Z0Z_2 ));
    CascadeMux I__3734 (
            .O(N__30197),
            .I(N__30194));
    InMux I__3733 (
            .O(N__30194),
            .I(N__30191));
    LocalMux I__3732 (
            .O(N__30191),
            .I(N__30188));
    Odrv4 I__3731 (
            .O(N__30188),
            .I(\ALU.d_RNIRJ3VHZ0Z_1 ));
    InMux I__3730 (
            .O(N__30185),
            .I(\ALU.mult_1_c6 ));
    InMux I__3729 (
            .O(N__30182),
            .I(N__30179));
    LocalMux I__3728 (
            .O(N__30179),
            .I(N__30176));
    Span4Mux_h I__3727 (
            .O(N__30176),
            .I(N__30173));
    Odrv4 I__3726 (
            .O(N__30173),
            .I(\ALU.d_RNI990621Z0Z_0 ));
    InMux I__3725 (
            .O(N__30170),
            .I(\ALU.mult_1_c7 ));
    InMux I__3724 (
            .O(N__30167),
            .I(N__30164));
    LocalMux I__3723 (
            .O(N__30164),
            .I(\ALU.d_RNIH49MHZ0Z_1 ));
    InMux I__3722 (
            .O(N__30161),
            .I(bfn_13_12_0_));
    CascadeMux I__3721 (
            .O(N__30158),
            .I(N__30155));
    InMux I__3720 (
            .O(N__30155),
            .I(N__30152));
    LocalMux I__3719 (
            .O(N__30152),
            .I(N__30149));
    Odrv4 I__3718 (
            .O(N__30149),
            .I(\ALU.d_RNISP66IZ0Z_1 ));
    InMux I__3717 (
            .O(N__30146),
            .I(\ALU.mult_1_c9 ));
    InMux I__3716 (
            .O(N__30143),
            .I(N__30140));
    LocalMux I__3715 (
            .O(N__30140),
            .I(N__30137));
    Span4Mux_h I__3714 (
            .O(N__30137),
            .I(N__30134));
    Odrv4 I__3713 (
            .O(N__30134),
            .I(\ALU.d_RNI0LDMJZ0Z_1 ));
    CascadeMux I__3712 (
            .O(N__30131),
            .I(N__30128));
    InMux I__3711 (
            .O(N__30128),
            .I(N__30125));
    LocalMux I__3710 (
            .O(N__30125),
            .I(\ALU.d_RNIK8R951Z0Z_0 ));
    InMux I__3709 (
            .O(N__30122),
            .I(\ALU.mult_1_c10 ));
    InMux I__3708 (
            .O(N__30119),
            .I(\ALU.mult_1_c11 ));
    InMux I__3707 (
            .O(N__30116),
            .I(N__30113));
    LocalMux I__3706 (
            .O(N__30113),
            .I(N__30110));
    Span4Mux_v I__3705 (
            .O(N__30110),
            .I(N__30107));
    Odrv4 I__3704 (
            .O(N__30107),
            .I(\ALU.d_RNI9UI0KZ0Z_1 ));
    InMux I__3703 (
            .O(N__30104),
            .I(\ALU.mult_1_c12 ));
    InMux I__3702 (
            .O(N__30101),
            .I(\ALU.mult_1_c13 ));
    CascadeMux I__3701 (
            .O(N__30098),
            .I(N__30095));
    InMux I__3700 (
            .O(N__30095),
            .I(N__30092));
    LocalMux I__3699 (
            .O(N__30092),
            .I(N__30089));
    Odrv4 I__3698 (
            .O(N__30089),
            .I(\ALU.d_RNIA6P2IZ0Z_7 ));
    InMux I__3697 (
            .O(N__30086),
            .I(\ALU.mult_1_c1 ));
    CascadeMux I__3696 (
            .O(N__30083),
            .I(N__30080));
    InMux I__3695 (
            .O(N__30080),
            .I(N__30077));
    LocalMux I__3694 (
            .O(N__30077),
            .I(\ALU.d_RNIFBJI61Z0Z_0 ));
    InMux I__3693 (
            .O(N__30074),
            .I(\ALU.mult_1_c2 ));
    InMux I__3692 (
            .O(N__30071),
            .I(N__30068));
    LocalMux I__3691 (
            .O(N__30068),
            .I(\ALU.d_RNIIOGRGZ0Z_1 ));
    CascadeMux I__3690 (
            .O(N__30065),
            .I(N__30062));
    InMux I__3689 (
            .O(N__30062),
            .I(N__30059));
    LocalMux I__3688 (
            .O(N__30059),
            .I(N__30056));
    Span4Mux_h I__3687 (
            .O(N__30056),
            .I(N__30053));
    Odrv4 I__3686 (
            .O(N__30053),
            .I(\ALU.d_RNI67HQ21Z0Z_0 ));
    InMux I__3685 (
            .O(N__30050),
            .I(\ALU.mult_1_c3 ));
    InMux I__3684 (
            .O(N__30047),
            .I(N__30044));
    LocalMux I__3683 (
            .O(N__30044),
            .I(N__30041));
    Span4Mux_h I__3682 (
            .O(N__30041),
            .I(N__30038));
    Odrv4 I__3681 (
            .O(N__30038),
            .I(\ALU.d_RNI8Q43IZ0Z_1 ));
    CascadeMux I__3680 (
            .O(N__30035),
            .I(N__30032));
    InMux I__3679 (
            .O(N__30032),
            .I(N__30029));
    LocalMux I__3678 (
            .O(N__30029),
            .I(N__30026));
    Odrv4 I__3677 (
            .O(N__30026),
            .I(\ALU.d_RNIITFA41Z0Z_0 ));
    InMux I__3676 (
            .O(N__30023),
            .I(\ALU.mult_1_c4 ));
    InMux I__3675 (
            .O(N__30020),
            .I(N__30017));
    LocalMux I__3674 (
            .O(N__30017),
            .I(N__30014));
    Span4Mux_h I__3673 (
            .O(N__30014),
            .I(N__30011));
    Odrv4 I__3672 (
            .O(N__30011),
            .I(\ALU.d_RNI5NE641Z0Z_0 ));
    CascadeMux I__3671 (
            .O(N__30008),
            .I(N__30005));
    InMux I__3670 (
            .O(N__30005),
            .I(N__30002));
    LocalMux I__3669 (
            .O(N__30002),
            .I(N__29999));
    Odrv12 I__3668 (
            .O(N__29999),
            .I(\ALU.d_RNIUEFBIZ0Z_1 ));
    InMux I__3667 (
            .O(N__29996),
            .I(\ALU.mult_1_c5 ));
    InMux I__3666 (
            .O(N__29993),
            .I(N__29990));
    LocalMux I__3665 (
            .O(N__29990),
            .I(\ALU.d_RNIUFQIGZ0Z_7 ));
    CascadeMux I__3664 (
            .O(N__29987),
            .I(N__29984));
    InMux I__3663 (
            .O(N__29984),
            .I(N__29981));
    LocalMux I__3662 (
            .O(N__29981),
            .I(N__29978));
    Span4Mux_v I__3661 (
            .O(N__29978),
            .I(N__29975));
    Span4Mux_h I__3660 (
            .O(N__29975),
            .I(N__29972));
    Odrv4 I__3659 (
            .O(N__29972),
            .I(\ALU.d_RNI8JFO21Z0Z_6 ));
    InMux I__3658 (
            .O(N__29969),
            .I(\ALU.mult_7_c9 ));
    InMux I__3657 (
            .O(N__29966),
            .I(N__29963));
    LocalMux I__3656 (
            .O(N__29963),
            .I(N__29960));
    Span4Mux_h I__3655 (
            .O(N__29960),
            .I(N__29957));
    Span4Mux_v I__3654 (
            .O(N__29957),
            .I(N__29954));
    Odrv4 I__3653 (
            .O(N__29954),
            .I(\ALU.d_RNIKHEQHZ0Z_7 ));
    CascadeMux I__3652 (
            .O(N__29951),
            .I(N__29948));
    InMux I__3651 (
            .O(N__29948),
            .I(N__29945));
    LocalMux I__3650 (
            .O(N__29945),
            .I(N__29942));
    Span4Mux_v I__3649 (
            .O(N__29942),
            .I(N__29939));
    Sp12to4 I__3648 (
            .O(N__29939),
            .I(N__29936));
    Odrv12 I__3647 (
            .O(N__29936),
            .I(\ALU.d_RNIK9E841Z0Z_6 ));
    InMux I__3646 (
            .O(N__29933),
            .I(\ALU.mult_7_c10 ));
    InMux I__3645 (
            .O(N__29930),
            .I(N__29927));
    LocalMux I__3644 (
            .O(N__29927),
            .I(N__29924));
    Span4Mux_v I__3643 (
            .O(N__29924),
            .I(N__29921));
    Span4Mux_h I__3642 (
            .O(N__29921),
            .I(N__29918));
    Odrv4 I__3641 (
            .O(N__29918),
            .I(\ALU.d_RNI73D441Z0Z_6 ));
    InMux I__3640 (
            .O(N__29915),
            .I(\ALU.mult_7_c11 ));
    InMux I__3639 (
            .O(N__29912),
            .I(N__29909));
    LocalMux I__3638 (
            .O(N__29909),
            .I(N__29906));
    Span4Mux_v I__3637 (
            .O(N__29906),
            .I(N__29903));
    Odrv4 I__3636 (
            .O(N__29903),
            .I(\ALU.d_RNI7BDMHZ0Z_7 ));
    InMux I__3635 (
            .O(N__29900),
            .I(\ALU.mult_7_c12 ));
    InMux I__3634 (
            .O(N__29897),
            .I(N__29894));
    LocalMux I__3633 (
            .O(N__29894),
            .I(N__29891));
    Span4Mux_v I__3632 (
            .O(N__29891),
            .I(N__29888));
    Odrv4 I__3631 (
            .O(N__29888),
            .I(\ALU.d_RNIBLU321Z0Z_6 ));
    InMux I__3630 (
            .O(N__29885),
            .I(\ALU.mult_7_c13 ));
    InMux I__3629 (
            .O(N__29882),
            .I(bfn_13_10_0_));
    CascadeMux I__3628 (
            .O(N__29879),
            .I(N__29876));
    InMux I__3627 (
            .O(N__29876),
            .I(N__29873));
    LocalMux I__3626 (
            .O(N__29873),
            .I(\ALU.d_RNIHNHG61Z0Z_6 ));
    CascadeMux I__3625 (
            .O(N__29870),
            .I(N__29867));
    InMux I__3624 (
            .O(N__29867),
            .I(N__29864));
    LocalMux I__3623 (
            .O(N__29864),
            .I(\ALU.d_RNI4LU7E1Z0Z_6 ));
    CascadeMux I__3622 (
            .O(N__29861),
            .I(\ALU.d_RNILJMRC1Z0Z_8_cascade_ ));
    InMux I__3621 (
            .O(N__29858),
            .I(\ALU.mult_7_c7 ));
    InMux I__3620 (
            .O(N__29855),
            .I(N__29852));
    LocalMux I__3619 (
            .O(N__29852),
            .I(\ALU.d_RNITLGILZ0Z_7 ));
    InMux I__3618 (
            .O(N__29849),
            .I(\ALU.mult_7_c8 ));
    InMux I__3617 (
            .O(N__29846),
            .I(N__29843));
    LocalMux I__3616 (
            .O(N__29843),
            .I(N__29839));
    InMux I__3615 (
            .O(N__29842),
            .I(N__29836));
    Span4Mux_v I__3614 (
            .O(N__29839),
            .I(N__29833));
    LocalMux I__3613 (
            .O(N__29836),
            .I(N__29830));
    Odrv4 I__3612 (
            .O(N__29833),
            .I(\CONTROL.programCounter_1_10 ));
    Odrv4 I__3611 (
            .O(N__29830),
            .I(\CONTROL.programCounter_1_10 ));
    InMux I__3610 (
            .O(N__29825),
            .I(N__29818));
    InMux I__3609 (
            .O(N__29824),
            .I(N__29815));
    InMux I__3608 (
            .O(N__29823),
            .I(N__29808));
    InMux I__3607 (
            .O(N__29822),
            .I(N__29808));
    InMux I__3606 (
            .O(N__29821),
            .I(N__29808));
    LocalMux I__3605 (
            .O(N__29818),
            .I(\CONTROL.programCounter11_reto_rep1 ));
    LocalMux I__3604 (
            .O(N__29815),
            .I(\CONTROL.programCounter11_reto_rep1 ));
    LocalMux I__3603 (
            .O(N__29808),
            .I(\CONTROL.programCounter11_reto_rep1 ));
    InMux I__3602 (
            .O(N__29801),
            .I(N__29798));
    LocalMux I__3601 (
            .O(N__29798),
            .I(\CONTROL.programCounter_1_reto_10 ));
    InMux I__3600 (
            .O(N__29795),
            .I(N__29792));
    LocalMux I__3599 (
            .O(N__29792),
            .I(\CONTROL.N_425 ));
    InMux I__3598 (
            .O(N__29789),
            .I(N__29786));
    LocalMux I__3597 (
            .O(N__29786),
            .I(N__29783));
    Span4Mux_h I__3596 (
            .O(N__29783),
            .I(N__29780));
    Odrv4 I__3595 (
            .O(N__29780),
            .I(\CONTROL.programCounter_1_axb_1 ));
    CascadeMux I__3594 (
            .O(N__29777),
            .I(N__29774));
    InMux I__3593 (
            .O(N__29774),
            .I(N__29771));
    LocalMux I__3592 (
            .O(N__29771),
            .I(N__29768));
    Odrv12 I__3591 (
            .O(N__29768),
            .I(\CONTROL.addrstackptr_8_1 ));
    CascadeMux I__3590 (
            .O(N__29765),
            .I(N__29762));
    InMux I__3589 (
            .O(N__29762),
            .I(N__29759));
    LocalMux I__3588 (
            .O(N__29759),
            .I(N__29756));
    Odrv12 I__3587 (
            .O(N__29756),
            .I(\CONTROL.addrstackptr_RNI19JNL91Z0Z_0 ));
    InMux I__3586 (
            .O(N__29753),
            .I(N__29750));
    LocalMux I__3585 (
            .O(N__29750),
            .I(\CONTROL.dout_reto_9 ));
    CascadeMux I__3584 (
            .O(N__29747),
            .I(N__29744));
    InMux I__3583 (
            .O(N__29744),
            .I(N__29741));
    LocalMux I__3582 (
            .O(N__29741),
            .I(N__29737));
    InMux I__3581 (
            .O(N__29740),
            .I(N__29734));
    Span4Mux_v I__3580 (
            .O(N__29737),
            .I(N__29731));
    LocalMux I__3579 (
            .O(N__29734),
            .I(progRomAddress_15));
    Odrv4 I__3578 (
            .O(N__29731),
            .I(progRomAddress_15));
    InMux I__3577 (
            .O(N__29726),
            .I(N__29723));
    LocalMux I__3576 (
            .O(N__29723),
            .I(N__29719));
    InMux I__3575 (
            .O(N__29722),
            .I(N__29716));
    Span4Mux_v I__3574 (
            .O(N__29719),
            .I(N__29713));
    LocalMux I__3573 (
            .O(N__29716),
            .I(\CONTROL.programCounter_1_11 ));
    Odrv4 I__3572 (
            .O(N__29713),
            .I(\CONTROL.programCounter_1_11 ));
    InMux I__3571 (
            .O(N__29708),
            .I(N__29704));
    InMux I__3570 (
            .O(N__29707),
            .I(N__29701));
    LocalMux I__3569 (
            .O(N__29704),
            .I(N__29695));
    LocalMux I__3568 (
            .O(N__29701),
            .I(N__29695));
    CascadeMux I__3567 (
            .O(N__29700),
            .I(N__29692));
    Span4Mux_v I__3566 (
            .O(N__29695),
            .I(N__29689));
    InMux I__3565 (
            .O(N__29692),
            .I(N__29686));
    Odrv4 I__3564 (
            .O(N__29689),
            .I(\CONTROL.addrstack_1_4 ));
    LocalMux I__3563 (
            .O(N__29686),
            .I(\CONTROL.addrstack_1_4 ));
    InMux I__3562 (
            .O(N__29681),
            .I(N__29678));
    LocalMux I__3561 (
            .O(N__29678),
            .I(\CONTROL.N_4_1 ));
    InMux I__3560 (
            .O(N__29675),
            .I(N__29671));
    InMux I__3559 (
            .O(N__29674),
            .I(N__29668));
    LocalMux I__3558 (
            .O(N__29671),
            .I(\CONTROL.un1_addrstackptr_c4_0 ));
    LocalMux I__3557 (
            .O(N__29668),
            .I(\CONTROL.un1_addrstackptr_c4_0 ));
    CascadeMux I__3556 (
            .O(N__29663),
            .I(N__29660));
    InMux I__3555 (
            .O(N__29660),
            .I(N__29657));
    LocalMux I__3554 (
            .O(N__29657),
            .I(N__29654));
    Span4Mux_h I__3553 (
            .O(N__29654),
            .I(N__29651));
    Odrv4 I__3552 (
            .O(N__29651),
            .I(\CONTROL.addrstackptr_8_4 ));
    InMux I__3551 (
            .O(N__29648),
            .I(N__29644));
    InMux I__3550 (
            .O(N__29647),
            .I(N__29641));
    LocalMux I__3549 (
            .O(N__29644),
            .I(N__29638));
    LocalMux I__3548 (
            .O(N__29641),
            .I(\CONTROL.programCounter_1_14 ));
    Odrv4 I__3547 (
            .O(N__29638),
            .I(\CONTROL.programCounter_1_14 ));
    InMux I__3546 (
            .O(N__29633),
            .I(N__29630));
    LocalMux I__3545 (
            .O(N__29630),
            .I(\CONTROL.programCounter_1_reto_14 ));
    InMux I__3544 (
            .O(N__29627),
            .I(N__29624));
    LocalMux I__3543 (
            .O(N__29624),
            .I(\CONTROL.programCounter_1_reto_11 ));
    InMux I__3542 (
            .O(N__29621),
            .I(N__29618));
    LocalMux I__3541 (
            .O(N__29618),
            .I(\CONTROL.dout_reto_11 ));
    InMux I__3540 (
            .O(N__29615),
            .I(N__29612));
    LocalMux I__3539 (
            .O(N__29612),
            .I(N__29609));
    Span4Mux_h I__3538 (
            .O(N__29609),
            .I(N__29606));
    Odrv4 I__3537 (
            .O(N__29606),
            .I(\PROM.ROMDATA.m470_am ));
    InMux I__3536 (
            .O(N__29603),
            .I(N__29600));
    LocalMux I__3535 (
            .O(N__29600),
            .I(\CONTROL.dout_reto_14 ));
    InMux I__3534 (
            .O(N__29597),
            .I(N__29593));
    InMux I__3533 (
            .O(N__29596),
            .I(N__29590));
    LocalMux I__3532 (
            .O(N__29593),
            .I(N__29587));
    LocalMux I__3531 (
            .O(N__29590),
            .I(N__29584));
    Odrv4 I__3530 (
            .O(N__29587),
            .I(controlWord_18));
    Odrv4 I__3529 (
            .O(N__29584),
            .I(controlWord_18));
    CascadeMux I__3528 (
            .O(N__29579),
            .I(controlWord_18_cascade_));
    IoInMux I__3527 (
            .O(N__29576),
            .I(N__29573));
    LocalMux I__3526 (
            .O(N__29573),
            .I(N__29570));
    IoSpan4Mux I__3525 (
            .O(N__29570),
            .I(N__29567));
    Span4Mux_s0_h I__3524 (
            .O(N__29567),
            .I(N__29564));
    Sp12to4 I__3523 (
            .O(N__29564),
            .I(N__29561));
    Span12Mux_s8_h I__3522 (
            .O(N__29561),
            .I(N__29558));
    Span12Mux_h I__3521 (
            .O(N__29558),
            .I(N__29554));
    InMux I__3520 (
            .O(N__29557),
            .I(N__29551));
    Odrv12 I__3519 (
            .O(N__29554),
            .I(A2_c));
    LocalMux I__3518 (
            .O(N__29551),
            .I(A2_c));
    CascadeMux I__3517 (
            .O(N__29546),
            .I(\CONTROL.g0_3_i_1_0_cascade_ ));
    CascadeMux I__3516 (
            .O(N__29543),
            .I(\CONTROL.N_4_1_cascade_ ));
    CascadeMux I__3515 (
            .O(N__29540),
            .I(N__29536));
    CascadeMux I__3514 (
            .O(N__29539),
            .I(N__29533));
    InMux I__3513 (
            .O(N__29536),
            .I(N__29528));
    InMux I__3512 (
            .O(N__29533),
            .I(N__29528));
    LocalMux I__3511 (
            .O(N__29528),
            .I(N__29525));
    Span4Mux_v I__3510 (
            .O(N__29525),
            .I(N__29522));
    Span4Mux_h I__3509 (
            .O(N__29522),
            .I(N__29519));
    Odrv4 I__3508 (
            .O(N__29519),
            .I(\CONTROL.N_81_0 ));
    InMux I__3507 (
            .O(N__29516),
            .I(N__29513));
    LocalMux I__3506 (
            .O(N__29513),
            .I(\CONTROL.g0_3_i_a7_2_0 ));
    InMux I__3505 (
            .O(N__29510),
            .I(N__29507));
    LocalMux I__3504 (
            .O(N__29507),
            .I(\CONTROL.N_429 ));
    InMux I__3503 (
            .O(N__29504),
            .I(N__29501));
    LocalMux I__3502 (
            .O(N__29501),
            .I(\CONTROL.dout_reto_8 ));
    CascadeMux I__3501 (
            .O(N__29498),
            .I(\CONTROL.gpuWrite_RNOZ0Z_2_cascade_ ));
    CascadeMux I__3500 (
            .O(N__29495),
            .I(\CONTROL.busState96_cascade_ ));
    InMux I__3499 (
            .O(N__29492),
            .I(N__29489));
    LocalMux I__3498 (
            .O(N__29489),
            .I(\CONTROL.busState96 ));
    InMux I__3497 (
            .O(N__29486),
            .I(N__29483));
    LocalMux I__3496 (
            .O(N__29483),
            .I(\CONTROL.N_66_0 ));
    InMux I__3495 (
            .O(N__29480),
            .I(N__29477));
    LocalMux I__3494 (
            .O(N__29477),
            .I(\CONTROL.gpuWrite_RNOZ0Z_0 ));
    InMux I__3493 (
            .O(N__29474),
            .I(N__29470));
    CascadeMux I__3492 (
            .O(N__29473),
            .I(N__29467));
    LocalMux I__3491 (
            .O(N__29470),
            .I(N__29464));
    InMux I__3490 (
            .O(N__29467),
            .I(N__29461));
    Odrv12 I__3489 (
            .O(N__29464),
            .I(gpuWrite));
    LocalMux I__3488 (
            .O(N__29461),
            .I(gpuWrite));
    CascadeMux I__3487 (
            .O(N__29456),
            .I(N__29452));
    InMux I__3486 (
            .O(N__29455),
            .I(N__29448));
    InMux I__3485 (
            .O(N__29452),
            .I(N__29445));
    CascadeMux I__3484 (
            .O(N__29451),
            .I(N__29442));
    LocalMux I__3483 (
            .O(N__29448),
            .I(N__29439));
    LocalMux I__3482 (
            .O(N__29445),
            .I(N__29436));
    InMux I__3481 (
            .O(N__29442),
            .I(N__29433));
    Span4Mux_v I__3480 (
            .O(N__29439),
            .I(N__29430));
    Span4Mux_h I__3479 (
            .O(N__29436),
            .I(N__29425));
    LocalMux I__3478 (
            .O(N__29433),
            .I(N__29425));
    Span4Mux_h I__3477 (
            .O(N__29430),
            .I(N__29420));
    Span4Mux_v I__3476 (
            .O(N__29425),
            .I(N__29420));
    Odrv4 I__3475 (
            .O(N__29420),
            .I(controlWord_21));
    CascadeMux I__3474 (
            .O(N__29417),
            .I(\RAM.un1_WR_105_0Z0Z_3_cascade_ ));
    IoInMux I__3473 (
            .O(N__29414),
            .I(N__29411));
    LocalMux I__3472 (
            .O(N__29411),
            .I(N__29408));
    Span4Mux_s2_v I__3471 (
            .O(N__29408),
            .I(N__29405));
    Span4Mux_h I__3470 (
            .O(N__29405),
            .I(N__29402));
    Sp12to4 I__3469 (
            .O(N__29402),
            .I(N__29399));
    Span12Mux_h I__3468 (
            .O(N__29399),
            .I(N__29395));
    InMux I__3467 (
            .O(N__29398),
            .I(N__29392));
    Odrv12 I__3466 (
            .O(N__29395),
            .I(A5_c));
    LocalMux I__3465 (
            .O(N__29392),
            .I(A5_c));
    CascadeMux I__3464 (
            .O(N__29387),
            .I(N__29384));
    InMux I__3463 (
            .O(N__29384),
            .I(N__29381));
    LocalMux I__3462 (
            .O(N__29381),
            .I(N__29378));
    Span4Mux_v I__3461 (
            .O(N__29378),
            .I(N__29375));
    Span4Mux_h I__3460 (
            .O(N__29375),
            .I(N__29372));
    Odrv4 I__3459 (
            .O(N__29372),
            .I(\RAM.un1_WR_105_0Z0Z_11 ));
    InMux I__3458 (
            .O(N__29369),
            .I(N__29365));
    InMux I__3457 (
            .O(N__29368),
            .I(N__29362));
    LocalMux I__3456 (
            .O(N__29365),
            .I(N__29359));
    LocalMux I__3455 (
            .O(N__29362),
            .I(controlWord_23));
    Odrv4 I__3454 (
            .O(N__29359),
            .I(controlWord_23));
    IoInMux I__3453 (
            .O(N__29354),
            .I(N__29351));
    LocalMux I__3452 (
            .O(N__29351),
            .I(N__29348));
    Span12Mux_s8_h I__3451 (
            .O(N__29348),
            .I(N__29345));
    Span12Mux_h I__3450 (
            .O(N__29345),
            .I(N__29341));
    InMux I__3449 (
            .O(N__29344),
            .I(N__29338));
    Odrv12 I__3448 (
            .O(N__29341),
            .I(A7_c));
    LocalMux I__3447 (
            .O(N__29338),
            .I(A7_c));
    IoInMux I__3446 (
            .O(N__29333),
            .I(N__29330));
    LocalMux I__3445 (
            .O(N__29330),
            .I(N__29327));
    IoSpan4Mux I__3444 (
            .O(N__29327),
            .I(N__29324));
    Span4Mux_s3_h I__3443 (
            .O(N__29324),
            .I(N__29321));
    Sp12to4 I__3442 (
            .O(N__29321),
            .I(N__29318));
    Span12Mux_s11_h I__3441 (
            .O(N__29318),
            .I(N__29315));
    Odrv12 I__3440 (
            .O(N__29315),
            .I(gpuAddress_3));
    IoInMux I__3439 (
            .O(N__29312),
            .I(N__29309));
    LocalMux I__3438 (
            .O(N__29309),
            .I(N__29306));
    IoSpan4Mux I__3437 (
            .O(N__29306),
            .I(N__29303));
    Span4Mux_s0_h I__3436 (
            .O(N__29303),
            .I(N__29300));
    Sp12to4 I__3435 (
            .O(N__29300),
            .I(N__29297));
    Span12Mux_s11_h I__3434 (
            .O(N__29297),
            .I(N__29294));
    Span12Mux_v I__3433 (
            .O(N__29294),
            .I(N__29291));
    Odrv12 I__3432 (
            .O(N__29291),
            .I(gpuAddress_4));
    IoInMux I__3431 (
            .O(N__29288),
            .I(N__29285));
    LocalMux I__3430 (
            .O(N__29285),
            .I(N__29282));
    Span4Mux_s0_h I__3429 (
            .O(N__29282),
            .I(N__29279));
    Span4Mux_h I__3428 (
            .O(N__29279),
            .I(N__29276));
    Sp12to4 I__3427 (
            .O(N__29276),
            .I(N__29273));
    Span12Mux_v I__3426 (
            .O(N__29273),
            .I(N__29270));
    Odrv12 I__3425 (
            .O(N__29270),
            .I(gpuAddress_5));
    IoInMux I__3424 (
            .O(N__29267),
            .I(N__29264));
    LocalMux I__3423 (
            .O(N__29264),
            .I(N__29261));
    Span12Mux_s3_h I__3422 (
            .O(N__29261),
            .I(N__29258));
    Span12Mux_v I__3421 (
            .O(N__29258),
            .I(N__29255));
    Odrv12 I__3420 (
            .O(N__29255),
            .I(gpuAddress_6));
    IoInMux I__3419 (
            .O(N__29252),
            .I(N__29249));
    LocalMux I__3418 (
            .O(N__29249),
            .I(N__29246));
    Span12Mux_s2_h I__3417 (
            .O(N__29246),
            .I(N__29243));
    Span12Mux_h I__3416 (
            .O(N__29243),
            .I(N__29240));
    Span12Mux_v I__3415 (
            .O(N__29240),
            .I(N__29237));
    Odrv12 I__3414 (
            .O(N__29237),
            .I(gpuAddress_7));
    IoInMux I__3413 (
            .O(N__29234),
            .I(N__29231));
    LocalMux I__3412 (
            .O(N__29231),
            .I(N__29228));
    IoSpan4Mux I__3411 (
            .O(N__29228),
            .I(N__29225));
    Span4Mux_s2_h I__3410 (
            .O(N__29225),
            .I(N__29222));
    Span4Mux_v I__3409 (
            .O(N__29222),
            .I(N__29219));
    Span4Mux_v I__3408 (
            .O(N__29219),
            .I(N__29216));
    Span4Mux_h I__3407 (
            .O(N__29216),
            .I(N__29213));
    Span4Mux_h I__3406 (
            .O(N__29213),
            .I(N__29210));
    Odrv4 I__3405 (
            .O(N__29210),
            .I(gpuAddress_8));
    CascadeMux I__3404 (
            .O(N__29207),
            .I(\CONTROL.un1_busState119_1_i_0_1_cascade_ ));
    InMux I__3403 (
            .O(N__29204),
            .I(N__29201));
    LocalMux I__3402 (
            .O(N__29201),
            .I(N__29198));
    Span4Mux_v I__3401 (
            .O(N__29198),
            .I(N__29195));
    Span4Mux_v I__3400 (
            .O(N__29195),
            .I(N__29192));
    Span4Mux_v I__3399 (
            .O(N__29192),
            .I(N__29189));
    IoSpan4Mux I__3398 (
            .O(N__29189),
            .I(N__29186));
    Odrv4 I__3397 (
            .O(N__29186),
            .I(gpuOut_c_7));
    InMux I__3396 (
            .O(N__29183),
            .I(N__29180));
    LocalMux I__3395 (
            .O(N__29180),
            .I(N_168));
    CascadeMux I__3394 (
            .O(N__29177),
            .I(N_168_cascade_));
    CascadeMux I__3393 (
            .O(N__29174),
            .I(N__29170));
    InMux I__3392 (
            .O(N__29173),
            .I(N__29165));
    InMux I__3391 (
            .O(N__29170),
            .I(N__29165));
    LocalMux I__3390 (
            .O(N__29165),
            .I(N__29162));
    Span4Mux_v I__3389 (
            .O(N__29162),
            .I(N__29159));
    Span4Mux_v I__3388 (
            .O(N__29159),
            .I(N__29156));
    Span4Mux_v I__3387 (
            .O(N__29156),
            .I(N__29153));
    Span4Mux_v I__3386 (
            .O(N__29153),
            .I(N__29150));
    IoSpan4Mux I__3385 (
            .O(N__29150),
            .I(N__29147));
    Odrv4 I__3384 (
            .O(N__29147),
            .I(D7_in_c));
    CascadeMux I__3383 (
            .O(N__29144),
            .I(\CONTROL.bus_7_ns_1_7_cascade_ ));
    InMux I__3382 (
            .O(N__29141),
            .I(N__29135));
    InMux I__3381 (
            .O(N__29140),
            .I(N__29135));
    LocalMux I__3380 (
            .O(N__29135),
            .I(N__29132));
    Span4Mux_v I__3379 (
            .O(N__29132),
            .I(N__29129));
    Span4Mux_h I__3378 (
            .O(N__29129),
            .I(N__29126));
    Odrv4 I__3377 (
            .O(N__29126),
            .I(PROM_ROMDATA_dintern_23ro));
    CascadeMux I__3376 (
            .O(N__29123),
            .I(\CONTROL.bus_7_a1_1_8_cascade_ ));
    InMux I__3375 (
            .O(N__29120),
            .I(N__29117));
    LocalMux I__3374 (
            .O(N__29117),
            .I(N__29114));
    Span4Mux_v I__3373 (
            .O(N__29114),
            .I(N__29111));
    Odrv4 I__3372 (
            .O(N__29111),
            .I(\CONTROL.bus_sx_8 ));
    IoInMux I__3371 (
            .O(N__29108),
            .I(N__29105));
    LocalMux I__3370 (
            .O(N__29105),
            .I(N__29102));
    Span4Mux_s3_h I__3369 (
            .O(N__29102),
            .I(N__29099));
    Span4Mux_h I__3368 (
            .O(N__29099),
            .I(N__29096));
    Sp12to4 I__3367 (
            .O(N__29096),
            .I(N__29093));
    Span12Mux_v I__3366 (
            .O(N__29093),
            .I(N__29090));
    Odrv12 I__3365 (
            .O(N__29090),
            .I(gpuAddress_2));
    InMux I__3364 (
            .O(N__29087),
            .I(N__29084));
    LocalMux I__3363 (
            .O(N__29084),
            .I(\ALU.c_RNI3MHFZ0Z_11 ));
    InMux I__3362 (
            .O(N__29081),
            .I(N__29078));
    LocalMux I__3361 (
            .O(N__29078),
            .I(\ALU.dout_3_ns_1_11 ));
    CascadeMux I__3360 (
            .O(N__29075),
            .I(\ALU.dout_3_ns_1_10_cascade_ ));
    CascadeMux I__3359 (
            .O(N__29072),
            .I(\ALU.dout_6_ns_1_10_cascade_ ));
    CascadeMux I__3358 (
            .O(N__29069),
            .I(\ALU.N_1143_cascade_ ));
    InMux I__3357 (
            .O(N__29066),
            .I(N__29063));
    LocalMux I__3356 (
            .O(N__29063),
            .I(\ALU.N_1095 ));
    CascadeMux I__3355 (
            .O(N__29060),
            .I(aluOut_10_cascade_));
    InMux I__3354 (
            .O(N__29057),
            .I(N__29053));
    InMux I__3353 (
            .O(N__29056),
            .I(N__29050));
    LocalMux I__3352 (
            .O(N__29053),
            .I(N__29047));
    LocalMux I__3351 (
            .O(N__29050),
            .I(N__29044));
    Span4Mux_v I__3350 (
            .O(N__29047),
            .I(N__29041));
    Span4Mux_h I__3349 (
            .O(N__29044),
            .I(N__29038));
    Odrv4 I__3348 (
            .O(N__29041),
            .I(\CONTROL.bus_0_10 ));
    Odrv4 I__3347 (
            .O(N__29038),
            .I(\CONTROL.bus_0_10 ));
    InMux I__3346 (
            .O(N__29033),
            .I(N__29030));
    LocalMux I__3345 (
            .O(N__29030),
            .I(ALU_N_1141));
    InMux I__3344 (
            .O(N__29027),
            .I(N__29023));
    InMux I__3343 (
            .O(N__29026),
            .I(N__29020));
    LocalMux I__3342 (
            .O(N__29023),
            .I(ALU_N_1093));
    LocalMux I__3341 (
            .O(N__29020),
            .I(ALU_N_1093));
    InMux I__3340 (
            .O(N__29015),
            .I(N__29012));
    LocalMux I__3339 (
            .O(N__29012),
            .I(\ALU.N_1144 ));
    CascadeMux I__3338 (
            .O(N__29009),
            .I(\ALU.N_1096_cascade_ ));
    InMux I__3337 (
            .O(N__29006),
            .I(N__29003));
    LocalMux I__3336 (
            .O(N__29003),
            .I(N__29000));
    Span4Mux_h I__3335 (
            .O(N__29000),
            .I(N__28997));
    Odrv4 I__3334 (
            .O(N__28997),
            .I(DROM_ROMDATA_dintern_11ro));
    CascadeMux I__3333 (
            .O(N__28994),
            .I(aluOut_11_cascade_));
    CascadeMux I__3332 (
            .O(N__28991),
            .I(\ALU.operand2_7_ns_1_11_cascade_ ));
    InMux I__3331 (
            .O(N__28988),
            .I(N__28985));
    LocalMux I__3330 (
            .O(N__28985),
            .I(N__28982));
    Odrv4 I__3329 (
            .O(N__28982),
            .I(\ALU.b_RNI2TJC1Z0Z_11 ));
    CascadeMux I__3328 (
            .O(N__28979),
            .I(\ALU.operand2_11_cascade_ ));
    CascadeMux I__3327 (
            .O(N__28976),
            .I(\ALU.d_RNIMR627Z0Z_11_cascade_ ));
    CascadeMux I__3326 (
            .O(N__28973),
            .I(N__28970));
    InMux I__3325 (
            .O(N__28970),
            .I(N__28967));
    LocalMux I__3324 (
            .O(N__28967),
            .I(\ALU.a_RNIV5PUZ0Z_11 ));
    CascadeMux I__3323 (
            .O(N__28964),
            .I(N__28961));
    InMux I__3322 (
            .O(N__28961),
            .I(N__28958));
    LocalMux I__3321 (
            .O(N__28958),
            .I(N__28955));
    Odrv12 I__3320 (
            .O(N__28955),
            .I(\ALU.d_RNI9IN2HZ0Z_3 ));
    InMux I__3319 (
            .O(N__28952),
            .I(N__28949));
    LocalMux I__3318 (
            .O(N__28949),
            .I(N__28946));
    Span4Mux_v I__3317 (
            .O(N__28946),
            .I(N__28943));
    Odrv4 I__3316 (
            .O(N__28943),
            .I(\ALU.a_RNI2N741Z0Z_12 ));
    InMux I__3315 (
            .O(N__28940),
            .I(N__28937));
    LocalMux I__3314 (
            .O(N__28937),
            .I(N__28934));
    Span4Mux_v I__3313 (
            .O(N__28934),
            .I(N__28930));
    InMux I__3312 (
            .O(N__28933),
            .I(N__28927));
    Odrv4 I__3311 (
            .O(N__28930),
            .I(\ALU.d_RNIJRM75Z0Z_5 ));
    LocalMux I__3310 (
            .O(N__28927),
            .I(\ALU.d_RNIJRM75Z0Z_5 ));
    CascadeMux I__3309 (
            .O(N__28922),
            .I(N__28917));
    CascadeMux I__3308 (
            .O(N__28921),
            .I(N__28914));
    InMux I__3307 (
            .O(N__28920),
            .I(N__28911));
    InMux I__3306 (
            .O(N__28917),
            .I(N__28908));
    InMux I__3305 (
            .O(N__28914),
            .I(N__28905));
    LocalMux I__3304 (
            .O(N__28911),
            .I(N__28902));
    LocalMux I__3303 (
            .O(N__28908),
            .I(N__28899));
    LocalMux I__3302 (
            .O(N__28905),
            .I(N__28896));
    Span4Mux_h I__3301 (
            .O(N__28902),
            .I(N__28891));
    Span4Mux_h I__3300 (
            .O(N__28899),
            .I(N__28891));
    Span4Mux_h I__3299 (
            .O(N__28896),
            .I(N__28888));
    Span4Mux_v I__3298 (
            .O(N__28891),
            .I(N__28885));
    Span4Mux_v I__3297 (
            .O(N__28888),
            .I(N__28882));
    Odrv4 I__3296 (
            .O(N__28885),
            .I(DROM_ROMDATA_dintern_5ro));
    Odrv4 I__3295 (
            .O(N__28882),
            .I(DROM_ROMDATA_dintern_5ro));
    InMux I__3294 (
            .O(N__28877),
            .I(N__28873));
    InMux I__3293 (
            .O(N__28876),
            .I(N__28870));
    LocalMux I__3292 (
            .O(N__28873),
            .I(N__28867));
    LocalMux I__3291 (
            .O(N__28870),
            .I(N__28864));
    Odrv4 I__3290 (
            .O(N__28867),
            .I(\ALU.d_RNIC0VE6Z0Z_5 ));
    Odrv4 I__3289 (
            .O(N__28864),
            .I(\ALU.d_RNIC0VE6Z0Z_5 ));
    CascadeMux I__3288 (
            .O(N__28859),
            .I(N__28856));
    InMux I__3287 (
            .O(N__28856),
            .I(N__28853));
    LocalMux I__3286 (
            .O(N__28853),
            .I(N__28850));
    Odrv12 I__3285 (
            .O(N__28850),
            .I(\ALU.d_RNI693UNZ0Z_3 ));
    CascadeMux I__3284 (
            .O(N__28847),
            .I(N__28844));
    InMux I__3283 (
            .O(N__28844),
            .I(N__28841));
    LocalMux I__3282 (
            .O(N__28841),
            .I(N__28838));
    Odrv12 I__3281 (
            .O(N__28838),
            .I(\ALU.mult_95_c_RNOZ0Z_0 ));
    CascadeMux I__3280 (
            .O(N__28835),
            .I(\ALU.dout_6_ns_1_11_cascade_ ));
    InMux I__3279 (
            .O(N__28832),
            .I(\ALU.mult_3_c14 ));
    CascadeMux I__3278 (
            .O(N__28829),
            .I(N__28826));
    InMux I__3277 (
            .O(N__28826),
            .I(N__28823));
    LocalMux I__3276 (
            .O(N__28823),
            .I(\ALU.d_RNI2IA441Z0Z_2 ));
    CascadeMux I__3275 (
            .O(N__28820),
            .I(N__28817));
    InMux I__3274 (
            .O(N__28817),
            .I(N__28814));
    LocalMux I__3273 (
            .O(N__28814),
            .I(N__28811));
    Odrv4 I__3272 (
            .O(N__28811),
            .I(\ALU.d_RNI7SQI21Z0Z_2 ));
    CascadeMux I__3271 (
            .O(N__28808),
            .I(N__28805));
    InMux I__3270 (
            .O(N__28805),
            .I(N__28802));
    LocalMux I__3269 (
            .O(N__28802),
            .I(N__28799));
    Odrv12 I__3268 (
            .O(N__28799),
            .I(\ALU.d_RNID31VFZ0Z_3 ));
    InMux I__3267 (
            .O(N__28796),
            .I(N__28793));
    LocalMux I__3266 (
            .O(N__28793),
            .I(\ALU.d_RNIBRFE41Z0Z_2 ));
    InMux I__3265 (
            .O(N__28790),
            .I(N__28787));
    LocalMux I__3264 (
            .O(N__28787),
            .I(\ALU.d_RNI9DAEHZ0Z_3 ));
    CascadeMux I__3263 (
            .O(N__28784),
            .I(N__28781));
    InMux I__3262 (
            .O(N__28781),
            .I(N__28778));
    LocalMux I__3261 (
            .O(N__28778),
            .I(N__28775));
    Odrv4 I__3260 (
            .O(N__28775),
            .I(\ALU.d_RNI07V431Z0Z_2 ));
    InMux I__3259 (
            .O(N__28772),
            .I(\ALU.mult_3_c6 ));
    InMux I__3258 (
            .O(N__28769),
            .I(N__28766));
    LocalMux I__3257 (
            .O(N__28766),
            .I(\ALU.d_RNIJ0U031Z0Z_2 ));
    CascadeMux I__3256 (
            .O(N__28763),
            .I(N__28760));
    InMux I__3255 (
            .O(N__28760),
            .I(N__28757));
    LocalMux I__3254 (
            .O(N__28757),
            .I(\ALU.d_RNIV1LMHZ0Z_3 ));
    InMux I__3253 (
            .O(N__28754),
            .I(\ALU.mult_3_c7 ));
    InMux I__3252 (
            .O(N__28751),
            .I(N__28748));
    LocalMux I__3251 (
            .O(N__28748),
            .I(\ALU.d_RNIS69AHZ0Z_3 ));
    CascadeMux I__3250 (
            .O(N__28745),
            .I(N__28742));
    InMux I__3249 (
            .O(N__28742),
            .I(N__28739));
    LocalMux I__3248 (
            .O(N__28739),
            .I(\ALU.d_RNI12A911Z0Z_2 ));
    InMux I__3247 (
            .O(N__28736),
            .I(\ALU.mult_3_c8 ));
    InMux I__3246 (
            .O(N__28733),
            .I(N__28730));
    LocalMux I__3245 (
            .O(N__28730),
            .I(\ALU.d_RNINIF011Z0Z_2 ));
    InMux I__3244 (
            .O(N__28727),
            .I(\ALU.mult_3_c9 ));
    InMux I__3243 (
            .O(N__28724),
            .I(N__28721));
    LocalMux I__3242 (
            .O(N__28721),
            .I(N__28718));
    Odrv4 I__3241 (
            .O(N__28718),
            .I(\ALU.d_RNIINE1HZ0Z_3 ));
    InMux I__3240 (
            .O(N__28715),
            .I(bfn_12_12_0_));
    InMux I__3239 (
            .O(N__28712),
            .I(N__28709));
    LocalMux I__3238 (
            .O(N__28709),
            .I(N__28706));
    Span4Mux_h I__3237 (
            .O(N__28706),
            .I(N__28703));
    Odrv4 I__3236 (
            .O(N__28703),
            .I(\ALU.d_RNIMCVI41Z0Z_2 ));
    CascadeMux I__3235 (
            .O(N__28700),
            .I(N__28697));
    InMux I__3234 (
            .O(N__28697),
            .I(N__28694));
    LocalMux I__3233 (
            .O(N__28694),
            .I(N__28691));
    Span4Mux_v I__3232 (
            .O(N__28691),
            .I(N__28688));
    Odrv4 I__3231 (
            .O(N__28688),
            .I(\ALU.d_RNITCCHHZ0Z_3 ));
    InMux I__3230 (
            .O(N__28685),
            .I(\ALU.mult_3_c11 ));
    InMux I__3229 (
            .O(N__28682),
            .I(N__28679));
    LocalMux I__3228 (
            .O(N__28679),
            .I(N__28676));
    Span4Mux_h I__3227 (
            .O(N__28676),
            .I(N__28673));
    Span4Mux_h I__3226 (
            .O(N__28673),
            .I(N__28670));
    Odrv4 I__3225 (
            .O(N__28670),
            .I(\ALU.d_RNI18J1JZ0Z_3 ));
    InMux I__3224 (
            .O(N__28667),
            .I(\ALU.mult_3_c12 ));
    InMux I__3223 (
            .O(N__28664),
            .I(\ALU.mult_3_c13 ));
    CascadeMux I__3222 (
            .O(N__28661),
            .I(\ALU.status_19_2_cascade_ ));
    CascadeMux I__3221 (
            .O(N__28658),
            .I(N__28655));
    InMux I__3220 (
            .O(N__28655),
            .I(N__28652));
    LocalMux I__3219 (
            .O(N__28652),
            .I(N__28649));
    Span4Mux_h I__3218 (
            .O(N__28649),
            .I(N__28646));
    Span4Mux_v I__3217 (
            .O(N__28646),
            .I(N__28643));
    Odrv4 I__3216 (
            .O(N__28643),
            .I(romOut_4));
    InMux I__3215 (
            .O(N__28640),
            .I(N__28637));
    LocalMux I__3214 (
            .O(N__28637),
            .I(N__28634));
    Odrv4 I__3213 (
            .O(N__28634),
            .I(\CONTROL.busState_1_RNI7U266Z0Z_2 ));
    InMux I__3212 (
            .O(N__28631),
            .I(\ALU.mult_3_c3 ));
    CascadeMux I__3211 (
            .O(N__28628),
            .I(N__28625));
    InMux I__3210 (
            .O(N__28625),
            .I(N__28622));
    LocalMux I__3209 (
            .O(N__28622),
            .I(\ALU.d_RNITK2D51Z0Z_2 ));
    InMux I__3208 (
            .O(N__28619),
            .I(\ALU.mult_3_c4 ));
    InMux I__3207 (
            .O(N__28616),
            .I(N__28613));
    LocalMux I__3206 (
            .O(N__28613),
            .I(\ALU.d_RNIJBM6GZ0Z_3 ));
    CascadeMux I__3205 (
            .O(N__28610),
            .I(N__28607));
    InMux I__3204 (
            .O(N__28607),
            .I(N__28604));
    LocalMux I__3203 (
            .O(N__28604),
            .I(\ALU.d_RNIKG0L11Z0Z_2 ));
    InMux I__3202 (
            .O(N__28601),
            .I(\ALU.mult_3_c5 ));
    InMux I__3201 (
            .O(N__28598),
            .I(N__28595));
    LocalMux I__3200 (
            .O(N__28595),
            .I(N__28592));
    Span4Mux_v I__3199 (
            .O(N__28592),
            .I(N__28589));
    Odrv4 I__3198 (
            .O(N__28589),
            .I(\ALU.status_17_I_1_c_RNOZ0 ));
    CascadeMux I__3197 (
            .O(N__28586),
            .I(\ALU.N_834_cascade_ ));
    InMux I__3196 (
            .O(N__28583),
            .I(N__28580));
    LocalMux I__3195 (
            .O(N__28580),
            .I(N__28577));
    Span4Mux_v I__3194 (
            .O(N__28577),
            .I(N__28573));
    InMux I__3193 (
            .O(N__28576),
            .I(N__28570));
    Span4Mux_v I__3192 (
            .O(N__28573),
            .I(N__28567));
    LocalMux I__3191 (
            .O(N__28570),
            .I(busState_1_RNIDU0U1_2));
    Odrv4 I__3190 (
            .O(N__28567),
            .I(busState_1_RNIDU0U1_2));
    InMux I__3189 (
            .O(N__28562),
            .I(N__28559));
    LocalMux I__3188 (
            .O(N__28559),
            .I(\CONTROL.programCounter_1_reto_9 ));
    InMux I__3187 (
            .O(N__28556),
            .I(N__28553));
    LocalMux I__3186 (
            .O(N__28553),
            .I(\CONTROL.addrstack_reto_9 ));
    CascadeMux I__3185 (
            .O(N__28550),
            .I(\CONTROL.N_424_cascade_ ));
    InMux I__3184 (
            .O(N__28547),
            .I(N__28544));
    LocalMux I__3183 (
            .O(N__28544),
            .I(N__28541));
    Odrv12 I__3182 (
            .O(N__28541),
            .I(progRomAddress_9));
    InMux I__3181 (
            .O(N__28538),
            .I(N__28532));
    InMux I__3180 (
            .O(N__28537),
            .I(N__28532));
    LocalMux I__3179 (
            .O(N__28532),
            .I(CONTROL_addrstack_reto_8));
    InMux I__3178 (
            .O(N__28529),
            .I(N__28526));
    LocalMux I__3177 (
            .O(N__28526),
            .I(N_423));
    CascadeMux I__3176 (
            .O(N__28523),
            .I(progRomAddress_9_cascade_));
    InMux I__3175 (
            .O(N__28520),
            .I(N__28514));
    InMux I__3174 (
            .O(N__28519),
            .I(N__28514));
    LocalMux I__3173 (
            .O(N__28514),
            .I(N__28511));
    Span4Mux_v I__3172 (
            .O(N__28511),
            .I(N__28508));
    Odrv4 I__3171 (
            .O(N__28508),
            .I(\PROM.ROMDATA.dintern_adfltZ0Z_3 ));
    InMux I__3170 (
            .O(N__28505),
            .I(N__28502));
    LocalMux I__3169 (
            .O(N__28502),
            .I(N__28499));
    Odrv12 I__3168 (
            .O(N__28499),
            .I(\CONTROL.tempCounterZ0Z_10 ));
    InMux I__3167 (
            .O(N__28496),
            .I(N__28492));
    InMux I__3166 (
            .O(N__28495),
            .I(N__28489));
    LocalMux I__3165 (
            .O(N__28492),
            .I(N__28484));
    LocalMux I__3164 (
            .O(N__28489),
            .I(N__28484));
    Odrv12 I__3163 (
            .O(N__28484),
            .I(\CONTROL.programCounter_1_9 ));
    InMux I__3162 (
            .O(N__28481),
            .I(N__28478));
    LocalMux I__3161 (
            .O(N__28478),
            .I(N__28475));
    Odrv4 I__3160 (
            .O(N__28475),
            .I(\CONTROL.tempCounterZ0Z_9 ));
    CascadeMux I__3159 (
            .O(N__28472),
            .I(N__28469));
    InMux I__3158 (
            .O(N__28469),
            .I(N__28466));
    LocalMux I__3157 (
            .O(N__28466),
            .I(\ALU.rshift_3_ns_1_2 ));
    InMux I__3156 (
            .O(N__28463),
            .I(N__28460));
    LocalMux I__3155 (
            .O(N__28460),
            .I(N__28457));
    Span4Mux_v I__3154 (
            .O(N__28457),
            .I(N__28454));
    Span4Mux_h I__3153 (
            .O(N__28454),
            .I(N__28451));
    Odrv4 I__3152 (
            .O(N__28451),
            .I(\CONTROL.addrstack_13 ));
    InMux I__3151 (
            .O(N__28448),
            .I(N__28445));
    LocalMux I__3150 (
            .O(N__28445),
            .I(\CONTROL.addrstack_reto_13 ));
    InMux I__3149 (
            .O(N__28442),
            .I(N__28435));
    InMux I__3148 (
            .O(N__28441),
            .I(N__28435));
    InMux I__3147 (
            .O(N__28440),
            .I(N__28432));
    LocalMux I__3146 (
            .O(N__28435),
            .I(N__28429));
    LocalMux I__3145 (
            .O(N__28432),
            .I(progRomAddress_10));
    Odrv12 I__3144 (
            .O(N__28429),
            .I(progRomAddress_10));
    InMux I__3143 (
            .O(N__28424),
            .I(N__28421));
    LocalMux I__3142 (
            .O(N__28421),
            .I(\CONTROL.addrstack_reto_12 ));
    InMux I__3141 (
            .O(N__28418),
            .I(N__28414));
    InMux I__3140 (
            .O(N__28417),
            .I(N__28411));
    LocalMux I__3139 (
            .O(N__28414),
            .I(N__28408));
    LocalMux I__3138 (
            .O(N__28411),
            .I(progRomAddress_12));
    Odrv12 I__3137 (
            .O(N__28408),
            .I(progRomAddress_12));
    InMux I__3136 (
            .O(N__28403),
            .I(N__28400));
    LocalMux I__3135 (
            .O(N__28400),
            .I(N__28397));
    Span4Mux_h I__3134 (
            .O(N__28397),
            .I(N__28394));
    Odrv4 I__3133 (
            .O(N__28394),
            .I(\CONTROL.addrstack_10 ));
    InMux I__3132 (
            .O(N__28391),
            .I(N__28388));
    LocalMux I__3131 (
            .O(N__28388),
            .I(\CONTROL.addrstack_reto_10 ));
    InMux I__3130 (
            .O(N__28385),
            .I(N__28382));
    LocalMux I__3129 (
            .O(N__28382),
            .I(\CONTROL.programCounter_1_reto_8 ));
    CascadeMux I__3128 (
            .O(N__28379),
            .I(N_423_cascade_));
    InMux I__3127 (
            .O(N__28376),
            .I(N__28373));
    LocalMux I__3126 (
            .O(N__28373),
            .I(N__28370));
    Odrv4 I__3125 (
            .O(N__28370),
            .I(\CONTROL.programCounter_1_axb_8 ));
    CEMux I__3124 (
            .O(N__28367),
            .I(N__28364));
    LocalMux I__3123 (
            .O(N__28364),
            .I(N__28361));
    Span4Mux_v I__3122 (
            .O(N__28361),
            .I(N__28358));
    Odrv4 I__3121 (
            .O(N__28358),
            .I(\CONTROL.programCounter10 ));
    InMux I__3120 (
            .O(N__28355),
            .I(\CONTROL.programCounter_1_cry_11 ));
    InMux I__3119 (
            .O(N__28352),
            .I(\CONTROL.programCounter_1_cry_12 ));
    InMux I__3118 (
            .O(N__28349),
            .I(\CONTROL.programCounter_1_cry_13 ));
    InMux I__3117 (
            .O(N__28346),
            .I(\CONTROL.programCounter_1_cry_14 ));
    InMux I__3116 (
            .O(N__28343),
            .I(N__28339));
    InMux I__3115 (
            .O(N__28342),
            .I(N__28336));
    LocalMux I__3114 (
            .O(N__28339),
            .I(N__28333));
    LocalMux I__3113 (
            .O(N__28336),
            .I(N__28328));
    Span4Mux_h I__3112 (
            .O(N__28333),
            .I(N__28328));
    Odrv4 I__3111 (
            .O(N__28328),
            .I(\CONTROL.programCounter_1_13 ));
    InMux I__3110 (
            .O(N__28325),
            .I(N__28322));
    LocalMux I__3109 (
            .O(N__28322),
            .I(\CONTROL.programCounter_1_reto_13 ));
    InMux I__3108 (
            .O(N__28319),
            .I(N__28316));
    LocalMux I__3107 (
            .O(N__28316),
            .I(\CONTROL.dout_reto_13 ));
    CascadeMux I__3106 (
            .O(N__28313),
            .I(\CONTROL.N_428_cascade_ ));
    InMux I__3105 (
            .O(N__28310),
            .I(N__28306));
    InMux I__3104 (
            .O(N__28309),
            .I(N__28303));
    LocalMux I__3103 (
            .O(N__28306),
            .I(N__28300));
    LocalMux I__3102 (
            .O(N__28303),
            .I(progRomAddress_13));
    Odrv12 I__3101 (
            .O(N__28300),
            .I(progRomAddress_13));
    CascadeMux I__3100 (
            .O(N__28295),
            .I(N__28292));
    InMux I__3099 (
            .O(N__28292),
            .I(N__28289));
    LocalMux I__3098 (
            .O(N__28289),
            .I(\CONTROL.addrstack_reto_14 ));
    InMux I__3097 (
            .O(N__28286),
            .I(N__28282));
    InMux I__3096 (
            .O(N__28285),
            .I(N__28279));
    LocalMux I__3095 (
            .O(N__28282),
            .I(N__28276));
    LocalMux I__3094 (
            .O(N__28279),
            .I(progRomAddress_14));
    Odrv12 I__3093 (
            .O(N__28276),
            .I(progRomAddress_14));
    InMux I__3092 (
            .O(N__28271),
            .I(N__28268));
    LocalMux I__3091 (
            .O(N__28268),
            .I(N__28265));
    Span4Mux_v I__3090 (
            .O(N__28265),
            .I(N__28262));
    Odrv4 I__3089 (
            .O(N__28262),
            .I(\CONTROL.programCounter_1_axb_3 ));
    InMux I__3088 (
            .O(N__28259),
            .I(\CONTROL.programCounter_1_cry_2 ));
    InMux I__3087 (
            .O(N__28256),
            .I(\CONTROL.programCounter_1_cry_3 ));
    InMux I__3086 (
            .O(N__28253),
            .I(\CONTROL.programCounter_1_cry_4 ));
    InMux I__3085 (
            .O(N__28250),
            .I(\CONTROL.programCounter_1_cry_5 ));
    InMux I__3084 (
            .O(N__28247),
            .I(\CONTROL.programCounter_1_cry_6 ));
    InMux I__3083 (
            .O(N__28244),
            .I(bfn_11_22_0_));
    InMux I__3082 (
            .O(N__28241),
            .I(\CONTROL.programCounter_1_cry_8 ));
    InMux I__3081 (
            .O(N__28238),
            .I(\CONTROL.programCounter_1_cry_9 ));
    InMux I__3080 (
            .O(N__28235),
            .I(\CONTROL.programCounter_1_cry_10 ));
    CascadeMux I__3079 (
            .O(N__28232),
            .I(controlWord_29_cascade_));
    CascadeMux I__3078 (
            .O(N__28229),
            .I(N__28225));
    InMux I__3077 (
            .O(N__28228),
            .I(N__28222));
    InMux I__3076 (
            .O(N__28225),
            .I(N__28219));
    LocalMux I__3075 (
            .O(N__28222),
            .I(N__28216));
    LocalMux I__3074 (
            .O(N__28219),
            .I(N__28213));
    Odrv4 I__3073 (
            .O(N__28216),
            .I(controlWord_28));
    Odrv4 I__3072 (
            .O(N__28213),
            .I(controlWord_28));
    CascadeMux I__3071 (
            .O(N__28208),
            .I(controlWord_28_cascade_));
    IoInMux I__3070 (
            .O(N__28205),
            .I(N__28202));
    LocalMux I__3069 (
            .O(N__28202),
            .I(N__28199));
    IoSpan4Mux I__3068 (
            .O(N__28199),
            .I(N__28196));
    Span4Mux_s2_h I__3067 (
            .O(N__28196),
            .I(N__28193));
    Sp12to4 I__3066 (
            .O(N__28193),
            .I(N__28190));
    Span12Mux_h I__3065 (
            .O(N__28190),
            .I(N__28187));
    Span12Mux_v I__3064 (
            .O(N__28187),
            .I(N__28183));
    InMux I__3063 (
            .O(N__28186),
            .I(N__28180));
    Odrv12 I__3062 (
            .O(N__28183),
            .I(A12_c));
    LocalMux I__3061 (
            .O(N__28180),
            .I(A12_c));
    IoInMux I__3060 (
            .O(N__28175),
            .I(N__28172));
    LocalMux I__3059 (
            .O(N__28172),
            .I(N__28169));
    Span4Mux_s3_v I__3058 (
            .O(N__28169),
            .I(N__28166));
    Span4Mux_h I__3057 (
            .O(N__28166),
            .I(N__28163));
    Sp12to4 I__3056 (
            .O(N__28163),
            .I(N__28160));
    Span12Mux_h I__3055 (
            .O(N__28160),
            .I(N__28156));
    InMux I__3054 (
            .O(N__28159),
            .I(N__28153));
    Odrv12 I__3053 (
            .O(N__28156),
            .I(A13_c));
    LocalMux I__3052 (
            .O(N__28153),
            .I(A13_c));
    InMux I__3051 (
            .O(N__28148),
            .I(N__28145));
    LocalMux I__3050 (
            .O(N__28145),
            .I(N__28142));
    Span4Mux_v I__3049 (
            .O(N__28142),
            .I(N__28139));
    Odrv4 I__3048 (
            .O(N__28139),
            .I(\RAM.un1_WR_105_0Z0Z_10 ));
    InMux I__3047 (
            .O(N__28136),
            .I(\CONTROL.programCounter_1_cry_0 ));
    InMux I__3046 (
            .O(N__28133),
            .I(\CONTROL.programCounter_1_cry_1 ));
    CascadeMux I__3045 (
            .O(N__28130),
            .I(\CONTROL.busState_1_e_1_0_cascade_ ));
    CascadeMux I__3044 (
            .O(N__28127),
            .I(\CONTROL.un1_busState_1_sqmuxa_iZ0Z_0_cascade_ ));
    CEMux I__3043 (
            .O(N__28124),
            .I(N__28119));
    CEMux I__3042 (
            .O(N__28123),
            .I(N__28116));
    CEMux I__3041 (
            .O(N__28122),
            .I(N__28113));
    LocalMux I__3040 (
            .O(N__28119),
            .I(N__28105));
    LocalMux I__3039 (
            .O(N__28116),
            .I(N__28105));
    LocalMux I__3038 (
            .O(N__28113),
            .I(N__28102));
    CEMux I__3037 (
            .O(N__28112),
            .I(N__28099));
    CEMux I__3036 (
            .O(N__28111),
            .I(N__28096));
    CEMux I__3035 (
            .O(N__28110),
            .I(N__28093));
    Span4Mux_v I__3034 (
            .O(N__28105),
            .I(N__28086));
    Span4Mux_v I__3033 (
            .O(N__28102),
            .I(N__28086));
    LocalMux I__3032 (
            .O(N__28099),
            .I(N__28086));
    LocalMux I__3031 (
            .O(N__28096),
            .I(N_29));
    LocalMux I__3030 (
            .O(N__28093),
            .I(N_29));
    Odrv4 I__3029 (
            .O(N__28086),
            .I(N_29));
    InMux I__3028 (
            .O(N__28079),
            .I(N__28076));
    LocalMux I__3027 (
            .O(N__28076),
            .I(\CONTROL.N_352 ));
    InMux I__3026 (
            .O(N__28073),
            .I(N__28070));
    LocalMux I__3025 (
            .O(N__28070),
            .I(\CONTROL.un1_busState_1_sqmuxa_iZ0Z_0 ));
    InMux I__3024 (
            .O(N__28067),
            .I(N__28064));
    LocalMux I__3023 (
            .O(N__28064),
            .I(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_3 ));
    InMux I__3022 (
            .O(N__28061),
            .I(N__28058));
    LocalMux I__3021 (
            .O(N__28058),
            .I(N__28054));
    InMux I__3020 (
            .O(N__28057),
            .I(N__28051));
    Span4Mux_h I__3019 (
            .O(N__28054),
            .I(N__28048));
    LocalMux I__3018 (
            .O(N__28051),
            .I(N__28045));
    Odrv4 I__3017 (
            .O(N__28048),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_3 ));
    Odrv4 I__3016 (
            .O(N__28045),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_3 ));
    InMux I__3015 (
            .O(N__28040),
            .I(N__28037));
    LocalMux I__3014 (
            .O(N__28037),
            .I(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_0 ));
    InMux I__3013 (
            .O(N__28034),
            .I(N__28030));
    InMux I__3012 (
            .O(N__28033),
            .I(N__28027));
    LocalMux I__3011 (
            .O(N__28030),
            .I(N__28024));
    LocalMux I__3010 (
            .O(N__28027),
            .I(N__28021));
    Span4Mux_h I__3009 (
            .O(N__28024),
            .I(N__28018));
    Odrv4 I__3008 (
            .O(N__28021),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_0 ));
    Odrv4 I__3007 (
            .O(N__28018),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_0 ));
    InMux I__3006 (
            .O(N__28013),
            .I(N__28007));
    InMux I__3005 (
            .O(N__28012),
            .I(N__28007));
    LocalMux I__3004 (
            .O(N__28007),
            .I(N__28004));
    Span4Mux_h I__3003 (
            .O(N__28004),
            .I(N__28000));
    InMux I__3002 (
            .O(N__28003),
            .I(N__27997));
    Span4Mux_v I__3001 (
            .O(N__28000),
            .I(N__27994));
    LocalMux I__3000 (
            .O(N__27997),
            .I(DROM_ROMDATA_dintern_4ro));
    Odrv4 I__2999 (
            .O(N__27994),
            .I(DROM_ROMDATA_dintern_4ro));
    InMux I__2998 (
            .O(N__27989),
            .I(N__27985));
    InMux I__2997 (
            .O(N__27988),
            .I(N__27982));
    LocalMux I__2996 (
            .O(N__27985),
            .I(N__27979));
    LocalMux I__2995 (
            .O(N__27982),
            .I(N__27976));
    Odrv4 I__2994 (
            .O(N__27979),
            .I(controlWord_29));
    Odrv4 I__2993 (
            .O(N__27976),
            .I(controlWord_29));
    CascadeMux I__2992 (
            .O(N__27971),
            .I(\ALU.dout_3_ns_1_8_cascade_ ));
    InMux I__2991 (
            .O(N__27968),
            .I(N__27965));
    LocalMux I__2990 (
            .O(N__27965),
            .I(\ALU.c_RNIFT2SZ0Z_8 ));
    InMux I__2989 (
            .O(N__27962),
            .I(N__27959));
    LocalMux I__2988 (
            .O(N__27959),
            .I(N__27956));
    Span4Mux_h I__2987 (
            .O(N__27956),
            .I(N__27950));
    InMux I__2986 (
            .O(N__27955),
            .I(N__27943));
    InMux I__2985 (
            .O(N__27954),
            .I(N__27943));
    InMux I__2984 (
            .O(N__27953),
            .I(N__27943));
    Odrv4 I__2983 (
            .O(N__27950),
            .I(dataRomAddress_10));
    LocalMux I__2982 (
            .O(N__27943),
            .I(dataRomAddress_10));
    CascadeMux I__2981 (
            .O(N__27938),
            .I(N__27933));
    CascadeMux I__2980 (
            .O(N__27937),
            .I(N__27930));
    InMux I__2979 (
            .O(N__27936),
            .I(N__27927));
    InMux I__2978 (
            .O(N__27933),
            .I(N__27922));
    InMux I__2977 (
            .O(N__27930),
            .I(N__27922));
    LocalMux I__2976 (
            .O(N__27927),
            .I(dataRomAddress_12));
    LocalMux I__2975 (
            .O(N__27922),
            .I(dataRomAddress_12));
    CascadeMux I__2974 (
            .O(N__27917),
            .I(\PROM.ROMDATA.dintern_adfltZ0Z_4_cascade_ ));
    CascadeMux I__2973 (
            .O(N__27914),
            .I(\PROM.ROMDATA.dintern_12dflt_0Z0Z_1_cascade_ ));
    InMux I__2972 (
            .O(N__27911),
            .I(N__27908));
    LocalMux I__2971 (
            .O(N__27908),
            .I(\PROM.ROMDATA.dintern_adfltZ0Z_4 ));
    InMux I__2970 (
            .O(N__27905),
            .I(N__27902));
    LocalMux I__2969 (
            .O(N__27902),
            .I(N__27899));
    Span12Mux_v I__2968 (
            .O(N__27899),
            .I(N__27893));
    InMux I__2967 (
            .O(N__27898),
            .I(N__27890));
    InMux I__2966 (
            .O(N__27897),
            .I(N__27885));
    InMux I__2965 (
            .O(N__27896),
            .I(N__27885));
    Odrv12 I__2964 (
            .O(N__27893),
            .I(dataRomAddress_11));
    LocalMux I__2963 (
            .O(N__27890),
            .I(dataRomAddress_11));
    LocalMux I__2962 (
            .O(N__27885),
            .I(dataRomAddress_11));
    InMux I__2961 (
            .O(N__27878),
            .I(N__27875));
    LocalMux I__2960 (
            .O(N__27875),
            .I(\ALU.c_RNIAMVQZ0Z_6 ));
    InMux I__2959 (
            .O(N__27872),
            .I(N__27869));
    LocalMux I__2958 (
            .O(N__27869),
            .I(\ALU.d_RNIDV8EZ0Z_6 ));
    InMux I__2957 (
            .O(N__27866),
            .I(N__27863));
    LocalMux I__2956 (
            .O(N__27863),
            .I(\ALU.c_RNI230LZ0Z_10 ));
    CascadeMux I__2955 (
            .O(N__27860),
            .I(\ALU.a_RNIUI741Z0Z_10_cascade_ ));
    InMux I__2954 (
            .O(N__27857),
            .I(N__27854));
    LocalMux I__2953 (
            .O(N__27854),
            .I(\ALU.operand2_7_ns_1_10 ));
    CascadeMux I__2952 (
            .O(N__27851),
            .I(\ALU.dout_6_ns_1_8_cascade_ ));
    CascadeMux I__2951 (
            .O(N__27848),
            .I(ALU_N_1141_cascade_));
    CascadeMux I__2950 (
            .O(N__27845),
            .I(\CONTROL.bus_0_sx_8_cascade_ ));
    CascadeMux I__2949 (
            .O(N__27842),
            .I(N__27839));
    InMux I__2948 (
            .O(N__27839),
            .I(N__27836));
    LocalMux I__2947 (
            .O(N__27836),
            .I(N__27832));
    InMux I__2946 (
            .O(N__27835),
            .I(N__27829));
    Odrv4 I__2945 (
            .O(N__27832),
            .I(CONTROL_bus_0_8));
    LocalMux I__2944 (
            .O(N__27829),
            .I(CONTROL_bus_0_8));
    CascadeMux I__2943 (
            .O(N__27824),
            .I(\ALU.status_19_8_cascade_ ));
    CascadeMux I__2942 (
            .O(N__27821),
            .I(\ALU.operand2_7_ns_1_6_cascade_ ));
    InMux I__2941 (
            .O(N__27818),
            .I(N__27815));
    LocalMux I__2940 (
            .O(N__27815),
            .I(\ALU.operand2_6 ));
    InMux I__2939 (
            .O(N__27812),
            .I(N__27809));
    LocalMux I__2938 (
            .O(N__27809),
            .I(\ALU.b_RNI9JSPZ0Z_6 ));
    InMux I__2937 (
            .O(N__27806),
            .I(N__27803));
    LocalMux I__2936 (
            .O(N__27803),
            .I(\ALU.e_RNI6AJMZ0Z_6 ));
    CascadeMux I__2935 (
            .O(N__27800),
            .I(\ALU.operand2_7_ns_1_4_cascade_ ));
    InMux I__2934 (
            .O(N__27797),
            .I(N__27794));
    LocalMux I__2933 (
            .O(N__27794),
            .I(\ALU.operand2_4 ));
    InMux I__2932 (
            .O(N__27791),
            .I(N__27788));
    LocalMux I__2931 (
            .O(N__27788),
            .I(\ALU.c_RNI6IVQZ0Z_4 ));
    CascadeMux I__2930 (
            .O(N__27785),
            .I(\ALU.dout_6_ns_1_4_cascade_ ));
    InMux I__2929 (
            .O(N__27782),
            .I(N__27778));
    InMux I__2928 (
            .O(N__27781),
            .I(N__27775));
    LocalMux I__2927 (
            .O(N__27778),
            .I(\ALU.aZ0Z_4 ));
    LocalMux I__2926 (
            .O(N__27775),
            .I(\ALU.aZ0Z_4 ));
    CascadeMux I__2925 (
            .O(N__27770),
            .I(\ALU.dout_3_ns_1_4_cascade_ ));
    CascadeMux I__2924 (
            .O(N__27767),
            .I(\ALU.N_1089_cascade_ ));
    InMux I__2923 (
            .O(N__27764),
            .I(N__27761));
    LocalMux I__2922 (
            .O(N__27761),
            .I(\ALU.N_1137 ));
    CascadeMux I__2921 (
            .O(N__27758),
            .I(aluOut_4_cascade_));
    InMux I__2920 (
            .O(N__27755),
            .I(N__27749));
    InMux I__2919 (
            .O(N__27754),
            .I(N__27749));
    LocalMux I__2918 (
            .O(N__27749),
            .I(\ALU.d_RNIBJM75Z0Z_4 ));
    CascadeMux I__2917 (
            .O(N__27746),
            .I(\ALU.addsub_cry_3_c_RNIGCKVJZ0Z5_cascade_ ));
    CascadeMux I__2916 (
            .O(N__27743),
            .I(\ALU.addsub_cry_3_c_RNIM4CUTZ0Z9_cascade_ ));
    CascadeMux I__2915 (
            .O(N__27740),
            .I(\ALU.e_RNI26JMZ0Z_4_cascade_ ));
    InMux I__2914 (
            .O(N__27737),
            .I(N__27734));
    LocalMux I__2913 (
            .O(N__27734),
            .I(N__27731));
    Span4Mux_h I__2912 (
            .O(N__27731),
            .I(N__27728));
    Odrv4 I__2911 (
            .O(N__27728),
            .I(\CONTROL.tempCounterZ0Z_11 ));
    InMux I__2910 (
            .O(N__27725),
            .I(N__27722));
    LocalMux I__2909 (
            .O(N__27722),
            .I(N__27719));
    Span4Mux_v I__2908 (
            .O(N__27719),
            .I(N__27716));
    Odrv4 I__2907 (
            .O(N__27716),
            .I(\CONTROL.tempCounterZ0Z_15 ));
    InMux I__2906 (
            .O(N__27713),
            .I(N__27710));
    LocalMux I__2905 (
            .O(N__27710),
            .I(N__27707));
    Span4Mux_v I__2904 (
            .O(N__27707),
            .I(N__27704));
    Odrv4 I__2903 (
            .O(N__27704),
            .I(\CONTROL.tempCounterZ0Z_14 ));
    InMux I__2902 (
            .O(N__27701),
            .I(N__27698));
    LocalMux I__2901 (
            .O(N__27698),
            .I(N__27695));
    Odrv4 I__2900 (
            .O(N__27695),
            .I(\CONTROL.addrstack_8 ));
    InMux I__2899 (
            .O(N__27692),
            .I(N__27689));
    LocalMux I__2898 (
            .O(N__27689),
            .I(N__27686));
    Odrv4 I__2897 (
            .O(N__27686),
            .I(\CONTROL.addrstack_9 ));
    CascadeMux I__2896 (
            .O(N__27683),
            .I(N__27680));
    InMux I__2895 (
            .O(N__27680),
            .I(N__27677));
    LocalMux I__2894 (
            .O(N__27677),
            .I(N__27674));
    Odrv4 I__2893 (
            .O(N__27674),
            .I(\ALU.status_17_I_9_c_RNOZ0 ));
    InMux I__2892 (
            .O(N__27671),
            .I(N__27668));
    LocalMux I__2891 (
            .O(N__27668),
            .I(\CONTROL.g0_3_iZ0Z_1 ));
    InMux I__2890 (
            .O(N__27665),
            .I(N__27662));
    LocalMux I__2889 (
            .O(N__27662),
            .I(\CONTROL.g0_3_i_a7Z0Z_2 ));
    CascadeMux I__2888 (
            .O(N__27659),
            .I(N__27656));
    InMux I__2887 (
            .O(N__27656),
            .I(N__27653));
    LocalMux I__2886 (
            .O(N__27653),
            .I(N__27650));
    Odrv4 I__2885 (
            .O(N__27650),
            .I(\CONTROL.g0_0_2 ));
    InMux I__2884 (
            .O(N__27647),
            .I(N__27644));
    LocalMux I__2883 (
            .O(N__27644),
            .I(N__27641));
    Span4Mux_v I__2882 (
            .O(N__27641),
            .I(N__27638));
    Span4Mux_h I__2881 (
            .O(N__27638),
            .I(N__27635));
    Odrv4 I__2880 (
            .O(N__27635),
            .I(\CONTROL.addrstack_12 ));
    InMux I__2879 (
            .O(N__27632),
            .I(N__27629));
    LocalMux I__2878 (
            .O(N__27629),
            .I(N__27626));
    Span4Mux_h I__2877 (
            .O(N__27626),
            .I(N__27623));
    Odrv4 I__2876 (
            .O(N__27623),
            .I(\CONTROL.addrstack_11 ));
    InMux I__2875 (
            .O(N__27620),
            .I(N__27617));
    LocalMux I__2874 (
            .O(N__27617),
            .I(N__27614));
    Span4Mux_h I__2873 (
            .O(N__27614),
            .I(N__27611));
    Odrv4 I__2872 (
            .O(N__27611),
            .I(\CONTROL.addrstack_7 ));
    InMux I__2871 (
            .O(N__27608),
            .I(N__27605));
    LocalMux I__2870 (
            .O(N__27605),
            .I(N__27602));
    Span4Mux_h I__2869 (
            .O(N__27602),
            .I(N__27599));
    Odrv4 I__2868 (
            .O(N__27599),
            .I(\CONTROL.addrstack_14 ));
    InMux I__2867 (
            .O(N__27596),
            .I(N__27593));
    LocalMux I__2866 (
            .O(N__27593),
            .I(N__27590));
    Span4Mux_v I__2865 (
            .O(N__27590),
            .I(N__27587));
    Span4Mux_v I__2864 (
            .O(N__27587),
            .I(N__27584));
    Span4Mux_v I__2863 (
            .O(N__27584),
            .I(N__27581));
    Sp12to4 I__2862 (
            .O(N__27581),
            .I(N__27578));
    Odrv12 I__2861 (
            .O(N__27578),
            .I(D6_in_c));
    CascadeMux I__2860 (
            .O(N__27575),
            .I(\CONTROL.N_167_cascade_ ));
    InMux I__2859 (
            .O(N__27572),
            .I(N__27568));
    InMux I__2858 (
            .O(N__27571),
            .I(N__27565));
    LocalMux I__2857 (
            .O(N__27568),
            .I(N__27562));
    LocalMux I__2856 (
            .O(N__27565),
            .I(N_183));
    Odrv12 I__2855 (
            .O(N__27562),
            .I(N_183));
    CascadeMux I__2854 (
            .O(N__27557),
            .I(\CONTROL.addrstackptr_N_8_mux_1_0_cascade_ ));
    CascadeMux I__2853 (
            .O(N__27554),
            .I(N__27551));
    InMux I__2852 (
            .O(N__27551),
            .I(N__27548));
    LocalMux I__2851 (
            .O(N__27548),
            .I(N__27545));
    Span4Mux_v I__2850 (
            .O(N__27545),
            .I(N__27542));
    Odrv4 I__2849 (
            .O(N__27542),
            .I(\CONTROL.addrstackptr_N_6_0_1_i ));
    CascadeMux I__2848 (
            .O(N__27539),
            .I(\CONTROL.g0_3_i_2_cascade_ ));
    InMux I__2847 (
            .O(N__27536),
            .I(N__27533));
    LocalMux I__2846 (
            .O(N__27533),
            .I(\CONTROL.N_4_0 ));
    InMux I__2845 (
            .O(N__27530),
            .I(N__27523));
    InMux I__2844 (
            .O(N__27529),
            .I(N__27523));
    CascadeMux I__2843 (
            .O(N__27528),
            .I(N__27520));
    LocalMux I__2842 (
            .O(N__27523),
            .I(N__27517));
    InMux I__2841 (
            .O(N__27520),
            .I(N__27514));
    Odrv4 I__2840 (
            .O(N__27517),
            .I(\CONTROL.addrstack_1_5 ));
    LocalMux I__2839 (
            .O(N__27514),
            .I(\CONTROL.addrstack_1_5 ));
    CascadeMux I__2838 (
            .O(N__27509),
            .I(\CONTROL.N_4_0_cascade_ ));
    InMux I__2837 (
            .O(N__27506),
            .I(N__27503));
    LocalMux I__2836 (
            .O(N__27503),
            .I(\CONTROL.addrstackptr_N_8_mux_1_0 ));
    InMux I__2835 (
            .O(N__27500),
            .I(N__27495));
    InMux I__2834 (
            .O(N__27499),
            .I(N__27488));
    InMux I__2833 (
            .O(N__27498),
            .I(N__27488));
    LocalMux I__2832 (
            .O(N__27495),
            .I(N__27485));
    InMux I__2831 (
            .O(N__27494),
            .I(N__27480));
    InMux I__2830 (
            .O(N__27493),
            .I(N__27480));
    LocalMux I__2829 (
            .O(N__27488),
            .I(N__27477));
    Span4Mux_h I__2828 (
            .O(N__27485),
            .I(N__27474));
    LocalMux I__2827 (
            .O(N__27480),
            .I(\CONTROL.addrstackptrZ0Z_5 ));
    Odrv4 I__2826 (
            .O(N__27477),
            .I(\CONTROL.addrstackptrZ0Z_5 ));
    Odrv4 I__2825 (
            .O(N__27474),
            .I(\CONTROL.addrstackptrZ0Z_5 ));
    InMux I__2824 (
            .O(N__27467),
            .I(N__27463));
    InMux I__2823 (
            .O(N__27466),
            .I(N__27460));
    LocalMux I__2822 (
            .O(N__27463),
            .I(N__27457));
    LocalMux I__2821 (
            .O(N__27460),
            .I(N__27454));
    Span4Mux_v I__2820 (
            .O(N__27457),
            .I(N__27451));
    Span4Mux_h I__2819 (
            .O(N__27454),
            .I(N__27448));
    Odrv4 I__2818 (
            .O(N__27451),
            .I(\DROM.ROMDATA.dintern_0_2_NEW_1 ));
    Odrv4 I__2817 (
            .O(N__27448),
            .I(\DROM.ROMDATA.dintern_0_2_NEW_1 ));
    InMux I__2816 (
            .O(N__27443),
            .I(N__27440));
    LocalMux I__2815 (
            .O(N__27440),
            .I(N__27437));
    Odrv4 I__2814 (
            .O(N__27437),
            .I(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_1 ));
    InMux I__2813 (
            .O(N__27434),
            .I(N__27430));
    InMux I__2812 (
            .O(N__27433),
            .I(N__27427));
    LocalMux I__2811 (
            .O(N__27430),
            .I(N__27424));
    LocalMux I__2810 (
            .O(N__27427),
            .I(N__27421));
    Span4Mux_h I__2809 (
            .O(N__27424),
            .I(N__27418));
    Span4Mux_h I__2808 (
            .O(N__27421),
            .I(N__27415));
    Odrv4 I__2807 (
            .O(N__27418),
            .I(\DROM.ROMDATA.dintern_0_2_NEW_2 ));
    Odrv4 I__2806 (
            .O(N__27415),
            .I(\DROM.ROMDATA.dintern_0_2_NEW_2 ));
    InMux I__2805 (
            .O(N__27410),
            .I(N__27407));
    LocalMux I__2804 (
            .O(N__27407),
            .I(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_2 ));
    InMux I__2803 (
            .O(N__27404),
            .I(N__27401));
    LocalMux I__2802 (
            .O(N__27401),
            .I(N__27397));
    InMux I__2801 (
            .O(N__27400),
            .I(N__27394));
    Span4Mux_h I__2800 (
            .O(N__27397),
            .I(N__27391));
    LocalMux I__2799 (
            .O(N__27394),
            .I(N__27388));
    Odrv4 I__2798 (
            .O(N__27391),
            .I(\DROM.ROMDATA.dintern_0_2_NEW_3 ));
    Odrv4 I__2797 (
            .O(N__27388),
            .I(\DROM.ROMDATA.dintern_0_2_NEW_3 ));
    InMux I__2796 (
            .O(N__27383),
            .I(N__27380));
    LocalMux I__2795 (
            .O(N__27380),
            .I(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_3 ));
    InMux I__2794 (
            .O(N__27377),
            .I(N__27373));
    InMux I__2793 (
            .O(N__27376),
            .I(N__27370));
    LocalMux I__2792 (
            .O(N__27373),
            .I(N__27367));
    LocalMux I__2791 (
            .O(N__27370),
            .I(N__27364));
    Span12Mux_v I__2790 (
            .O(N__27367),
            .I(N__27361));
    Span4Mux_v I__2789 (
            .O(N__27364),
            .I(N__27358));
    Odrv12 I__2788 (
            .O(N__27361),
            .I(\DROM.ROMDATA.dintern_0_3_NEW_0 ));
    Odrv4 I__2787 (
            .O(N__27358),
            .I(\DROM.ROMDATA.dintern_0_3_NEW_0 ));
    InMux I__2786 (
            .O(N__27353),
            .I(N__27350));
    LocalMux I__2785 (
            .O(N__27350),
            .I(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_0 ));
    CascadeMux I__2784 (
            .O(N__27347),
            .I(N__27342));
    CascadeMux I__2783 (
            .O(N__27346),
            .I(N__27339));
    InMux I__2782 (
            .O(N__27345),
            .I(N__27334));
    InMux I__2781 (
            .O(N__27342),
            .I(N__27334));
    InMux I__2780 (
            .O(N__27339),
            .I(N__27331));
    LocalMux I__2779 (
            .O(N__27334),
            .I(N__27328));
    LocalMux I__2778 (
            .O(N__27331),
            .I(N__27325));
    Span4Mux_h I__2777 (
            .O(N__27328),
            .I(N__27322));
    Span4Mux_v I__2776 (
            .O(N__27325),
            .I(N__27317));
    Span4Mux_v I__2775 (
            .O(N__27322),
            .I(N__27317));
    Odrv4 I__2774 (
            .O(N__27317),
            .I(DROM_ROMDATA_dintern_6ro));
    CascadeMux I__2773 (
            .O(N__27314),
            .I(\CONTROL.N_199_cascade_ ));
    InMux I__2772 (
            .O(N__27311),
            .I(N__27308));
    LocalMux I__2771 (
            .O(N__27308),
            .I(N__27305));
    Span4Mux_h I__2770 (
            .O(N__27305),
            .I(N__27302));
    Sp12to4 I__2769 (
            .O(N__27302),
            .I(N__27299));
    Span12Mux_v I__2768 (
            .O(N__27299),
            .I(N__27296));
    Odrv12 I__2767 (
            .O(N__27296),
            .I(gpuOut_c_6));
    CascadeMux I__2766 (
            .O(N__27293),
            .I(DROM_ROMDATA_dintern_13ro_cascade_));
    CascadeMux I__2765 (
            .O(N__27290),
            .I(N__27287));
    InMux I__2764 (
            .O(N__27287),
            .I(N__27278));
    InMux I__2763 (
            .O(N__27286),
            .I(N__27278));
    InMux I__2762 (
            .O(N__27285),
            .I(N__27271));
    InMux I__2761 (
            .O(N__27284),
            .I(N__27271));
    InMux I__2760 (
            .O(N__27283),
            .I(N__27271));
    LocalMux I__2759 (
            .O(N__27278),
            .I(N__27265));
    LocalMux I__2758 (
            .O(N__27271),
            .I(N__27262));
    InMux I__2757 (
            .O(N__27270),
            .I(N__27255));
    InMux I__2756 (
            .O(N__27269),
            .I(N__27255));
    InMux I__2755 (
            .O(N__27268),
            .I(N__27255));
    Odrv4 I__2754 (
            .O(N__27265),
            .I(\CONTROL.bus_7_a0_2_8 ));
    Odrv4 I__2753 (
            .O(N__27262),
            .I(\CONTROL.bus_7_a0_2_8 ));
    LocalMux I__2752 (
            .O(N__27255),
            .I(\CONTROL.bus_7_a0_2_8 ));
    InMux I__2751 (
            .O(N__27248),
            .I(N__27245));
    LocalMux I__2750 (
            .O(N__27245),
            .I(DROM_ROMDATA_dintern_13ro));
    IoInMux I__2749 (
            .O(N__27242),
            .I(N__27239));
    LocalMux I__2748 (
            .O(N__27239),
            .I(N__27236));
    IoSpan4Mux I__2747 (
            .O(N__27236),
            .I(N__27232));
    IoInMux I__2746 (
            .O(N__27235),
            .I(N__27229));
    Span4Mux_s0_h I__2745 (
            .O(N__27232),
            .I(N__27226));
    LocalMux I__2744 (
            .O(N__27229),
            .I(N__27223));
    Span4Mux_h I__2743 (
            .O(N__27226),
            .I(N__27220));
    IoSpan4Mux I__2742 (
            .O(N__27223),
            .I(N__27217));
    Span4Mux_h I__2741 (
            .O(N__27220),
            .I(N__27214));
    IoSpan4Mux I__2740 (
            .O(N__27217),
            .I(N__27211));
    Sp12to4 I__2739 (
            .O(N__27214),
            .I(N__27208));
    Span4Mux_s2_h I__2738 (
            .O(N__27211),
            .I(N__27205));
    Span12Mux_h I__2737 (
            .O(N__27208),
            .I(N__27202));
    Span4Mux_h I__2736 (
            .O(N__27205),
            .I(N__27199));
    Odrv12 I__2735 (
            .O(N__27202),
            .I(bus_13));
    Odrv4 I__2734 (
            .O(N__27199),
            .I(bus_13));
    InMux I__2733 (
            .O(N__27194),
            .I(N__27190));
    InMux I__2732 (
            .O(N__27193),
            .I(N__27187));
    LocalMux I__2731 (
            .O(N__27190),
            .I(N__27184));
    LocalMux I__2730 (
            .O(N__27187),
            .I(DROM_ROMDATA_dintern_10ro));
    Odrv4 I__2729 (
            .O(N__27184),
            .I(DROM_ROMDATA_dintern_10ro));
    InMux I__2728 (
            .O(N__27179),
            .I(N__27175));
    InMux I__2727 (
            .O(N__27178),
            .I(N__27172));
    LocalMux I__2726 (
            .O(N__27175),
            .I(N__27169));
    LocalMux I__2725 (
            .O(N__27172),
            .I(N__27166));
    Span4Mux_h I__2724 (
            .O(N__27169),
            .I(N__27163));
    Span4Mux_h I__2723 (
            .O(N__27166),
            .I(N__27160));
    Odrv4 I__2722 (
            .O(N__27163),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_1 ));
    Odrv4 I__2721 (
            .O(N__27160),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_1 ));
    InMux I__2720 (
            .O(N__27155),
            .I(N__27152));
    LocalMux I__2719 (
            .O(N__27152),
            .I(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_1 ));
    InMux I__2718 (
            .O(N__27149),
            .I(N__27146));
    LocalMux I__2717 (
            .O(N__27146),
            .I(N__27142));
    InMux I__2716 (
            .O(N__27145),
            .I(N__27139));
    Span4Mux_h I__2715 (
            .O(N__27142),
            .I(N__27136));
    LocalMux I__2714 (
            .O(N__27139),
            .I(N__27133));
    Odrv4 I__2713 (
            .O(N__27136),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_2 ));
    Odrv4 I__2712 (
            .O(N__27133),
            .I(\DROM.ROMDATA.dintern_0_1_NEW_2 ));
    InMux I__2711 (
            .O(N__27128),
            .I(N__27125));
    LocalMux I__2710 (
            .O(N__27125),
            .I(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_2 ));
    CascadeMux I__2709 (
            .O(N__27122),
            .I(\DROM.ROMDATA.dintern_adfltZ0Z_3_cascade_ ));
    InMux I__2708 (
            .O(N__27119),
            .I(N__27116));
    LocalMux I__2707 (
            .O(N__27116),
            .I(\DROM.ROMDATA.dintern_adflt_sxZ0 ));
    InMux I__2706 (
            .O(N__27113),
            .I(N__27104));
    InMux I__2705 (
            .O(N__27112),
            .I(N__27104));
    InMux I__2704 (
            .O(N__27111),
            .I(N__27104));
    LocalMux I__2703 (
            .O(N__27104),
            .I(dataRomAddress_13));
    InMux I__2702 (
            .O(N__27101),
            .I(N__27092));
    InMux I__2701 (
            .O(N__27100),
            .I(N__27092));
    InMux I__2700 (
            .O(N__27099),
            .I(N__27092));
    LocalMux I__2699 (
            .O(N__27092),
            .I(dataRomAddress_14));
    CascadeMux I__2698 (
            .O(N__27089),
            .I(N__27084));
    InMux I__2697 (
            .O(N__27088),
            .I(N__27077));
    InMux I__2696 (
            .O(N__27087),
            .I(N__27077));
    InMux I__2695 (
            .O(N__27084),
            .I(N__27077));
    LocalMux I__2694 (
            .O(N__27077),
            .I(dataRomAddress_15));
    InMux I__2693 (
            .O(N__27074),
            .I(N__27071));
    LocalMux I__2692 (
            .O(N__27071),
            .I(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_1 ));
    InMux I__2691 (
            .O(N__27068),
            .I(N__27064));
    InMux I__2690 (
            .O(N__27067),
            .I(N__27061));
    LocalMux I__2689 (
            .O(N__27064),
            .I(N__27058));
    LocalMux I__2688 (
            .O(N__27061),
            .I(N__27055));
    Span4Mux_v I__2687 (
            .O(N__27058),
            .I(N__27050));
    Span4Mux_h I__2686 (
            .O(N__27055),
            .I(N__27050));
    Span4Mux_v I__2685 (
            .O(N__27050),
            .I(N__27047));
    Odrv4 I__2684 (
            .O(N__27047),
            .I(\DROM.ROMDATA.dintern_0_3_NEW_1 ));
    CascadeMux I__2683 (
            .O(N__27044),
            .I(N__27041));
    InMux I__2682 (
            .O(N__27041),
            .I(N__27038));
    LocalMux I__2681 (
            .O(N__27038),
            .I(N__27035));
    Sp12to4 I__2680 (
            .O(N__27035),
            .I(N__27032));
    Odrv12 I__2679 (
            .O(N__27032),
            .I(\ALU.status_18_cry_3_c_RNOZ0 ));
    CascadeMux I__2678 (
            .O(N__27029),
            .I(N_228_0_cascade_));
    InMux I__2677 (
            .O(N__27026),
            .I(N__27023));
    LocalMux I__2676 (
            .O(N__27023),
            .I(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_3 ));
    InMux I__2675 (
            .O(N__27020),
            .I(N__27014));
    InMux I__2674 (
            .O(N__27019),
            .I(N__27014));
    LocalMux I__2673 (
            .O(N__27014),
            .I(N__27011));
    Odrv4 I__2672 (
            .O(N__27011),
            .I(\DROM.ROMDATA.dintern_0_0_NEW_3 ));
    CascadeMux I__2671 (
            .O(N__27008),
            .I(DROM_ROMDATA_dintern_3ro_cascade_));
    InMux I__2670 (
            .O(N__27005),
            .I(N__27002));
    LocalMux I__2669 (
            .O(N__27002),
            .I(DROM_ROMDATA_dintern_1ro));
    CascadeMux I__2668 (
            .O(N__26999),
            .I(DROM_ROMDATA_dintern_adflt_cascade_));
    CascadeMux I__2667 (
            .O(N__26996),
            .I(N__26993));
    InMux I__2666 (
            .O(N__26993),
            .I(N__26990));
    LocalMux I__2665 (
            .O(N__26990),
            .I(N__26987));
    Span4Mux_v I__2664 (
            .O(N__26987),
            .I(N__26984));
    Odrv4 I__2663 (
            .O(N__26984),
            .I(\DROM.ROMDATA.dintern_adfltZ0Z_3 ));
    CascadeMux I__2662 (
            .O(N__26981),
            .I(\ALU.operand2_10_cascade_ ));
    CascadeMux I__2661 (
            .O(N__26978),
            .I(\ALU.status_19_9_cascade_ ));
    CascadeMux I__2660 (
            .O(N__26975),
            .I(\ALU.e_RNIBHMNZ0Z_8_cascade_ ));
    InMux I__2659 (
            .O(N__26972),
            .I(N__26969));
    LocalMux I__2658 (
            .O(N__26969),
            .I(\ALU.d_RNIIINJZ0Z_8 ));
    InMux I__2657 (
            .O(N__26966),
            .I(N__26963));
    LocalMux I__2656 (
            .O(N__26963),
            .I(\ALU.operand2_7_ns_1_8 ));
    CascadeMux I__2655 (
            .O(N__26960),
            .I(\ALU.b_RNIE6BVZ0Z_8_cascade_ ));
    InMux I__2654 (
            .O(N__26957),
            .I(N__26954));
    LocalMux I__2653 (
            .O(N__26954),
            .I(N__26951));
    Odrv12 I__2652 (
            .O(N__26951),
            .I(\ALU.operand2_8 ));
    InMux I__2651 (
            .O(N__26948),
            .I(N__26945));
    LocalMux I__2650 (
            .O(N__26945),
            .I(busState_1_RNI05PC2_0));
    CascadeMux I__2649 (
            .O(N__26942),
            .I(\ALU.operand2_8_cascade_ ));
    InMux I__2648 (
            .O(N__26939),
            .I(N__26936));
    LocalMux I__2647 (
            .O(N__26936),
            .I(N_182));
    InMux I__2646 (
            .O(N__26933),
            .I(N__26927));
    InMux I__2645 (
            .O(N__26932),
            .I(N__26927));
    LocalMux I__2644 (
            .O(N__26927),
            .I(N__26924));
    Odrv4 I__2643 (
            .O(N__26924),
            .I(\ALU.combOperand2_0_0_6 ));
    InMux I__2642 (
            .O(N__26921),
            .I(N__26918));
    LocalMux I__2641 (
            .O(N__26918),
            .I(\ALU.b_RNI4VJC1Z0Z_12 ));
    InMux I__2640 (
            .O(N__26915),
            .I(N__26912));
    LocalMux I__2639 (
            .O(N__26912),
            .I(\ALU.d_RNI4BCTZ0Z_10 ));
    CascadeMux I__2638 (
            .O(N__26909),
            .I(\ALU.b_RNI0RJC1Z0Z_10_cascade_ ));
    CascadeMux I__2637 (
            .O(N__26906),
            .I(N__26902));
    CascadeMux I__2636 (
            .O(N__26905),
            .I(N__26899));
    InMux I__2635 (
            .O(N__26902),
            .I(N__26896));
    InMux I__2634 (
            .O(N__26899),
            .I(N__26892));
    LocalMux I__2633 (
            .O(N__26896),
            .I(N__26889));
    InMux I__2632 (
            .O(N__26895),
            .I(N__26886));
    LocalMux I__2631 (
            .O(N__26892),
            .I(N__26883));
    Odrv4 I__2630 (
            .O(N__26889),
            .I(\ALU.operand2_10 ));
    LocalMux I__2629 (
            .O(N__26886),
            .I(\ALU.operand2_10 ));
    Odrv4 I__2628 (
            .O(N__26883),
            .I(\ALU.operand2_10 ));
    CascadeMux I__2627 (
            .O(N__26876),
            .I(\ALU.combOperand2_0_4_cascade_ ));
    CascadeMux I__2626 (
            .O(N__26873),
            .I(N_181_cascade_));
    InMux I__2625 (
            .O(N__26870),
            .I(N__26867));
    LocalMux I__2624 (
            .O(N__26867),
            .I(\ALU.d_RNIVKK66Z0Z_4 ));
    CascadeMux I__2623 (
            .O(N__26864),
            .I(\ALU.d_RNIVKK66Z0Z_4_cascade_ ));
    CascadeMux I__2622 (
            .O(N__26861),
            .I(N__26858));
    InMux I__2621 (
            .O(N__26858),
            .I(N__26854));
    CascadeMux I__2620 (
            .O(N__26857),
            .I(N__26851));
    LocalMux I__2619 (
            .O(N__26854),
            .I(N__26848));
    InMux I__2618 (
            .O(N__26851),
            .I(N__26845));
    Span4Mux_h I__2617 (
            .O(N__26848),
            .I(N__26841));
    LocalMux I__2616 (
            .O(N__26845),
            .I(N__26838));
    InMux I__2615 (
            .O(N__26844),
            .I(N__26835));
    Odrv4 I__2614 (
            .O(N__26841),
            .I(\ALU.combOperand2_0_4 ));
    Odrv4 I__2613 (
            .O(N__26838),
            .I(\ALU.combOperand2_0_4 ));
    LocalMux I__2612 (
            .O(N__26835),
            .I(\ALU.combOperand2_0_4 ));
    CascadeMux I__2611 (
            .O(N__26828),
            .I(N__26825));
    InMux I__2610 (
            .O(N__26825),
            .I(N__26822));
    LocalMux I__2609 (
            .O(N__26822),
            .I(N__26819));
    Sp12to4 I__2608 (
            .O(N__26819),
            .I(N__26816));
    Odrv12 I__2607 (
            .O(N__26816),
            .I(\ALU.status_17_I_33_c_RNOZ0 ));
    InMux I__2606 (
            .O(N__26813),
            .I(N__26809));
    InMux I__2605 (
            .O(N__26812),
            .I(N__26806));
    LocalMux I__2604 (
            .O(N__26809),
            .I(\ALU.combOperand2_0_6 ));
    LocalMux I__2603 (
            .O(N__26806),
            .I(\ALU.combOperand2_0_6 ));
    CascadeMux I__2602 (
            .O(N__26801),
            .I(\ALU.combOperand2_0_6_cascade_ ));
    CascadeMux I__2601 (
            .O(N__26798),
            .I(\ALU.status_19_5_cascade_ ));
    CascadeMux I__2600 (
            .O(N__26795),
            .I(\ALU.dout_6_ns_1_5_cascade_ ));
    CascadeMux I__2599 (
            .O(N__26792),
            .I(\ALU.N_1138_cascade_ ));
    InMux I__2598 (
            .O(N__26789),
            .I(N__26786));
    LocalMux I__2597 (
            .O(N__26786),
            .I(\ALU.N_1090 ));
    CascadeMux I__2596 (
            .O(N__26783),
            .I(aluOut_5_cascade_));
    CascadeMux I__2595 (
            .O(N__26780),
            .I(\ALU.status_19_4_cascade_ ));
    InMux I__2594 (
            .O(N__26777),
            .I(N__26774));
    LocalMux I__2593 (
            .O(N__26774),
            .I(N__26771));
    Odrv4 I__2592 (
            .O(N__26771),
            .I(\ALU.status_17_I_15_c_RNOZ0 ));
    InMux I__2591 (
            .O(N__26768),
            .I(\CONTROL.addrstack_1_cry_0 ));
    InMux I__2590 (
            .O(N__26765),
            .I(\CONTROL.addrstack_1_cry_1 ));
    InMux I__2589 (
            .O(N__26762),
            .I(\CONTROL.addrstack_1_cry_2 ));
    InMux I__2588 (
            .O(N__26759),
            .I(\CONTROL.addrstack_1_cry_3 ));
    InMux I__2587 (
            .O(N__26756),
            .I(\CONTROL.addrstack_1_cry_4 ));
    CascadeMux I__2586 (
            .O(N__26753),
            .I(N__26747));
    CascadeMux I__2585 (
            .O(N__26752),
            .I(N__26744));
    InMux I__2584 (
            .O(N__26751),
            .I(N__26737));
    InMux I__2583 (
            .O(N__26750),
            .I(N__26737));
    InMux I__2582 (
            .O(N__26747),
            .I(N__26737));
    InMux I__2581 (
            .O(N__26744),
            .I(N__26734));
    LocalMux I__2580 (
            .O(N__26737),
            .I(N__26729));
    LocalMux I__2579 (
            .O(N__26734),
            .I(N__26729));
    Odrv4 I__2578 (
            .O(N__26729),
            .I(\CONTROL.addrstackptrZ0Z_6 ));
    InMux I__2577 (
            .O(N__26726),
            .I(N__26719));
    InMux I__2576 (
            .O(N__26725),
            .I(N__26719));
    CascadeMux I__2575 (
            .O(N__26724),
            .I(N__26716));
    LocalMux I__2574 (
            .O(N__26719),
            .I(N__26713));
    InMux I__2573 (
            .O(N__26716),
            .I(N__26710));
    Odrv12 I__2572 (
            .O(N__26713),
            .I(\CONTROL.addrstack_1_6 ));
    LocalMux I__2571 (
            .O(N__26710),
            .I(\CONTROL.addrstack_1_6 ));
    InMux I__2570 (
            .O(N__26705),
            .I(\CONTROL.addrstack_1_cry_5 ));
    InMux I__2569 (
            .O(N__26702),
            .I(\CONTROL.addrstack_1_cry_6 ));
    CascadeMux I__2568 (
            .O(N__26699),
            .I(\ALU.dout_3_ns_1_5_cascade_ ));
    CascadeMux I__2567 (
            .O(N__26696),
            .I(\CONTROL.g0_3_cascade_ ));
    CascadeMux I__2566 (
            .O(N__26693),
            .I(\CONTROL.addrstackptr_N_10_mux_0_0_0_cascade_ ));
    CascadeMux I__2565 (
            .O(N__26690),
            .I(N__26687));
    InMux I__2564 (
            .O(N__26687),
            .I(N__26684));
    LocalMux I__2563 (
            .O(N__26684),
            .I(N__26681));
    Span4Mux_v I__2562 (
            .O(N__26681),
            .I(N__26678));
    Odrv4 I__2561 (
            .O(N__26678),
            .I(\CONTROL.addrstackptr_N_7_0_i ));
    CascadeMux I__2560 (
            .O(N__26675),
            .I(\CONTROL.N_6_1_cascade_ ));
    InMux I__2559 (
            .O(N__26672),
            .I(N__26669));
    LocalMux I__2558 (
            .O(N__26669),
            .I(\CONTROL.N_4_2 ));
    CascadeMux I__2557 (
            .O(N__26666),
            .I(\CONTROL.N_4_2_cascade_ ));
    InMux I__2556 (
            .O(N__26663),
            .I(N__26660));
    LocalMux I__2555 (
            .O(N__26660),
            .I(\CONTROL.addrstackptr_N_10_mux_0_0_0 ));
    InMux I__2554 (
            .O(N__26657),
            .I(N__26654));
    LocalMux I__2553 (
            .O(N__26654),
            .I(\CONTROL.tempCounterZ0Z_13 ));
    InMux I__2552 (
            .O(N__26651),
            .I(N__26648));
    LocalMux I__2551 (
            .O(N__26648),
            .I(N__26645));
    Odrv4 I__2550 (
            .O(N__26645),
            .I(\CONTROL.tempCounterZ0Z_6 ));
    CascadeMux I__2549 (
            .O(N__26642),
            .I(PROM_ROMDATA_dintern_23ro_cascade_));
    CascadeMux I__2548 (
            .O(N__26639),
            .I(N__26636));
    CascadeBuf I__2547 (
            .O(N__26636),
            .I(N__26633));
    CascadeMux I__2546 (
            .O(N__26633),
            .I(N__26630));
    CascadeBuf I__2545 (
            .O(N__26630),
            .I(N__26627));
    CascadeMux I__2544 (
            .O(N__26627),
            .I(N__26624));
    CascadeBuf I__2543 (
            .O(N__26624),
            .I(N__26621));
    CascadeMux I__2542 (
            .O(N__26621),
            .I(N__26618));
    InMux I__2541 (
            .O(N__26618),
            .I(N__26615));
    LocalMux I__2540 (
            .O(N__26615),
            .I(N__26612));
    Span4Mux_h I__2539 (
            .O(N__26612),
            .I(N__26609));
    Odrv4 I__2538 (
            .O(N__26609),
            .I(CONTROL_romAddReg_7_7));
    CascadeMux I__2537 (
            .O(N__26606),
            .I(N__26603));
    CascadeBuf I__2536 (
            .O(N__26603),
            .I(N__26600));
    CascadeMux I__2535 (
            .O(N__26600),
            .I(N__26597));
    CascadeBuf I__2534 (
            .O(N__26597),
            .I(N__26594));
    CascadeMux I__2533 (
            .O(N__26594),
            .I(N__26591));
    CascadeBuf I__2532 (
            .O(N__26591),
            .I(N__26588));
    CascadeMux I__2531 (
            .O(N__26588),
            .I(N__26585));
    InMux I__2530 (
            .O(N__26585),
            .I(N__26582));
    LocalMux I__2529 (
            .O(N__26582),
            .I(N__26579));
    Odrv4 I__2528 (
            .O(N__26579),
            .I(CONTROL_romAddReg_7_6));
    CascadeMux I__2527 (
            .O(N__26576),
            .I(\PROM.ROMDATA.m465_bm_cascade_ ));
    CascadeMux I__2526 (
            .O(N__26573),
            .I(\PROM.ROMDATA.m471_ns_1_cascade_ ));
    CascadeMux I__2525 (
            .O(N__26570),
            .I(\PROM.ROMDATA.m471_ns_cascade_ ));
    CascadeMux I__2524 (
            .O(N__26567),
            .I(controlWord_24_cascade_));
    CascadeMux I__2523 (
            .O(N__26564),
            .I(N__26561));
    CascadeBuf I__2522 (
            .O(N__26561),
            .I(N__26558));
    CascadeMux I__2521 (
            .O(N__26558),
            .I(N__26555));
    CascadeBuf I__2520 (
            .O(N__26555),
            .I(N__26552));
    CascadeMux I__2519 (
            .O(N__26552),
            .I(N__26549));
    CascadeBuf I__2518 (
            .O(N__26549),
            .I(N__26546));
    CascadeMux I__2517 (
            .O(N__26546),
            .I(N__26543));
    InMux I__2516 (
            .O(N__26543),
            .I(N__26540));
    LocalMux I__2515 (
            .O(N__26540),
            .I(CONTROL_romAddReg_7_8));
    CascadeMux I__2514 (
            .O(N__26537),
            .I(N__26534));
    CascadeBuf I__2513 (
            .O(N__26534),
            .I(N__26531));
    CascadeMux I__2512 (
            .O(N__26531),
            .I(N__26528));
    CascadeBuf I__2511 (
            .O(N__26528),
            .I(N__26525));
    CascadeMux I__2510 (
            .O(N__26525),
            .I(N__26522));
    CascadeBuf I__2509 (
            .O(N__26522),
            .I(N__26519));
    CascadeMux I__2508 (
            .O(N__26519),
            .I(N__26516));
    InMux I__2507 (
            .O(N__26516),
            .I(N__26513));
    LocalMux I__2506 (
            .O(N__26513),
            .I(CONTROL_romAddReg_7_4));
    IoInMux I__2505 (
            .O(N__26510),
            .I(N__26507));
    LocalMux I__2504 (
            .O(N__26507),
            .I(N__26504));
    Span4Mux_s1_h I__2503 (
            .O(N__26504),
            .I(N__26501));
    Span4Mux_v I__2502 (
            .O(N__26501),
            .I(N__26498));
    Span4Mux_h I__2501 (
            .O(N__26498),
            .I(N__26495));
    Odrv4 I__2500 (
            .O(N__26495),
            .I(gpuAddress_10));
    IoInMux I__2499 (
            .O(N__26492),
            .I(N__26489));
    LocalMux I__2498 (
            .O(N__26489),
            .I(N__26486));
    IoSpan4Mux I__2497 (
            .O(N__26486),
            .I(N__26483));
    IoSpan4Mux I__2496 (
            .O(N__26483),
            .I(N__26480));
    Sp12to4 I__2495 (
            .O(N__26480),
            .I(N__26477));
    Odrv12 I__2494 (
            .O(N__26477),
            .I(gpuAddress_12));
    IoInMux I__2493 (
            .O(N__26474),
            .I(N__26471));
    LocalMux I__2492 (
            .O(N__26471),
            .I(N__26468));
    IoSpan4Mux I__2491 (
            .O(N__26468),
            .I(N__26465));
    IoSpan4Mux I__2490 (
            .O(N__26465),
            .I(N__26462));
    Span4Mux_s1_h I__2489 (
            .O(N__26462),
            .I(N__26459));
    Span4Mux_h I__2488 (
            .O(N__26459),
            .I(N__26456));
    Odrv4 I__2487 (
            .O(N__26456),
            .I(gpuAddress_13));
    IoInMux I__2486 (
            .O(N__26453),
            .I(N__26450));
    LocalMux I__2485 (
            .O(N__26450),
            .I(N__26447));
    IoSpan4Mux I__2484 (
            .O(N__26447),
            .I(N__26444));
    IoSpan4Mux I__2483 (
            .O(N__26444),
            .I(N__26441));
    Span4Mux_s2_h I__2482 (
            .O(N__26441),
            .I(N__26438));
    Span4Mux_h I__2481 (
            .O(N__26438),
            .I(N__26435));
    Odrv4 I__2480 (
            .O(N__26435),
            .I(gpuAddress_15));
    CascadeMux I__2479 (
            .O(N__26432),
            .I(N__26429));
    CascadeBuf I__2478 (
            .O(N__26429),
            .I(N__26426));
    CascadeMux I__2477 (
            .O(N__26426),
            .I(N__26423));
    CascadeBuf I__2476 (
            .O(N__26423),
            .I(N__26420));
    CascadeMux I__2475 (
            .O(N__26420),
            .I(N__26417));
    CascadeBuf I__2474 (
            .O(N__26417),
            .I(N__26414));
    CascadeMux I__2473 (
            .O(N__26414),
            .I(N__26411));
    InMux I__2472 (
            .O(N__26411),
            .I(N__26408));
    LocalMux I__2471 (
            .O(N__26408),
            .I(N__26405));
    Span4Mux_h I__2470 (
            .O(N__26405),
            .I(N__26402));
    Odrv4 I__2469 (
            .O(N__26402),
            .I(CONTROL_romAddReg_7_2));
    CascadeMux I__2468 (
            .O(N__26399),
            .I(N__26396));
    CascadeBuf I__2467 (
            .O(N__26396),
            .I(N__26393));
    CascadeMux I__2466 (
            .O(N__26393),
            .I(N__26390));
    CascadeBuf I__2465 (
            .O(N__26390),
            .I(N__26387));
    CascadeMux I__2464 (
            .O(N__26387),
            .I(N__26384));
    CascadeBuf I__2463 (
            .O(N__26384),
            .I(N__26381));
    CascadeMux I__2462 (
            .O(N__26381),
            .I(N__26378));
    InMux I__2461 (
            .O(N__26378),
            .I(N__26375));
    LocalMux I__2460 (
            .O(N__26375),
            .I(N__26372));
    Odrv4 I__2459 (
            .O(N__26372),
            .I(CONTROL_romAddReg_7_3));
    CascadeMux I__2458 (
            .O(N__26369),
            .I(N__26366));
    CascadeBuf I__2457 (
            .O(N__26366),
            .I(N__26363));
    CascadeMux I__2456 (
            .O(N__26363),
            .I(N__26360));
    CascadeBuf I__2455 (
            .O(N__26360),
            .I(N__26357));
    CascadeMux I__2454 (
            .O(N__26357),
            .I(N__26354));
    CascadeBuf I__2453 (
            .O(N__26354),
            .I(N__26351));
    CascadeMux I__2452 (
            .O(N__26351),
            .I(N__26348));
    InMux I__2451 (
            .O(N__26348),
            .I(N__26345));
    LocalMux I__2450 (
            .O(N__26345),
            .I(N__26342));
    Span4Mux_h I__2449 (
            .O(N__26342),
            .I(N__26339));
    Odrv4 I__2448 (
            .O(N__26339),
            .I(CONTROL_romAddReg_7_5));
    CascadeMux I__2447 (
            .O(N__26336),
            .I(DROM_ROMDATA_dintern_12ro_cascade_));
    InMux I__2446 (
            .O(N__26333),
            .I(N__26330));
    LocalMux I__2445 (
            .O(N__26330),
            .I(DROM_ROMDATA_dintern_12ro));
    IoInMux I__2444 (
            .O(N__26327),
            .I(N__26324));
    LocalMux I__2443 (
            .O(N__26324),
            .I(N__26321));
    Span4Mux_s3_h I__2442 (
            .O(N__26321),
            .I(N__26317));
    IoInMux I__2441 (
            .O(N__26320),
            .I(N__26314));
    Span4Mux_v I__2440 (
            .O(N__26317),
            .I(N__26311));
    LocalMux I__2439 (
            .O(N__26314),
            .I(N__26308));
    Sp12to4 I__2438 (
            .O(N__26311),
            .I(N__26305));
    Span4Mux_s3_h I__2437 (
            .O(N__26308),
            .I(N__26302));
    Span12Mux_s11_h I__2436 (
            .O(N__26305),
            .I(N__26299));
    Span4Mux_h I__2435 (
            .O(N__26302),
            .I(N__26296));
    Span12Mux_h I__2434 (
            .O(N__26299),
            .I(N__26293));
    Span4Mux_v I__2433 (
            .O(N__26296),
            .I(N__26290));
    Span12Mux_v I__2432 (
            .O(N__26293),
            .I(N__26287));
    Span4Mux_v I__2431 (
            .O(N__26290),
            .I(N__26284));
    Odrv12 I__2430 (
            .O(N__26287),
            .I(bus_12));
    Odrv4 I__2429 (
            .O(N__26284),
            .I(bus_12));
    InMux I__2428 (
            .O(N__26279),
            .I(N__26276));
    LocalMux I__2427 (
            .O(N__26276),
            .I(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_2 ));
    InMux I__2426 (
            .O(N__26273),
            .I(N__26270));
    LocalMux I__2425 (
            .O(N__26270),
            .I(N__26266));
    InMux I__2424 (
            .O(N__26269),
            .I(N__26263));
    Span4Mux_h I__2423 (
            .O(N__26266),
            .I(N__26258));
    LocalMux I__2422 (
            .O(N__26263),
            .I(N__26258));
    Span4Mux_v I__2421 (
            .O(N__26258),
            .I(N__26255));
    Odrv4 I__2420 (
            .O(N__26255),
            .I(\DROM.ROMDATA.dintern_0_3_NEW_2 ));
    InMux I__2419 (
            .O(N__26252),
            .I(N__26249));
    LocalMux I__2418 (
            .O(N__26249),
            .I(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_3 ));
    InMux I__2417 (
            .O(N__26246),
            .I(N__26242));
    InMux I__2416 (
            .O(N__26245),
            .I(N__26239));
    LocalMux I__2415 (
            .O(N__26242),
            .I(N__26234));
    LocalMux I__2414 (
            .O(N__26239),
            .I(N__26234));
    Span4Mux_v I__2413 (
            .O(N__26234),
            .I(N__26231));
    Odrv4 I__2412 (
            .O(N__26231),
            .I(\DROM.ROMDATA.dintern_0_3_NEW_3 ));
    IoInMux I__2411 (
            .O(N__26228),
            .I(N__26225));
    LocalMux I__2410 (
            .O(N__26225),
            .I(N__26221));
    IoInMux I__2409 (
            .O(N__26224),
            .I(N__26218));
    IoSpan4Mux I__2408 (
            .O(N__26221),
            .I(N__26215));
    LocalMux I__2407 (
            .O(N__26218),
            .I(N__26212));
    Span4Mux_s2_h I__2406 (
            .O(N__26215),
            .I(N__26209));
    IoSpan4Mux I__2405 (
            .O(N__26212),
            .I(N__26206));
    Sp12to4 I__2404 (
            .O(N__26209),
            .I(N__26203));
    Span4Mux_s0_h I__2403 (
            .O(N__26206),
            .I(N__26200));
    Span12Mux_s10_h I__2402 (
            .O(N__26203),
            .I(N__26197));
    Span4Mux_h I__2401 (
            .O(N__26200),
            .I(N__26194));
    Span12Mux_h I__2400 (
            .O(N__26197),
            .I(N__26191));
    Span4Mux_h I__2399 (
            .O(N__26194),
            .I(N__26188));
    Span12Mux_v I__2398 (
            .O(N__26191),
            .I(N__26185));
    Span4Mux_v I__2397 (
            .O(N__26188),
            .I(N__26182));
    Odrv12 I__2396 (
            .O(N__26185),
            .I(bus_10));
    Odrv4 I__2395 (
            .O(N__26182),
            .I(bus_10));
    IoInMux I__2394 (
            .O(N__26177),
            .I(N__26174));
    LocalMux I__2393 (
            .O(N__26174),
            .I(N__26171));
    Span4Mux_s0_h I__2392 (
            .O(N__26171),
            .I(N__26168));
    Span4Mux_h I__2391 (
            .O(N__26168),
            .I(N__26165));
    Span4Mux_h I__2390 (
            .O(N__26165),
            .I(N__26162));
    Odrv4 I__2389 (
            .O(N__26162),
            .I(gpuAddress_0));
    IoInMux I__2388 (
            .O(N__26159),
            .I(N__26156));
    LocalMux I__2387 (
            .O(N__26156),
            .I(N__26153));
    Span12Mux_s8_h I__2386 (
            .O(N__26153),
            .I(N__26150));
    Odrv12 I__2385 (
            .O(N__26150),
            .I(gpuAddress_1));
    InMux I__2384 (
            .O(N__26147),
            .I(N__26141));
    InMux I__2383 (
            .O(N__26146),
            .I(N__26141));
    LocalMux I__2382 (
            .O(N__26141),
            .I(DROM_ROMDATA_dintern_8ro));
    IoInMux I__2381 (
            .O(N__26138),
            .I(N__26135));
    LocalMux I__2380 (
            .O(N__26135),
            .I(N__26132));
    Span12Mux_s8_h I__2379 (
            .O(N__26132),
            .I(N__26128));
    IoInMux I__2378 (
            .O(N__26131),
            .I(N__26125));
    Span12Mux_v I__2377 (
            .O(N__26128),
            .I(N__26122));
    LocalMux I__2376 (
            .O(N__26125),
            .I(N__26119));
    Span12Mux_h I__2375 (
            .O(N__26122),
            .I(N__26116));
    Span12Mux_s8_h I__2374 (
            .O(N__26119),
            .I(N__26113));
    Odrv12 I__2373 (
            .O(N__26116),
            .I(bus_8));
    Odrv12 I__2372 (
            .O(N__26113),
            .I(bus_8));
    InMux I__2371 (
            .O(N__26108),
            .I(N__26102));
    InMux I__2370 (
            .O(N__26107),
            .I(N__26102));
    LocalMux I__2369 (
            .O(N__26102),
            .I(\DROM.ROMDATA.dintern_0_0_NEW_1 ));
    InMux I__2368 (
            .O(N__26099),
            .I(N__26096));
    LocalMux I__2367 (
            .O(N__26096),
            .I(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_1 ));
    InMux I__2366 (
            .O(N__26093),
            .I(N__26089));
    InMux I__2365 (
            .O(N__26092),
            .I(N__26086));
    LocalMux I__2364 (
            .O(N__26089),
            .I(N__26081));
    LocalMux I__2363 (
            .O(N__26086),
            .I(N__26081));
    Span4Mux_v I__2362 (
            .O(N__26081),
            .I(N__26078));
    Odrv4 I__2361 (
            .O(N__26078),
            .I(\DROM.ROMDATA.dintern_0_2_NEW_0 ));
    InMux I__2360 (
            .O(N__26075),
            .I(N__26072));
    LocalMux I__2359 (
            .O(N__26072),
            .I(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_0 ));
    InMux I__2358 (
            .O(N__26069),
            .I(N__26066));
    LocalMux I__2357 (
            .O(N__26066),
            .I(\ALU.log_1_3cf0_1_10 ));
    CascadeMux I__2356 (
            .O(N__26063),
            .I(\ALU.log_1_3cf0_10_cascade_ ));
    InMux I__2355 (
            .O(N__26060),
            .I(N__26057));
    LocalMux I__2354 (
            .O(N__26057),
            .I(\ALU.log_1_3cf1_10 ));
    InMux I__2353 (
            .O(N__26054),
            .I(N__26051));
    LocalMux I__2352 (
            .O(N__26051),
            .I(\ALU.log_1_3cf1_1_10 ));
    CascadeMux I__2351 (
            .O(N__26048),
            .I(\CONTROL.bus_7_a0_2_8_cascade_ ));
    CascadeMux I__2350 (
            .O(N__26045),
            .I(N__26042));
    InMux I__2349 (
            .O(N__26042),
            .I(N__26039));
    LocalMux I__2348 (
            .O(N__26039),
            .I(N__26036));
    Odrv12 I__2347 (
            .O(N__26036),
            .I(\ALU.status_18_cry_8_c_RNOZ0 ));
    CascadeMux I__2346 (
            .O(N__26033),
            .I(DROM_ROMDATA_dintern_8ro_cascade_));
    CascadeMux I__2345 (
            .O(N__26030),
            .I(\ALU.operand2_12_cascade_ ));
    CascadeMux I__2344 (
            .O(N__26027),
            .I(\ALU.N_126_cascade_ ));
    CascadeMux I__2343 (
            .O(N__26024),
            .I(\ALU.c_RNI670LZ0Z_12_cascade_ ));
    InMux I__2342 (
            .O(N__26021),
            .I(N__26018));
    LocalMux I__2341 (
            .O(N__26018),
            .I(\ALU.operand2_7_ns_1_12 ));
    CascadeMux I__2340 (
            .O(N__26015),
            .I(N__26012));
    InMux I__2339 (
            .O(N__26012),
            .I(N__26009));
    LocalMux I__2338 (
            .O(N__26009),
            .I(\ALU.d_RNI8FCTZ0Z_12 ));
    CascadeMux I__2337 (
            .O(N__26006),
            .I(N__26003));
    InMux I__2336 (
            .O(N__26003),
            .I(N__26000));
    LocalMux I__2335 (
            .O(N__26000),
            .I(\ALU.operand2_12 ));
    CascadeMux I__2334 (
            .O(N__25997),
            .I(N__25994));
    InMux I__2333 (
            .O(N__25994),
            .I(N__25991));
    LocalMux I__2332 (
            .O(N__25991),
            .I(N__25988));
    Span4Mux_v I__2331 (
            .O(N__25988),
            .I(N__25985));
    Odrv4 I__2330 (
            .O(N__25985),
            .I(\ALU.status_18_cry_12_c_RNOZ0 ));
    CascadeMux I__2329 (
            .O(N__25982),
            .I(N__25979));
    InMux I__2328 (
            .O(N__25979),
            .I(N__25976));
    LocalMux I__2327 (
            .O(N__25976),
            .I(\ALU.status_18_cry_10_c_RNOZ0 ));
    CascadeMux I__2326 (
            .O(N__25973),
            .I(N__25970));
    InMux I__2325 (
            .O(N__25970),
            .I(N__25967));
    LocalMux I__2324 (
            .O(N__25967),
            .I(\ALU.status_18_cry_13_c_RNOZ0 ));
    CascadeMux I__2323 (
            .O(N__25964),
            .I(\CONTROL.busState_1_RNIG7366Z0Z_2_cascade_ ));
    InMux I__2322 (
            .O(N__25961),
            .I(N__25958));
    LocalMux I__2321 (
            .O(N__25958),
            .I(\CONTROL.busState_1_RNI1JVK1_0Z0Z_2 ));
    InMux I__2320 (
            .O(N__25955),
            .I(N__25952));
    LocalMux I__2319 (
            .O(N__25952),
            .I(N__25949));
    Span4Mux_v I__2318 (
            .O(N__25949),
            .I(N__25946));
    Span4Mux_v I__2317 (
            .O(N__25946),
            .I(N__25943));
    Span4Mux_v I__2316 (
            .O(N__25943),
            .I(N__25940));
    Span4Mux_v I__2315 (
            .O(N__25940),
            .I(N__25937));
    IoSpan4Mux I__2314 (
            .O(N__25937),
            .I(N__25934));
    IoSpan4Mux I__2313 (
            .O(N__25934),
            .I(N__25931));
    Odrv4 I__2312 (
            .O(N__25931),
            .I(gpuOut_c_5));
    InMux I__2311 (
            .O(N__25928),
            .I(N__25925));
    LocalMux I__2310 (
            .O(N__25925),
            .I(\CONTROL.N_166 ));
    CascadeMux I__2309 (
            .O(N__25922),
            .I(N__25918));
    InMux I__2308 (
            .O(N__25921),
            .I(N__25915));
    InMux I__2307 (
            .O(N__25918),
            .I(N__25912));
    LocalMux I__2306 (
            .O(N__25915),
            .I(N__25909));
    LocalMux I__2305 (
            .O(N__25912),
            .I(N__25906));
    Span4Mux_v I__2304 (
            .O(N__25909),
            .I(N__25901));
    Span4Mux_v I__2303 (
            .O(N__25906),
            .I(N__25901));
    Sp12to4 I__2302 (
            .O(N__25901),
            .I(N__25898));
    Span12Mux_h I__2301 (
            .O(N__25898),
            .I(N__25895));
    Span12Mux_v I__2300 (
            .O(N__25895),
            .I(N__25892));
    Odrv12 I__2299 (
            .O(N__25892),
            .I(D5_in_c));
    CascadeMux I__2298 (
            .O(N__25889),
            .I(\CONTROL.N_166_cascade_ ));
    CascadeMux I__2297 (
            .O(N__25886),
            .I(N__25883));
    InMux I__2296 (
            .O(N__25883),
            .I(N__25880));
    LocalMux I__2295 (
            .O(N__25880),
            .I(romOut_5));
    CascadeMux I__2294 (
            .O(N__25877),
            .I(N__25874));
    InMux I__2293 (
            .O(N__25874),
            .I(N__25871));
    LocalMux I__2292 (
            .O(N__25871),
            .I(\ALU.combOperand2_i_11 ));
    CascadeMux I__2291 (
            .O(N__25868),
            .I(N__25865));
    InMux I__2290 (
            .O(N__25865),
            .I(N__25862));
    LocalMux I__2289 (
            .O(N__25862),
            .I(\ALU.combOperand2_i_14 ));
    CascadeMux I__2288 (
            .O(N__25859),
            .I(N__25856));
    InMux I__2287 (
            .O(N__25856),
            .I(N__25853));
    LocalMux I__2286 (
            .O(N__25853),
            .I(\ALU.combOperand2_i_15 ));
    InMux I__2285 (
            .O(N__25850),
            .I(bfn_9_13_0_));
    InMux I__2284 (
            .O(N__25847),
            .I(N__25844));
    LocalMux I__2283 (
            .O(N__25844),
            .I(\ALU.status_17_I_45_c_RNOZ0 ));
    InMux I__2282 (
            .O(N__25841),
            .I(N__25838));
    LocalMux I__2281 (
            .O(N__25838),
            .I(\ALU.combOperand2_i_1 ));
    CascadeMux I__2280 (
            .O(N__25835),
            .I(N__25832));
    InMux I__2279 (
            .O(N__25832),
            .I(N__25829));
    LocalMux I__2278 (
            .O(N__25829),
            .I(N__25826));
    Odrv4 I__2277 (
            .O(N__25826),
            .I(\ALU.status_17_I_27_c_RNOZ0 ));
    InMux I__2276 (
            .O(N__25823),
            .I(N__25820));
    LocalMux I__2275 (
            .O(N__25820),
            .I(\ALU.combOperand2_i_7 ));
    InMux I__2274 (
            .O(N__25817),
            .I(bfn_9_10_0_));
    InMux I__2273 (
            .O(N__25814),
            .I(clkdiv_cry_22));
    IoInMux I__2272 (
            .O(N__25811),
            .I(N__25808));
    LocalMux I__2271 (
            .O(N__25808),
            .I(N__25805));
    Span12Mux_s6_v I__2270 (
            .O(N__25805),
            .I(N__25801));
    InMux I__2269 (
            .O(N__25804),
            .I(N__25798));
    Odrv12 I__2268 (
            .O(N__25801),
            .I(GPIO3_c));
    LocalMux I__2267 (
            .O(N__25798),
            .I(GPIO3_c));
    IoInMux I__2266 (
            .O(N__25793),
            .I(N__25788));
    IoInMux I__2265 (
            .O(N__25792),
            .I(N__25785));
    IoInMux I__2264 (
            .O(N__25791),
            .I(N__25782));
    LocalMux I__2263 (
            .O(N__25788),
            .I(B_OE_c_i));
    LocalMux I__2262 (
            .O(N__25785),
            .I(B_OE_c_i));
    LocalMux I__2261 (
            .O(N__25782),
            .I(B_OE_c_i));
    IoInMux I__2260 (
            .O(N__25775),
            .I(N__25772));
    LocalMux I__2259 (
            .O(N__25772),
            .I(N__25769));
    Span4Mux_s2_h I__2258 (
            .O(N__25769),
            .I(N__25766));
    Sp12to4 I__2257 (
            .O(N__25766),
            .I(N__25762));
    InMux I__2256 (
            .O(N__25765),
            .I(N__25759));
    Span12Mux_s11_v I__2255 (
            .O(N__25762),
            .I(N__25756));
    LocalMux I__2254 (
            .O(N__25759),
            .I(N__25753));
    Odrv12 I__2253 (
            .O(N__25756),
            .I(B_OE_c));
    Odrv4 I__2252 (
            .O(N__25753),
            .I(B_OE_c));
    IoInMux I__2251 (
            .O(N__25748),
            .I(N__25745));
    LocalMux I__2250 (
            .O(N__25745),
            .I(N__25742));
    Span4Mux_s3_h I__2249 (
            .O(N__25742),
            .I(N__25739));
    Span4Mux_v I__2248 (
            .O(N__25739),
            .I(N__25736));
    Odrv4 I__2247 (
            .O(N__25736),
            .I(gpuAddress_11));
    IoInMux I__2246 (
            .O(N__25733),
            .I(N__25730));
    LocalMux I__2245 (
            .O(N__25730),
            .I(N__25727));
    Span4Mux_s2_h I__2244 (
            .O(N__25727),
            .I(N__25724));
    Span4Mux_v I__2243 (
            .O(N__25724),
            .I(N__25721));
    Span4Mux_h I__2242 (
            .O(N__25721),
            .I(N__25718));
    Odrv4 I__2241 (
            .O(N__25718),
            .I(gpuAddress_14));
    IoInMux I__2240 (
            .O(N__25715),
            .I(N__25712));
    LocalMux I__2239 (
            .O(N__25712),
            .I(N__25709));
    Span12Mux_s6_h I__2238 (
            .O(N__25709),
            .I(N__25706));
    Odrv12 I__2237 (
            .O(N__25706),
            .I(gpuAddress_9));
    IoInMux I__2236 (
            .O(N__25703),
            .I(N__25700));
    LocalMux I__2235 (
            .O(N__25700),
            .I(N__25697));
    IoSpan4Mux I__2234 (
            .O(N__25697),
            .I(N__25694));
    Span4Mux_s3_h I__2233 (
            .O(N__25694),
            .I(N__25691));
    Odrv4 I__2232 (
            .O(N__25691),
            .I(N_6_0));
    IoInMux I__2231 (
            .O(N__25688),
            .I(N__25685));
    LocalMux I__2230 (
            .O(N__25685),
            .I(N__25681));
    IoInMux I__2229 (
            .O(N__25684),
            .I(N__25678));
    IoSpan4Mux I__2228 (
            .O(N__25681),
            .I(N__25673));
    LocalMux I__2227 (
            .O(N__25678),
            .I(N__25673));
    Span4Mux_s2_h I__2226 (
            .O(N__25673),
            .I(N__25669));
    IoInMux I__2225 (
            .O(N__25672),
            .I(N__25666));
    Span4Mux_h I__2224 (
            .O(N__25669),
            .I(N__25663));
    LocalMux I__2223 (
            .O(N__25666),
            .I(N__25660));
    Odrv4 I__2222 (
            .O(N__25663),
            .I(RAM_un1_WR_i));
    Odrv12 I__2221 (
            .O(N__25660),
            .I(RAM_un1_WR_i));
    InMux I__2220 (
            .O(N__25655),
            .I(N__25652));
    LocalMux I__2219 (
            .O(N__25652),
            .I(clkdivZ0Z_15));
    InMux I__2218 (
            .O(N__25649),
            .I(clkdiv_cry_14));
    InMux I__2217 (
            .O(N__25646),
            .I(N__25643));
    LocalMux I__2216 (
            .O(N__25643),
            .I(clkdivZ0Z_16));
    InMux I__2215 (
            .O(N__25640),
            .I(bfn_1_19_0_));
    InMux I__2214 (
            .O(N__25637),
            .I(N__25634));
    LocalMux I__2213 (
            .O(N__25634),
            .I(clkdivZ0Z_17));
    InMux I__2212 (
            .O(N__25631),
            .I(clkdiv_cry_16));
    InMux I__2211 (
            .O(N__25628),
            .I(N__25625));
    LocalMux I__2210 (
            .O(N__25625),
            .I(clkdivZ0Z_18));
    InMux I__2209 (
            .O(N__25622),
            .I(clkdiv_cry_17));
    InMux I__2208 (
            .O(N__25619),
            .I(N__25616));
    LocalMux I__2207 (
            .O(N__25616),
            .I(clkdivZ0Z_19));
    InMux I__2206 (
            .O(N__25613),
            .I(clkdiv_cry_18));
    InMux I__2205 (
            .O(N__25610),
            .I(N__25607));
    LocalMux I__2204 (
            .O(N__25607),
            .I(clkdivZ0Z_20));
    InMux I__2203 (
            .O(N__25604),
            .I(clkdiv_cry_19));
    InMux I__2202 (
            .O(N__25601),
            .I(N__25598));
    LocalMux I__2201 (
            .O(N__25598),
            .I(clkdivZ0Z_21));
    InMux I__2200 (
            .O(N__25595),
            .I(clkdiv_cry_20));
    InMux I__2199 (
            .O(N__25592),
            .I(N__25589));
    LocalMux I__2198 (
            .O(N__25589),
            .I(clkdivZ0Z_22));
    InMux I__2197 (
            .O(N__25586),
            .I(clkdiv_cry_21));
    InMux I__2196 (
            .O(N__25583),
            .I(N__25580));
    LocalMux I__2195 (
            .O(N__25580),
            .I(clkdivZ0Z_7));
    InMux I__2194 (
            .O(N__25577),
            .I(clkdiv_cry_6));
    InMux I__2193 (
            .O(N__25574),
            .I(N__25571));
    LocalMux I__2192 (
            .O(N__25571),
            .I(clkdivZ0Z_8));
    InMux I__2191 (
            .O(N__25568),
            .I(bfn_1_18_0_));
    InMux I__2190 (
            .O(N__25565),
            .I(N__25562));
    LocalMux I__2189 (
            .O(N__25562),
            .I(clkdivZ0Z_9));
    InMux I__2188 (
            .O(N__25559),
            .I(clkdiv_cry_8));
    InMux I__2187 (
            .O(N__25556),
            .I(N__25553));
    LocalMux I__2186 (
            .O(N__25553),
            .I(clkdivZ0Z_10));
    InMux I__2185 (
            .O(N__25550),
            .I(clkdiv_cry_9));
    InMux I__2184 (
            .O(N__25547),
            .I(N__25544));
    LocalMux I__2183 (
            .O(N__25544),
            .I(clkdivZ0Z_11));
    InMux I__2182 (
            .O(N__25541),
            .I(clkdiv_cry_10));
    InMux I__2181 (
            .O(N__25538),
            .I(N__25535));
    LocalMux I__2180 (
            .O(N__25535),
            .I(clkdivZ0Z_12));
    InMux I__2179 (
            .O(N__25532),
            .I(clkdiv_cry_11));
    InMux I__2178 (
            .O(N__25529),
            .I(N__25526));
    LocalMux I__2177 (
            .O(N__25526),
            .I(clkdivZ0Z_13));
    InMux I__2176 (
            .O(N__25523),
            .I(clkdiv_cry_12));
    InMux I__2175 (
            .O(N__25520),
            .I(N__25517));
    LocalMux I__2174 (
            .O(N__25517),
            .I(clkdivZ0Z_14));
    InMux I__2173 (
            .O(N__25514),
            .I(clkdiv_cry_13));
    InMux I__2172 (
            .O(N__25511),
            .I(N__25508));
    LocalMux I__2171 (
            .O(N__25508),
            .I(clkdivZ0Z_0));
    InMux I__2170 (
            .O(N__25505),
            .I(bfn_1_17_0_));
    InMux I__2169 (
            .O(N__25502),
            .I(N__25499));
    LocalMux I__2168 (
            .O(N__25499),
            .I(clkdivZ0Z_1));
    InMux I__2167 (
            .O(N__25496),
            .I(clkdiv_cry_0));
    InMux I__2166 (
            .O(N__25493),
            .I(N__25490));
    LocalMux I__2165 (
            .O(N__25490),
            .I(clkdivZ0Z_2));
    InMux I__2164 (
            .O(N__25487),
            .I(clkdiv_cry_1));
    InMux I__2163 (
            .O(N__25484),
            .I(N__25481));
    LocalMux I__2162 (
            .O(N__25481),
            .I(clkdivZ0Z_3));
    InMux I__2161 (
            .O(N__25478),
            .I(clkdiv_cry_2));
    InMux I__2160 (
            .O(N__25475),
            .I(N__25472));
    LocalMux I__2159 (
            .O(N__25472),
            .I(clkdivZ0Z_4));
    InMux I__2158 (
            .O(N__25469),
            .I(clkdiv_cry_3));
    InMux I__2157 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__2156 (
            .O(N__25463),
            .I(clkdivZ0Z_5));
    InMux I__2155 (
            .O(N__25460),
            .I(clkdiv_cry_4));
    InMux I__2154 (
            .O(N__25457),
            .I(N__25454));
    LocalMux I__2153 (
            .O(N__25454),
            .I(clkdivZ0Z_6));
    InMux I__2152 (
            .O(N__25451),
            .I(clkdiv_cry_5));
    INV \INVCONTROL.ramAddReg_6C  (
            .O(\INVCONTROL.ramAddReg_6C_net ),
            .I(N__73250));
    INV \INVCONTROL.results_2C  (
            .O(\INVCONTROL.results_2C_net ),
            .I(N__73249));
    INV \INVCONTROL.results_1C  (
            .O(\INVCONTROL.results_1C_net ),
            .I(N__73238));
    INV \INVCONTROL.increment_1C  (
            .O(\INVCONTROL.increment_1C_net ),
            .I(N__73207));
    INV \INVCONTROL.aluOperation_6C  (
            .O(\INVCONTROL.aluOperation_6C_net ),
            .I(N__73216));
    INV \INVCONTROL.ramAddReg_3C  (
            .O(\INVCONTROL.ramAddReg_3C_net ),
            .I(N__73206));
    INV \INVCONTROL.dout_13C  (
            .O(\INVCONTROL.dout_13C_net ),
            .I(N__73198));
    INV \INVCONTROL.increment_0C  (
            .O(\INVCONTROL.increment_0C_net ),
            .I(N__73245));
    INV \INVCONTROL.dout_9C  (
            .O(\INVCONTROL.dout_9C_net ),
            .I(N__73191));
    INV \INVCONTROL.operand2_fast_ne_1C  (
            .O(\INVCONTROL.operand2_fast_ne_1C_net ),
            .I(N__73182));
    INV \INVCONTROL.operand2_2_rep1_neC  (
            .O(\INVCONTROL.operand2_2_rep1_neC_net ),
            .I(N__73171));
    INV \INVCONTROL.addrstackptr_2C  (
            .O(\INVCONTROL.addrstackptr_2C_net ),
            .I(N__73215));
    INV \INVCONTROL.aluOperation_ne_5C  (
            .O(\INVCONTROL.aluOperation_ne_5C_net ),
            .I(N__73197));
    INV \INVCONTROL.dout_2C  (
            .O(\INVCONTROL.dout_2C_net ),
            .I(N__73201));
    INV \INVCONTROL.aluOperation_4C  (
            .O(\INVCONTROL.aluOperation_4C_net ),
            .I(N__73195));
    INV \INVCONTROL.aluParams_1_ne_1C  (
            .O(\INVCONTROL.aluParams_1_ne_1C_net ),
            .I(N__73189));
    INV \INVCONTROL.aluParams_1_0C  (
            .O(\INVCONTROL.aluParams_1_0C_net ),
            .I(N__73178));
    INV \INVCONTROL.operand1_ne_0C  (
            .O(\INVCONTROL.operand1_ne_0C_net ),
            .I(N__73167));
    INV \INVCONTROL.operand2_fast_ne_2C  (
            .O(\INVCONTROL.operand2_fast_ne_2C_net ),
            .I(N__73152));
    INV \INVCONTROL.ramWriteC  (
            .O(\INVCONTROL.ramWriteC_net ),
            .I(N__73223));
    INV \INVCONTROL.aluOperation_ne_1C  (
            .O(\INVCONTROL.aluOperation_ne_1C_net ),
            .I(N__73214));
    INV \INVCONTROL.addrstackptr_3C  (
            .O(\INVCONTROL.addrstackptr_3C_net ),
            .I(N__73205));
    INV \INVCONTROL.operand1_fast_ne_1C  (
            .O(\INVCONTROL.operand1_fast_ne_1C_net ),
            .I(N__73170));
    INV \INVCONTROL.tempCounter_4C  (
            .O(\INVCONTROL.tempCounter_4C_net ),
            .I(N__73255));
    INV \INVCONTROL.tempCounter_0C  (
            .O(\INVCONTROL.tempCounter_0C_net ),
            .I(N__73244));
    INV \INVCONTROL.dout_1C  (
            .O(\INVCONTROL.dout_1C_net ),
            .I(N__73222));
    INV \INVCONTROL.busState_1_1C  (
            .O(\INVCONTROL.busState_1_1C_net ),
            .I(N__73213));
    INV \INVCONTROL.busState_1_2C  (
            .O(\INVCONTROL.busState_1_2C_net ),
            .I(N__73204));
    INV \INVCONTROL.operand1_ne_1C  (
            .O(\INVCONTROL.operand1_ne_1C_net ),
            .I(N__73180));
    INV \INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C  (
            .O(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C_net ),
            .I(N__73149));
    INV \INVCONTROL.ramAddReg_14C  (
            .O(\INVCONTROL.ramAddReg_14C_net ),
            .I(N__73272));
    INV \INVCONTROL.addrstackptr_1C  (
            .O(\INVCONTROL.addrstackptr_1C_net ),
            .I(N__73254));
    INV \INVCONTROL.ramAddReg_0C  (
            .O(\INVCONTROL.ramAddReg_0C_net ),
            .I(N__73243));
    INV \INVCONTROL.dout_15C  (
            .O(\INVCONTROL.dout_15C_net ),
            .I(N__73231));
    INV \INVCONTROL.dout_10C  (
            .O(\INVCONTROL.dout_10C_net ),
            .I(N__73221));
    INV \INVCONTROL.aluReadBusC  (
            .O(\INVCONTROL.aluReadBusC_net ),
            .I(N__73203));
    INV \INVCONTROL.dout_11C  (
            .O(\INVCONTROL.dout_11C_net ),
            .I(N__73196));
    INV \INVCONTROL.dout_14C  (
            .O(\INVCONTROL.dout_14C_net ),
            .I(N__73179));
    INV \INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C  (
            .O(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C_net ),
            .I(N__73169));
    INV \INVCONTROL.addrstackptr_4C  (
            .O(\INVCONTROL.addrstackptr_4C_net ),
            .I(N__73242));
    INV \INVCONTROL.ramAddReg_5C  (
            .O(\INVCONTROL.ramAddReg_5C_net ),
            .I(N__73230));
    INV \INVCONTROL.gpuWriteC  (
            .O(\INVCONTROL.gpuWriteC_net ),
            .I(N__73220));
    INV \INVCONTROL.gpuAddReg_2C  (
            .O(\INVCONTROL.gpuAddReg_2C_net ),
            .I(N__73212));
    INV \INVCONTROL.dout_7C  (
            .O(\INVCONTROL.dout_7C_net ),
            .I(N__73202));
    INV \INVCONTROL.addrstackptr_0C  (
            .O(\INVCONTROL.addrstackptr_0C_net ),
            .I(N__73139));
    INV \INVCONTROL.tempCounter_10C  (
            .O(\INVCONTROL.tempCounter_10C_net ),
            .I(N__73276));
    INV \INVCONTROL.ramAddReg_13C  (
            .O(\INVCONTROL.ramAddReg_13C_net ),
            .I(N__73229));
    INV \INVCONTROL.busState_1_0C  (
            .O(\INVCONTROL.busState_1_0C_net ),
            .I(N__73219));
    INV \INVCONTROL.romAddReg_10C  (
            .O(\INVCONTROL.romAddReg_10C_net ),
            .I(N__73211));
    INV \INVCONTROL.tempCounter_11C  (
            .O(\INVCONTROL.tempCounter_11C_net ),
            .I(N__73275));
    INV \INVCONTROL.addrstackptr_5C  (
            .O(\INVCONTROL.addrstackptr_5C_net ),
            .I(N__73262));
    INV \INVCONTROL.dout_6C  (
            .O(\INVCONTROL.dout_6C_net ),
            .I(N__73252));
    INV \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C  (
            .O(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .I(N__73241));
    INV \INVCONTROL.aluOperation_ne_0C  (
            .O(\INVCONTROL.aluOperation_ne_0C_net ),
            .I(N__73228));
    INV \INVCONTROL.romAddReg_13C  (
            .O(\INVCONTROL.romAddReg_13C_net ),
            .I(N__73218));
    INV \INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C  (
            .O(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C_net ),
            .I(N__73210));
    INV \INVCONTROL.tempCounter_13C  (
            .O(\INVCONTROL.tempCounter_13C_net ),
            .I(N__73282));
    INV \INVCONTROL.addrstackptr_6C  (
            .O(\INVCONTROL.addrstackptr_6C_net ),
            .I(N__73277));
    INV \INVCONTROL.dout_3C  (
            .O(\INVCONTROL.dout_3C_net ),
            .I(N__73268));
    INV \INVCONTROL.gpuAddReg_0C  (
            .O(\INVCONTROL.gpuAddReg_0C_net ),
            .I(N__73261));
    INV \INVCONTROL.aluOperation_3C  (
            .O(\INVCONTROL.aluOperation_3C_net ),
            .I(N__73251));
    INV \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C  (
            .O(\INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net ),
            .I(N__73240));
    INV \INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C  (
            .O(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C_net ),
            .I(N__73227));
    INV \INVCONTROL.dout_5C  (
            .O(\INVCONTROL.dout_5C_net ),
            .I(N__73200));
    INV \INVCONTROL.gpuAddReg_9C  (
            .O(\INVCONTROL.gpuAddReg_9C_net ),
            .I(N__73273));
    INV \INVCONTROL.gpuAddReg_14C  (
            .O(\INVCONTROL.gpuAddReg_14C_net ),
            .I(N__73259));
    INV \INVCONTROL.gpuAddReg_11C  (
            .O(\INVCONTROL.gpuAddReg_11C_net ),
            .I(N__73280));
    INV \INVDROM.ROMDATA.dintern_0_0RCLKN  (
            .O(\INVDROM.ROMDATA.dintern_0_0RCLKN_net ),
            .I(N__73239));
    INV \INVDROM.ROMDATA.dintern_0_1RCLKN  (
            .O(\INVDROM.ROMDATA.dintern_0_1RCLKN_net ),
            .I(N__73260));
    INV \INVDROM.ROMDATA.dintern_0_2RCLKN  (
            .O(\INVDROM.ROMDATA.dintern_0_2RCLKN_net ),
            .I(N__73274));
    INV \INVDROM.ROMDATA.dintern_0_3RCLKN  (
            .O(\INVDROM.ROMDATA.dintern_0_3RCLKN_net ),
            .I(N__73281));
    INV \INVCONTROL.addrstack_addrstack_0_0RCLKN  (
            .O(\INVCONTROL.addrstack_addrstack_0_0RCLKN_net ),
            .I(N__73291));
    defparam IN_MUX_bfv_23_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_14_0_));
    defparam IN_MUX_bfv_23_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_15_0_ (
            .carryinitin(\ALU.addsub_cry_6 ),
            .carryinitout(bfn_23_15_0_));
    defparam IN_MUX_bfv_23_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_16_0_ (
            .carryinitin(\ALU.addsub_cry_14 ),
            .carryinitout(bfn_23_16_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\CONTROL.programCounter_1_cry_7 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\ALU.status_18_cry_7 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\ALU.status_18_4 ),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\ALU.status_17_data_tmp_7 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\ALU.mult_3_c10 ),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\ALU.mult_1_c8 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_20_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_10_0_));
    defparam IN_MUX_bfv_19_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_10_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\ALU.mult_7_c14 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\ALU.mult_5_c12 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(clkdiv_cry_7),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(clkdiv_cry_15),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_23_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_7_0_));
    defparam IN_MUX_bfv_23_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_8_0_ (
            .carryinitin(\ALU.status_19_cry_7 ),
            .carryinitout(bfn_23_8_0_));
    defparam IN_MUX_bfv_23_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_9_0_ (
            .carryinitin(\ALU.status_19Z0Z_5 ),
            .carryinitout(bfn_23_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\ALU.mult_17_c9 ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\ALU.mult_25_c11 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_19_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_9_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\ALU.mult_19_c13 ),
            .carryinitout(bfn_15_10_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam clkdiv_0_LC_1_17_0.C_ON=1'b1;
    defparam clkdiv_0_LC_1_17_0.SEQ_MODE=4'b1000;
    defparam clkdiv_0_LC_1_17_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_0_LC_1_17_0 (
            .in0(_gnd_net_),
            .in1(N__25511),
            .in2(_gnd_net_),
            .in3(N__25505),
            .lcout(clkdivZ0Z_0),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(clkdiv_cry_0),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_1_LC_1_17_1.C_ON=1'b1;
    defparam clkdiv_1_LC_1_17_1.SEQ_MODE=4'b1000;
    defparam clkdiv_1_LC_1_17_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_1_LC_1_17_1 (
            .in0(_gnd_net_),
            .in1(N__25502),
            .in2(_gnd_net_),
            .in3(N__25496),
            .lcout(clkdivZ0Z_1),
            .ltout(),
            .carryin(clkdiv_cry_0),
            .carryout(clkdiv_cry_1),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_2_LC_1_17_2.C_ON=1'b1;
    defparam clkdiv_2_LC_1_17_2.SEQ_MODE=4'b1000;
    defparam clkdiv_2_LC_1_17_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_2_LC_1_17_2 (
            .in0(_gnd_net_),
            .in1(N__25493),
            .in2(_gnd_net_),
            .in3(N__25487),
            .lcout(clkdivZ0Z_2),
            .ltout(),
            .carryin(clkdiv_cry_1),
            .carryout(clkdiv_cry_2),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_3_LC_1_17_3.C_ON=1'b1;
    defparam clkdiv_3_LC_1_17_3.SEQ_MODE=4'b1000;
    defparam clkdiv_3_LC_1_17_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_3_LC_1_17_3 (
            .in0(_gnd_net_),
            .in1(N__25484),
            .in2(_gnd_net_),
            .in3(N__25478),
            .lcout(clkdivZ0Z_3),
            .ltout(),
            .carryin(clkdiv_cry_2),
            .carryout(clkdiv_cry_3),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_4_LC_1_17_4.C_ON=1'b1;
    defparam clkdiv_4_LC_1_17_4.SEQ_MODE=4'b1000;
    defparam clkdiv_4_LC_1_17_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_4_LC_1_17_4 (
            .in0(_gnd_net_),
            .in1(N__25475),
            .in2(_gnd_net_),
            .in3(N__25469),
            .lcout(clkdivZ0Z_4),
            .ltout(),
            .carryin(clkdiv_cry_3),
            .carryout(clkdiv_cry_4),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_5_LC_1_17_5.C_ON=1'b1;
    defparam clkdiv_5_LC_1_17_5.SEQ_MODE=4'b1000;
    defparam clkdiv_5_LC_1_17_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_5_LC_1_17_5 (
            .in0(_gnd_net_),
            .in1(N__25466),
            .in2(_gnd_net_),
            .in3(N__25460),
            .lcout(clkdivZ0Z_5),
            .ltout(),
            .carryin(clkdiv_cry_4),
            .carryout(clkdiv_cry_5),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_6_LC_1_17_6.C_ON=1'b1;
    defparam clkdiv_6_LC_1_17_6.SEQ_MODE=4'b1000;
    defparam clkdiv_6_LC_1_17_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_6_LC_1_17_6 (
            .in0(_gnd_net_),
            .in1(N__25457),
            .in2(_gnd_net_),
            .in3(N__25451),
            .lcout(clkdivZ0Z_6),
            .ltout(),
            .carryin(clkdiv_cry_5),
            .carryout(clkdiv_cry_6),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_7_LC_1_17_7.C_ON=1'b1;
    defparam clkdiv_7_LC_1_17_7.SEQ_MODE=4'b1000;
    defparam clkdiv_7_LC_1_17_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_7_LC_1_17_7 (
            .in0(_gnd_net_),
            .in1(N__25583),
            .in2(_gnd_net_),
            .in3(N__25577),
            .lcout(clkdivZ0Z_7),
            .ltout(),
            .carryin(clkdiv_cry_6),
            .carryout(clkdiv_cry_7),
            .clk(N__73286),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_8_LC_1_18_0.C_ON=1'b1;
    defparam clkdiv_8_LC_1_18_0.SEQ_MODE=4'b1000;
    defparam clkdiv_8_LC_1_18_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_8_LC_1_18_0 (
            .in0(_gnd_net_),
            .in1(N__25574),
            .in2(_gnd_net_),
            .in3(N__25568),
            .lcout(clkdivZ0Z_8),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(clkdiv_cry_8),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_9_LC_1_18_1.C_ON=1'b1;
    defparam clkdiv_9_LC_1_18_1.SEQ_MODE=4'b1000;
    defparam clkdiv_9_LC_1_18_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_9_LC_1_18_1 (
            .in0(_gnd_net_),
            .in1(N__25565),
            .in2(_gnd_net_),
            .in3(N__25559),
            .lcout(clkdivZ0Z_9),
            .ltout(),
            .carryin(clkdiv_cry_8),
            .carryout(clkdiv_cry_9),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_10_LC_1_18_2.C_ON=1'b1;
    defparam clkdiv_10_LC_1_18_2.SEQ_MODE=4'b1000;
    defparam clkdiv_10_LC_1_18_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_10_LC_1_18_2 (
            .in0(_gnd_net_),
            .in1(N__25556),
            .in2(_gnd_net_),
            .in3(N__25550),
            .lcout(clkdivZ0Z_10),
            .ltout(),
            .carryin(clkdiv_cry_9),
            .carryout(clkdiv_cry_10),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_11_LC_1_18_3.C_ON=1'b1;
    defparam clkdiv_11_LC_1_18_3.SEQ_MODE=4'b1000;
    defparam clkdiv_11_LC_1_18_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_11_LC_1_18_3 (
            .in0(_gnd_net_),
            .in1(N__25547),
            .in2(_gnd_net_),
            .in3(N__25541),
            .lcout(clkdivZ0Z_11),
            .ltout(),
            .carryin(clkdiv_cry_10),
            .carryout(clkdiv_cry_11),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_12_LC_1_18_4.C_ON=1'b1;
    defparam clkdiv_12_LC_1_18_4.SEQ_MODE=4'b1000;
    defparam clkdiv_12_LC_1_18_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_12_LC_1_18_4 (
            .in0(_gnd_net_),
            .in1(N__25538),
            .in2(_gnd_net_),
            .in3(N__25532),
            .lcout(clkdivZ0Z_12),
            .ltout(),
            .carryin(clkdiv_cry_11),
            .carryout(clkdiv_cry_12),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_13_LC_1_18_5.C_ON=1'b1;
    defparam clkdiv_13_LC_1_18_5.SEQ_MODE=4'b1000;
    defparam clkdiv_13_LC_1_18_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_13_LC_1_18_5 (
            .in0(_gnd_net_),
            .in1(N__25529),
            .in2(_gnd_net_),
            .in3(N__25523),
            .lcout(clkdivZ0Z_13),
            .ltout(),
            .carryin(clkdiv_cry_12),
            .carryout(clkdiv_cry_13),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_14_LC_1_18_6.C_ON=1'b1;
    defparam clkdiv_14_LC_1_18_6.SEQ_MODE=4'b1000;
    defparam clkdiv_14_LC_1_18_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_14_LC_1_18_6 (
            .in0(_gnd_net_),
            .in1(N__25520),
            .in2(_gnd_net_),
            .in3(N__25514),
            .lcout(clkdivZ0Z_14),
            .ltout(),
            .carryin(clkdiv_cry_13),
            .carryout(clkdiv_cry_14),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_15_LC_1_18_7.C_ON=1'b1;
    defparam clkdiv_15_LC_1_18_7.SEQ_MODE=4'b1000;
    defparam clkdiv_15_LC_1_18_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_15_LC_1_18_7 (
            .in0(_gnd_net_),
            .in1(N__25655),
            .in2(_gnd_net_),
            .in3(N__25649),
            .lcout(clkdivZ0Z_15),
            .ltout(),
            .carryin(clkdiv_cry_14),
            .carryout(clkdiv_cry_15),
            .clk(N__73290),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_16_LC_1_19_0.C_ON=1'b1;
    defparam clkdiv_16_LC_1_19_0.SEQ_MODE=4'b1000;
    defparam clkdiv_16_LC_1_19_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_16_LC_1_19_0 (
            .in0(_gnd_net_),
            .in1(N__25646),
            .in2(_gnd_net_),
            .in3(N__25640),
            .lcout(clkdivZ0Z_16),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(clkdiv_cry_16),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_17_LC_1_19_1.C_ON=1'b1;
    defparam clkdiv_17_LC_1_19_1.SEQ_MODE=4'b1000;
    defparam clkdiv_17_LC_1_19_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_17_LC_1_19_1 (
            .in0(_gnd_net_),
            .in1(N__25637),
            .in2(_gnd_net_),
            .in3(N__25631),
            .lcout(clkdivZ0Z_17),
            .ltout(),
            .carryin(clkdiv_cry_16),
            .carryout(clkdiv_cry_17),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_18_LC_1_19_2.C_ON=1'b1;
    defparam clkdiv_18_LC_1_19_2.SEQ_MODE=4'b1000;
    defparam clkdiv_18_LC_1_19_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_18_LC_1_19_2 (
            .in0(_gnd_net_),
            .in1(N__25628),
            .in2(_gnd_net_),
            .in3(N__25622),
            .lcout(clkdivZ0Z_18),
            .ltout(),
            .carryin(clkdiv_cry_17),
            .carryout(clkdiv_cry_18),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_19_LC_1_19_3.C_ON=1'b1;
    defparam clkdiv_19_LC_1_19_3.SEQ_MODE=4'b1000;
    defparam clkdiv_19_LC_1_19_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_19_LC_1_19_3 (
            .in0(_gnd_net_),
            .in1(N__25619),
            .in2(_gnd_net_),
            .in3(N__25613),
            .lcout(clkdivZ0Z_19),
            .ltout(),
            .carryin(clkdiv_cry_18),
            .carryout(clkdiv_cry_19),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_20_LC_1_19_4.C_ON=1'b1;
    defparam clkdiv_20_LC_1_19_4.SEQ_MODE=4'b1000;
    defparam clkdiv_20_LC_1_19_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_20_LC_1_19_4 (
            .in0(_gnd_net_),
            .in1(N__25610),
            .in2(_gnd_net_),
            .in3(N__25604),
            .lcout(clkdivZ0Z_20),
            .ltout(),
            .carryin(clkdiv_cry_19),
            .carryout(clkdiv_cry_20),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_21_LC_1_19_5.C_ON=1'b1;
    defparam clkdiv_21_LC_1_19_5.SEQ_MODE=4'b1000;
    defparam clkdiv_21_LC_1_19_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_21_LC_1_19_5 (
            .in0(_gnd_net_),
            .in1(N__25601),
            .in2(_gnd_net_),
            .in3(N__25595),
            .lcout(clkdivZ0Z_21),
            .ltout(),
            .carryin(clkdiv_cry_20),
            .carryout(clkdiv_cry_21),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_22_LC_1_19_6.C_ON=1'b1;
    defparam clkdiv_22_LC_1_19_6.SEQ_MODE=4'b1000;
    defparam clkdiv_22_LC_1_19_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_22_LC_1_19_6 (
            .in0(_gnd_net_),
            .in1(N__25592),
            .in2(_gnd_net_),
            .in3(N__25586),
            .lcout(clkdivZ0Z_22),
            .ltout(),
            .carryin(clkdiv_cry_21),
            .carryout(clkdiv_cry_22),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_23_LC_1_19_7.C_ON=1'b0;
    defparam clkdiv_23_LC_1_19_7.SEQ_MODE=4'b1000;
    defparam clkdiv_23_LC_1_19_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 clkdiv_23_LC_1_19_7 (
            .in0(_gnd_net_),
            .in1(N__25804),
            .in2(_gnd_net_),
            .in3(N__25814),
            .lcout(GPIO3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73293),
            .ce(),
            .sr(_gnd_net_));
    defparam \GPU.BUFFER.B_OE_c_i_LC_1_20_4 .C_ON=1'b0;
    defparam \GPU.BUFFER.B_OE_c_i_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \GPU.BUFFER.B_OE_c_i_LC_1_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \GPU.BUFFER.B_OE_c_i_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25765),
            .lcout(B_OE_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \GPU.BUFFER.OE_LC_3_20_4 .C_ON=1'b0;
    defparam \GPU.BUFFER.OE_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \GPU.BUFFER.OE_LC_3_20_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \GPU.BUFFER.OE_LC_3_20_4  (
            .in0(N__29474),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73304),
            .lcout(B_OE_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_11_LC_5_20_3 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_11_LC_5_20_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_11_LC_5_20_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.gpuAddReg_11_LC_5_20_3  (
            .in0(N__31234),
            .in1(N__70795),
            .in2(N__58004),
            .in3(N__70552),
            .lcout(gpuAddress_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_11C_net ),
            .ce(N__30760),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_14_LC_7_18_5 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_14_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_14_LC_7_18_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.gpuAddReg_14_LC_7_18_5  (
            .in0(N__31411),
            .in1(N__70794),
            .in2(N__57869),
            .in3(N__70548),
            .lcout(gpuAddress_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_14C_net ),
            .ce(N__30761),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_25dflt_LC_7_19_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_25dflt_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_25dflt_LC_7_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PROM.ROMDATA.dintern_25dflt_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__72376),
            .in2(_gnd_net_),
            .in3(N__72248),
            .lcout(controlWord_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_9_LC_7_20_0 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_9_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_9_LC_7_20_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.gpuAddReg_9_LC_7_20_0  (
            .in0(N__31123),
            .in1(N__70761),
            .in2(N__37970),
            .in3(N__70535),
            .lcout(gpuAddress_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_9C_net ),
            .ce(N__30752),
            .sr(_gnd_net_));
    defparam \RAM.OE_i_LC_7_23_2 .C_ON=1'b0;
    defparam \RAM.OE_i_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \RAM.OE_i_LC_7_23_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \RAM.OE_i_LC_7_23_2  (
            .in0(N__73302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34989),
            .lcout(N_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RAM.un1_WR_i_LC_7_23_6 .C_ON=1'b0;
    defparam \RAM.un1_WR_i_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \RAM.un1_WR_i_LC_7_23_6 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \RAM.un1_WR_i_LC_7_23_6  (
            .in0(N__73303),
            .in1(N__34990),
            .in2(N__29387),
            .in3(N__28148),
            .lcout(RAM_un1_WR_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_1_c_LC_9_9_0 .C_ON=1'b1;
    defparam \ALU.status_17_I_1_c_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_1_c_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_1_c_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__28598),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\ALU.status_17_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_9_c_LC_9_9_1 .C_ON=1'b1;
    defparam \ALU.status_17_I_9_c_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_9_c_LC_9_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_9_c_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__32464),
            .in2(N__27683),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_17_data_tmp_0 ),
            .carryout(\ALU.status_17_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_15_c_LC_9_9_2 .C_ON=1'b1;
    defparam \ALU.status_17_I_15_c_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_15_c_LC_9_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_15_c_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__26777),
            .in2(N__32479),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_17_data_tmp_1 ),
            .carryout(\ALU.status_17_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_27_c_LC_9_9_3 .C_ON=1'b1;
    defparam \ALU.status_17_I_27_c_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_27_c_LC_9_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_27_c_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__32456),
            .in2(N__25835),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_17_data_tmp_2 ),
            .carryout(\ALU.status_17_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_45_c_LC_9_9_4 .C_ON=1'b1;
    defparam \ALU.status_17_I_45_c_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_45_c_LC_9_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_45_c_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__25847),
            .in2(N__32481),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_17_data_tmp_3 ),
            .carryout(\ALU.status_17_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_33_c_LC_9_9_5 .C_ON=1'b1;
    defparam \ALU.status_17_I_33_c_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_33_c_LC_9_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_33_c_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__32457),
            .in2(N__26828),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_17_data_tmp_4 ),
            .carryout(\ALU.status_17_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_39_c_LC_9_9_6 .C_ON=1'b1;
    defparam \ALU.status_17_I_39_c_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_39_c_LC_9_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_39_c_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__37403),
            .in2(N__32480),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_17_data_tmp_5 ),
            .carryout(\ALU.status_17_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_21_c_LC_9_9_7 .C_ON=1'b1;
    defparam \ALU.status_17_I_21_c_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_21_c_LC_9_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_17_I_21_c_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__53030),
            .in2(N__32482),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_17_data_tmp_6 ),
            .carryout(\ALU.status_17_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_0_3_LC_9_10_0 .C_ON=1'b0;
    defparam \ALU.status_0_3_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.status_0_3_LC_9_10_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.status_0_3_LC_9_10_0  (
            .in0(N__69529),
            .in1(N__45448),
            .in2(N__56627),
            .in3(N__25817),
            .lcout(aluStatus_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73166),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_45_c_RNO_LC_9_10_5 .C_ON=1'b0;
    defparam \ALU.status_17_I_45_c_RNO_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_45_c_RNO_LC_9_10_5 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \ALU.status_17_I_45_c_RNO_LC_9_10_5  (
            .in0(N__61935),
            .in1(N__62890),
            .in2(N__62956),
            .in3(N__55817),
            .lcout(\ALU.status_17_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_0_c_LC_9_11_0 .C_ON=1'b1;
    defparam \ALU.status_18_cry_0_c_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_0_c_LC_9_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_0_c_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__60617),
            .in2(N__35324),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\ALU.status_18_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_1_c_inv_LC_9_11_1 .C_ON=1'b1;
    defparam \ALU.status_18_cry_1_c_inv_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_1_c_inv_LC_9_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_18_cry_1_c_inv_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__25841),
            .in2(N__65574),
            .in3(N__66048),
            .lcout(\ALU.combOperand2_i_1 ),
            .ltout(),
            .carryin(\ALU.status_18_cry_0 ),
            .carryout(\ALU.status_18_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_2_c_LC_9_11_2 .C_ON=1'b1;
    defparam \ALU.status_18_cry_2_c_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_2_c_LC_9_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_2_c_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__66313),
            .in2(N__32378),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_1 ),
            .carryout(\ALU.status_18_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_3_c_LC_9_11_3 .C_ON=1'b1;
    defparam \ALU.status_18_cry_3_c_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_3_c_LC_9_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_3_c_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__60261),
            .in2(N__27044),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_2 ),
            .carryout(\ALU.status_18_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_4_c_LC_9_11_4 .C_ON=1'b1;
    defparam \ALU.status_18_cry_4_c_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_4_c_LC_9_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_4_c_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__59873),
            .in2(N__26861),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_3 ),
            .carryout(\ALU.status_18_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_5_c_LC_9_11_5 .C_ON=1'b1;
    defparam \ALU.status_18_cry_5_c_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_5_c_LC_9_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_5_c_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__59503),
            .in2(N__34016),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_4 ),
            .carryout(\ALU.status_18_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_27_c_RNO_LC_9_11_6 .C_ON=1'b1;
    defparam \ALU.status_17_I_27_c_RNO_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_27_c_RNO_LC_9_11_6 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \ALU.status_17_I_27_c_RNO_LC_9_11_6  (
            .in0(N__55993),
            .in1(N__26813),
            .in2(N__62579),
            .in3(N__62186),
            .lcout(\ALU.status_17_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(\ALU.status_18_cry_5 ),
            .carryout(\ALU.status_18_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_7_c_inv_LC_9_11_7 .C_ON=1'b1;
    defparam \ALU.status_18_cry_7_c_inv_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_7_c_inv_LC_9_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_18_cry_7_c_inv_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__25823),
            .in2(N__62234),
            .in3(N__55992),
            .lcout(\ALU.combOperand2_i_7 ),
            .ltout(),
            .carryin(\ALU.status_18_cry_6 ),
            .carryout(\ALU.status_18_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_8_c_LC_9_12_0 .C_ON=1'b1;
    defparam \ALU.status_18_cry_8_c_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_8_c_LC_9_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_8_c_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__61947),
            .in2(N__26045),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\ALU.status_18_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_9_c_LC_9_12_1 .C_ON=1'b1;
    defparam \ALU.status_18_cry_9_c_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_9_c_LC_9_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_9_c_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__62891),
            .in2(N__62957),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_8 ),
            .carryout(\ALU.status_18_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_10_c_LC_9_12_2 .C_ON=1'b1;
    defparam \ALU.status_18_cry_10_c_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_10_c_LC_9_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_10_c_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__61681),
            .in2(N__25982),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_9 ),
            .carryout(\ALU.status_18_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_11_c_inv_LC_9_12_3 .C_ON=1'b1;
    defparam \ALU.status_18_cry_11_c_inv_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_11_c_inv_LC_9_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_18_cry_11_c_inv_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__61433),
            .in2(N__25877),
            .in3(N__57031),
            .lcout(\ALU.combOperand2_i_11 ),
            .ltout(),
            .carryin(\ALU.status_18_cry_10 ),
            .carryout(\ALU.status_18_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_12_c_LC_9_12_4 .C_ON=1'b1;
    defparam \ALU.status_18_cry_12_c_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_12_c_LC_9_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_12_c_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__61193),
            .in2(N__25997),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_11 ),
            .carryout(\ALU.status_18_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_13_c_LC_9_12_5 .C_ON=1'b1;
    defparam \ALU.status_18_cry_13_c_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_13_c_LC_9_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.status_18_cry_13_c_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__60995),
            .in2(N__25973),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALU.status_18_cry_12 ),
            .carryout(\ALU.status_18_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_14_c_inv_LC_9_12_6 .C_ON=1'b1;
    defparam \ALU.status_18_cry_14_c_inv_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_14_c_inv_LC_9_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_18_cry_14_c_inv_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__63847),
            .in2(N__25868),
            .in3(N__56753),
            .lcout(\ALU.combOperand2_i_14 ),
            .ltout(),
            .carryin(\ALU.status_18_cry_13 ),
            .carryout(\ALU.status_18_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_15_c_inv_LC_9_12_7 .C_ON=1'b1;
    defparam \ALU.status_18_cry_15_c_inv_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_15_c_inv_LC_9_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_18_cry_15_c_inv_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__63674),
            .in2(N__25859),
            .in3(N__74608),
            .lcout(\ALU.combOperand2_i_15 ),
            .ltout(),
            .carryin(\ALU.status_18_cry_14 ),
            .carryout(\ALU.status_18_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_4_LC_9_13_0 .C_ON=1'b0;
    defparam \ALU.status_4_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \ALU.status_4_LC_9_13_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.status_4_LC_9_13_0  (
            .in0(N__69530),
            .in1(N__40729),
            .in2(N__56623),
            .in3(N__25850),
            .lcout(aluStatus_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73194),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_10_c_RNO_LC_9_13_2 .C_ON=1'b0;
    defparam \ALU.status_18_cry_10_c_RNO_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_10_c_RNO_LC_9_13_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \ALU.status_18_cry_10_c_RNO_LC_9_13_2  (
            .in0(N__61682),
            .in1(N__71452),
            .in2(N__26906),
            .in3(N__37120),
            .lcout(\ALU.status_18_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3D2O61_2_LC_9_13_3 .C_ON=1'b0;
    defparam \ALU.d_RNI3D2O61_2_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3D2O61_2_LC_9_13_3 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.d_RNI3D2O61_2_LC_9_13_3  (
            .in0(N__56900),
            .in1(N__60246),
            .in2(N__56824),
            .in3(N__66292),
            .lcout(\ALU.d_RNI3D2O61Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_13_c_RNO_LC_9_13_6 .C_ON=1'b0;
    defparam \ALU.status_18_cry_13_c_RNO_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_13_c_RNO_LC_9_13_6 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \ALU.status_18_cry_13_c_RNO_LC_9_13_6  (
            .in0(N__39674),
            .in1(N__39651),
            .in2(N__61013),
            .in3(N__71453),
            .lcout(\ALU.status_18_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIG7366_2_LC_9_14_0 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIG7366_2_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIG7366_2_LC_9_14_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \CONTROL.busState_1_RNIG7366_2_LC_9_14_0  (
            .in0(N__50225),
            .in1(N__59587),
            .in2(N__25886),
            .in3(N__49596),
            .lcout(),
            .ltout(\CONTROL.busState_1_RNIG7366Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI3G078_0_LC_9_14_1 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI3G078_0_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI3G078_0_LC_9_14_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \CONTROL.busState_1_RNI3G078_0_LC_9_14_1  (
            .in0(N__25961),
            .in1(_gnd_net_),
            .in2(N__25964),
            .in3(N__49829),
            .lcout(bus_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI1JVK1_0_2_LC_9_14_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI1JVK1_0_2_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI1JVK1_0_2_LC_9_14_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \CONTROL.busState_1_RNI1JVK1_0_2_LC_9_14_2  (
            .in0(N__50224),
            .in1(N__25928),
            .in2(N__25922),
            .in3(N__49595),
            .lcout(\CONTROL.busState_1_RNI1JVK1_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI6MOJ_5_LC_9_14_3 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI6MOJ_5_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI6MOJ_5_LC_9_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNI6MOJ_5_LC_9_14_3  (
            .in0(N__25955),
            .in1(N__45673),
            .in2(_gnd_net_),
            .in3(N__50222),
            .lcout(\CONTROL.N_166 ),
            .ltout(\CONTROL.N_166_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI1JVK1_2_LC_9_14_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI1JVK1_2_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI1JVK1_2_LC_9_14_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \CONTROL.busState_1_RNI1JVK1_2_LC_9_14_4  (
            .in0(N__50223),
            .in1(N__25921),
            .in2(N__25889),
            .in3(N__49594),
            .lcout(N_182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI6OIF1_1_LC_9_14_5 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI6OIF1_1_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI6OIF1_1_LC_9_14_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI6OIF1_1_LC_9_14_5  (
            .in0(N__28920),
            .in1(N__27905),
            .in2(N__26996),
            .in3(N__27962),
            .lcout(romOut_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_5_LC_9_14_6 .C_ON=1'b0;
    defparam \CONTROL.dout_5_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_5_LC_9_14_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \CONTROL.dout_5_LC_9_14_6  (
            .in0(N__40912),
            .in1(N__50620),
            .in2(N__79532),
            .in3(N__38801),
            .lcout(\CONTROL.ctrlOut_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_5C_net ),
            .ce(N__44461),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_21dflt_LC_9_14_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_21dflt_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_21dflt_LC_9_14_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_21dflt_LC_9_14_7  (
            .in0(N__38800),
            .in1(N__79523),
            .in2(N__50621),
            .in3(N__40911),
            .lcout(controlWord_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1C0D5_12_LC_9_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNI1C0D5_12_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1C0D5_12_LC_9_15_0 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \ALU.d_RNI1C0D5_12_LC_9_15_0  (
            .in0(N__53967),
            .in1(N__26921),
            .in2(N__26015),
            .in3(N__26021),
            .lcout(\ALU.operand2_12 ),
            .ltout(\ALU.operand2_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0UD4G_12_LC_9_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNI0UD4G_12_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0UD4G_12_LC_9_15_1 .LUT_INIT=16'b0011001111110000;
    LogicCell40 \ALU.d_RNI0UD4G_12_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__31755),
            .in2(N__26030),
            .in3(N__71449),
            .lcout(\ALU.N_126 ),
            .ltout(\ALU.N_126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9UI0K_1_LC_9_15_2 .C_ON=1'b0;
    defparam \ALU.d_RNI9UI0K_1_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9UI0K_1_LC_9_15_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNI9UI0K_1_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26027),
            .in3(N__65563),
            .lcout(\ALU.d_RNI9UI0KZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8I8I5_0_10_LC_9_15_3 .C_ON=1'b0;
    defparam \ALU.d_RNI8I8I5_0_10_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8I8I5_0_10_LC_9_15_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ALU.d_RNI8I8I5_0_10_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__26895),
            .in2(_gnd_net_),
            .in3(N__71450),
            .lcout(\ALU.log_1_3cf0_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI670L_12_LC_9_15_4 .C_ON=1'b0;
    defparam \ALU.c_RNI670L_12_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI670L_12_LC_9_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNI670L_12_LC_9_15_4  (
            .in0(N__52411),
            .in1(N__67556),
            .in2(_gnd_net_),
            .in3(N__43307),
            .lcout(),
            .ltout(\ALU.c_RNI670LZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIHJ2L2_12_LC_9_15_5 .C_ON=1'b0;
    defparam \ALU.c_RNIHJ2L2_12_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIHJ2L2_12_LC_9_15_5 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \ALU.c_RNIHJ2L2_12_LC_9_15_5  (
            .in0(N__46841),
            .in1(N__53966),
            .in2(N__26024),
            .in3(N__28952),
            .lcout(\ALU.operand2_7_ns_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8FCT_12_LC_9_15_6 .C_ON=1'b0;
    defparam \ALU.d_RNI8FCT_12_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8FCT_12_LC_9_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNI8FCT_12_LC_9_15_6  (
            .in0(N__57946),
            .in1(N__65096),
            .in2(_gnd_net_),
            .in3(N__43308),
            .lcout(\ALU.d_RNI8FCTZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_12_c_RNO_LC_9_15_7 .C_ON=1'b0;
    defparam \ALU.status_18_cry_12_c_RNO_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_12_c_RNO_LC_9_15_7 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \ALU.status_18_cry_12_c_RNO_LC_9_15_7  (
            .in0(N__61199),
            .in1(N__31756),
            .in2(N__26006),
            .in3(N__71451),
            .lcout(\ALU.status_18_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIIBVU9_10_LC_9_16_0 .C_ON=1'b0;
    defparam \ALU.c_RNIIBVU9_10_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIIBVU9_10_LC_9_16_0 .LUT_INIT=16'b1100101110010010;
    LogicCell40 \ALU.c_RNIIBVU9_10_LC_9_16_0  (
            .in0(N__63247),
            .in1(N__26069),
            .in2(N__74889),
            .in3(N__61662),
            .lcout(),
            .ltout(\ALU.log_1_3cf0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJPU5U_10_LC_9_16_1 .C_ON=1'b0;
    defparam \ALU.c_RNIJPU5U_10_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJPU5U_10_LC_9_16_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.c_RNIJPU5U_10_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__26060),
            .in2(N__26063),
            .in3(N__37113),
            .lcout(\ALU.log_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIIBVU9_0_10_LC_9_16_2 .C_ON=1'b0;
    defparam \ALU.c_RNIIBVU9_0_10_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIIBVU9_0_10_LC_9_16_2 .LUT_INIT=16'b0011111001101000;
    LogicCell40 \ALU.c_RNIIBVU9_0_10_LC_9_16_2  (
            .in0(N__63246),
            .in1(N__26054),
            .in2(N__74888),
            .in3(N__61661),
            .lcout(\ALU.log_1_3cf1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8I8I5_10_LC_9_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNI8I8I5_10_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8I8I5_10_LC_9_16_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ALU.d_RNI8I8I5_10_LC_9_16_3  (
            .in0(N__71424),
            .in1(_gnd_net_),
            .in2(N__26905),
            .in3(_gnd_net_),
            .lcout(\ALU.log_1_3cf1_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIMSAK1_0_LC_9_16_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIMSAK1_0_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIMSAK1_0_LC_9_16_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \CONTROL.busState_1_RNIMSAK1_0_LC_9_16_4  (
            .in0(N__49587),
            .in1(N__50298),
            .in2(N__49824),
            .in3(N__50190),
            .lcout(\CONTROL.bus_7_a0_2_8 ),
            .ltout(\CONTROL.bus_7_a0_2_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIF208A_0_0_LC_9_16_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIF208A_0_0_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIF208A_0_0_LC_9_16_5 .LUT_INIT=16'b0011111100000000;
    LogicCell40 \CONTROL.busState_1_RNIF208A_0_0_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__27194),
            .in2(N__26048),
            .in3(N__29056),
            .lcout(bus_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_8_c_RNO_LC_9_16_6 .C_ON=1'b0;
    defparam \ALU.status_18_cry_8_c_RNO_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_8_c_RNO_LC_9_16_6 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \ALU.status_18_cry_8_c_RNO_LC_9_16_6  (
            .in0(N__57094),
            .in1(N__26957),
            .in2(N__61948),
            .in3(N__71425),
            .lcout(\ALU.status_18_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIA8EO_0_LC_9_17_1 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIA8EO_0_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIA8EO_0_LC_9_17_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIA8EO_0_LC_9_17_1  (
            .in0(N__32308),
            .in1(N__26075),
            .in2(_gnd_net_),
            .in3(N__26092),
            .lcout(DROM_ROMDATA_dintern_8ro),
            .ltout(DROM_ROMDATA_dintern_8ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI05PC2_0_LC_9_17_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI05PC2_0_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI05PC2_0_LC_9_17_2 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \CONTROL.busState_1_RNI05PC2_0_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26033),
            .in3(N__27268),
            .lcout(busState_1_RNI05PC2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIA6749_0_LC_9_17_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIA6749_0_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIA6749_0_LC_9_17_3 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \CONTROL.busState_1_RNIA6749_0_LC_9_17_3  (
            .in0(N__27269),
            .in1(N__26146),
            .in2(_gnd_net_),
            .in3(N__29120),
            .lcout(bus_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIA6749_0_0_LC_9_17_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIA6749_0_0_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIA6749_0_0_LC_9_17_5 .LUT_INIT=16'b1000111110001111;
    LogicCell40 \CONTROL.busState_1_RNIA6749_0_0_LC_9_17_5  (
            .in0(N__27270),
            .in1(N__26147),
            .in2(N__27842),
            .in3(_gnd_net_),
            .lcout(bus_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI7LJL_1_LC_9_17_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI7LJL_1_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI7LJL_1_LC_9_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI7LJL_1_LC_9_17_6  (
            .in0(N__26099),
            .in1(N__26107),
            .in2(_gnd_net_),
            .in3(N__32307),
            .lcout(DROM_ROMDATA_dintern_1ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_1_LC_9_17_7 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_1_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_1_LC_9_17_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_1_LC_9_17_7  (
            .in0(N__26108),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C_net ),
            .ce(N__32324),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_1_LC_9_18_0 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_1_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_1_LC_9_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_1_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27068),
            .lcout(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net ),
            .ce(N__32321),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_2_LC_9_18_1 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_2_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_2_LC_9_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_2_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26273),
            .lcout(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net ),
            .ce(N__32321),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_3_LC_9_18_2 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_3_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_3_LC_9_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_3_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26246),
            .lcout(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net ),
            .ce(N__32321),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_0_LC_9_18_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_0_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_0_LC_9_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_0_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26093),
            .lcout(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net ),
            .ce(N__32321),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNICIR11_0_LC_9_19_0 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNICIR11_0_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNICIR11_0_LC_9_19_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_RNICIR11_0_LC_9_19_0  (
            .in0(N__27353),
            .in1(N__27376),
            .in2(_gnd_net_),
            .in3(N__32302),
            .lcout(DROM_ROMDATA_dintern_12ro),
            .ltout(DROM_ROMDATA_dintern_12ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI8R4IA_0_0_LC_9_19_1 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI8R4IA_0_0_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI8R4IA_0_0_LC_9_19_1 .LUT_INIT=16'b0000110011001100;
    LogicCell40 \CONTROL.busState_1_RNI8R4IA_0_0_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__30541),
            .in2(N__26336),
            .in3(N__27283),
            .lcout(bus_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_3_LC_9_19_2 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_3_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_3_LC_9_19_2 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \CONTROL.aluOperation_3_LC_9_19_2  (
            .in0(N__36689),
            .in1(N__69766),
            .in2(N__38140),
            .in3(N__41504),
            .lcout(aluOperation_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluOperation_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI8R4IA_0_LC_9_19_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI8R4IA_0_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI8R4IA_0_LC_9_19_3 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \CONTROL.busState_1_RNI8R4IA_0_LC_9_19_3  (
            .in0(N__26333),
            .in1(N__30542),
            .in2(_gnd_net_),
            .in3(N__27284),
            .lcout(bus_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIDBEO_3_LC_9_19_4 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIDBEO_3_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIDBEO_3_LC_9_19_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIDBEO_3_LC_9_19_4  (
            .in0(N__27383),
            .in1(N__27400),
            .in2(_gnd_net_),
            .in3(N__32300),
            .lcout(DROM_ROMDATA_dintern_11ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIEKR11_2_LC_9_19_5 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIEKR11_2_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIEKR11_2_LC_9_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIEKR11_2_LC_9_19_5  (
            .in0(N__32301),
            .in1(N__26279),
            .in2(_gnd_net_),
            .in3(N__26269),
            .lcout(DROM_ROMDATA_dintern_14ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIFLR11_3_LC_9_19_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIFLR11_3_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIFLR11_3_LC_9_19_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIFLR11_3_LC_9_19_6  (
            .in0(N__26252),
            .in1(N__26245),
            .in2(_gnd_net_),
            .in3(N__32303),
            .lcout(DROM_ROMDATA_dintern_15ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIF208A_0_LC_9_19_7 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIF208A_0_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIF208A_0_LC_9_19_7 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \CONTROL.busState_1_RNIF208A_0_LC_9_19_7  (
            .in0(N__29057),
            .in1(N__27193),
            .in2(_gnd_net_),
            .in3(N__27285),
            .lcout(bus_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_0_LC_9_20_0 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_0_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_0_LC_9_20_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \CONTROL.gpuAddReg_0_LC_9_20_0  (
            .in0(N__33317),
            .in1(N__70785),
            .in2(N__70544),
            .in3(N__37565),
            .lcout(gpuAddress_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_0C_net ),
            .ce(N__30739),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_1_LC_9_20_1 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_1_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_1_LC_9_20_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \CONTROL.gpuAddReg_1_LC_9_20_1  (
            .in0(N__70541),
            .in1(N__37520),
            .in2(N__70798),
            .in3(N__33257),
            .lcout(gpuAddress_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_0C_net ),
            .ce(N__30739),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_10_LC_9_20_2 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_10_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_10_LC_9_20_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.gpuAddReg_10_LC_9_20_2  (
            .in0(N__31276),
            .in1(N__70542),
            .in2(N__58241),
            .in3(N__70786),
            .lcout(gpuAddress_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_0C_net ),
            .ce(N__30739),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_12_LC_9_20_4 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_12_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_12_LC_9_20_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.gpuAddReg_12_LC_9_20_4  (
            .in0(N__57950),
            .in1(N__70543),
            .in2(N__28229),
            .in3(N__70787),
            .lcout(gpuAddress_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_0C_net ),
            .ce(N__30739),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_13_LC_9_20_5 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_13_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_13_LC_9_20_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \CONTROL.gpuAddReg_13_LC_9_20_5  (
            .in0(N__70539),
            .in1(N__27988),
            .in2(N__70796),
            .in3(N__57908),
            .lcout(gpuAddress_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_0C_net ),
            .ce(N__30739),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_15_LC_9_20_7 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_15_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_15_LC_9_20_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \CONTROL.gpuAddReg_15_LC_9_20_7  (
            .in0(N__70540),
            .in1(N__54194),
            .in2(N__70797),
            .in3(N__45010),
            .lcout(gpuAddress_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_0C_net ),
            .ce(N__30739),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_2_LC_9_21_0 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_2_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_2_LC_9_21_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.romAddReg_7_2_LC_9_21_0  (
            .in0(N__29596),
            .in1(N__72212),
            .in2(N__35570),
            .in3(N__71822),
            .lcout(CONTROL_romAddReg_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_3_LC_9_21_1 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_3_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_3_LC_9_21_1 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \CONTROL.romAddReg_7_3_LC_9_21_1  (
            .in0(N__71825),
            .in1(N__37745),
            .in2(N__72289),
            .in3(N__44278),
            .lcout(CONTROL_romAddReg_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_3_LC_9_21_2 .C_ON=1'b0;
    defparam \CONTROL.dout_3_LC_9_21_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_3_LC_9_21_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \CONTROL.dout_3_LC_9_21_2  (
            .in0(N__44279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__72220),
            .lcout(\CONTROL.ctrlOut_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_3C_net ),
            .ce(N__44462),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_5_LC_9_21_4 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_5_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_5_LC_9_21_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.romAddReg_7_5_LC_9_21_4  (
            .in0(N__40148),
            .in1(N__72213),
            .in2(N__29451),
            .in3(N__71823),
            .lcout(CONTROL_romAddReg_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m461_ns_LC_9_21_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m461_ns_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m461_ns_LC_9_21_5 .LUT_INIT=16'b1101000100010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m461_ns_LC_9_21_5  (
            .in0(N__47762),
            .in1(N__72773),
            .in2(N__55505),
            .in3(N__74072),
            .lcout(PROM_ROMDATA_dintern_23ro),
            .ltout(PROM_ROMDATA_dintern_23ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_7_LC_9_21_6 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_7_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_7_LC_9_21_6 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \CONTROL.romAddReg_7_7_LC_9_21_6  (
            .in0(N__72247),
            .in1(N__48872),
            .in2(N__26642),
            .in3(N__71824),
            .lcout(CONTROL_romAddReg_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_6_LC_9_21_7 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_6_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_6_LC_9_21_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \CONTROL.romAddReg_7_6_LC_9_21_7  (
            .in0(N__71826),
            .in1(N__35760),
            .in2(N__72288),
            .in3(N__70815),
            .lcout(CONTROL_romAddReg_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m465_bm_LC_9_22_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m465_bm_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m465_bm_LC_9_22_0 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m465_bm_LC_9_22_0  (
            .in0(N__64022),
            .in1(N__76625),
            .in2(N__65033),
            .in3(N__76015),
            .lcout(),
            .ltout(\PROM.ROMDATA.m465_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m471_ns_1_LC_9_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m471_ns_1_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m471_ns_1_LC_9_22_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m471_ns_1_LC_9_22_1  (
            .in0(N__33416),
            .in1(N__79500),
            .in2(N__26576),
            .in3(N__79896),
            .lcout(),
            .ltout(\PROM.ROMDATA.m471_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m471_ns_LC_9_22_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m471_ns_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m471_ns_LC_9_22_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m471_ns_LC_9_22_2  (
            .in0(N__79501),
            .in1(N__40985),
            .in2(N__26573),
            .in3(N__29615),
            .lcout(\PROM.ROMDATA.m471_ns ),
            .ltout(\PROM.ROMDATA.m471_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_24dflt_LC_9_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_24dflt_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_24dflt_LC_9_22_3 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_24dflt_LC_9_22_3  (
            .in0(N__47494),
            .in1(N__72774),
            .in2(N__26570),
            .in3(N__72221),
            .lcout(controlWord_24),
            .ltout(controlWord_24_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_8_LC_9_22_4 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_8_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_8_LC_9_22_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \CONTROL.romAddReg_7_8_LC_9_22_4  (
            .in0(N__71873),
            .in1(N__72223),
            .in2(N__26567),
            .in3(N__50438),
            .lcout(CONTROL_romAddReg_7_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_4_LC_9_22_7 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_4_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_4_LC_9_22_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.romAddReg_7_4_LC_9_22_7  (
            .in0(N__44178),
            .in1(N__72222),
            .in2(N__35807),
            .in3(N__71874),
            .lcout(CONTROL_romAddReg_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI2UPI1_5_LC_9_23_0 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI2UPI1_5_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI2UPI1_5_LC_9_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI2UPI1_5_LC_9_23_0  (
            .in0(N__34769),
            .in1(N__57819),
            .in2(N__60735),
            .in3(N__27499),
            .lcout(),
            .ltout(\CONTROL.g0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI6P3NN91_4_LC_9_23_1 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI6P3NN91_4_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI6P3NN91_4_LC_9_23_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI6P3NN91_4_LC_9_23_1  (
            .in0(N__38443),
            .in1(N__60813),
            .in2(N__26696),
            .in3(N__41986),
            .lcout(\CONTROL.addrstackptr_N_10_mux_0_0_0 ),
            .ltout(\CONTROL.addrstackptr_N_10_mux_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNIEKK1Q82_6_LC_9_23_2 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNIEKK1Q82_6_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNIEKK1Q82_6_LC_9_23_2 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \CONTROL.addrstackptr_RNIEKK1Q82_6_LC_9_23_2  (
            .in0(N__26750),
            .in1(N__26725),
            .in2(N__26693),
            .in3(N__26672),
            .lcout(\CONTROL.addrstackptr_N_7_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_19_LC_9_23_3 .C_ON=1'b0;
    defparam \CONTROL.g0_19_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_19_LC_9_23_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CONTROL.g0_19_LC_9_23_3  (
            .in0(N__36470),
            .in1(N__42261),
            .in2(N__45368),
            .in3(N__38184),
            .lcout(),
            .ltout(\CONTROL.N_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIDB191V_7_LC_9_23_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIDB191V_7_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIDB191V_7_LC_9_23_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIDB191V_7_LC_9_23_4  (
            .in0(N__38516),
            .in1(N__42044),
            .in2(N__26675),
            .in3(N__41503),
            .lcout(\CONTROL.N_4_2 ),
            .ltout(\CONTROL.N_4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_6_LC_9_23_5 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_6_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_6_LC_9_23_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \CONTROL.addrstackptr_6_LC_9_23_5  (
            .in0(N__26726),
            .in1(N__26751),
            .in2(N__26666),
            .in3(N__26663),
            .lcout(\CONTROL.addrstackptrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.addrstackptr_6C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI73QI1_6_LC_9_23_6 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI73QI1_6_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI73QI1_6_LC_9_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI73QI1_6_LC_9_23_6  (
            .in0(N__34770),
            .in1(N__27498),
            .in2(N__26753),
            .in3(N__38442),
            .lcout(\CONTROL.g1_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_13_LC_9_24_1 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_13_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_13_LC_9_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_13_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28343),
            .lcout(\CONTROL.tempCounterZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_13C_net ),
            .ce(N__34970),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_6_LC_9_24_2 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_6_LC_9_24_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_6_LC_9_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_6_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47839),
            .lcout(\CONTROL.tempCounterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_13C_net ),
            .ce(N__34970),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_0_c_LC_9_25_0 .C_ON=1'b1;
    defparam \CONTROL.addrstack_1_cry_0_c_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_0_c_LC_9_25_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \CONTROL.addrstack_1_cry_0_c_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(N__57791),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\CONTROL.addrstack_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_0_c_RNIDDJK_LC_9_25_1 .C_ON=1'b1;
    defparam \CONTROL.addrstack_1_cry_0_c_RNIDDJK_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_0_c_RNIDDJK_LC_9_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \CONTROL.addrstack_1_cry_0_c_RNIDDJK_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__38431),
            .in2(N__32567),
            .in3(N__26768),
            .lcout(\CONTROL.addrstack_1_1 ),
            .ltout(),
            .carryin(\CONTROL.addrstack_1_cry_0 ),
            .carryout(\CONTROL.addrstack_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_1_c_RNIFGKK_LC_9_25_2 .C_ON=1'b1;
    defparam \CONTROL.addrstack_1_cry_1_c_RNIFGKK_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_1_c_RNIFGKK_LC_9_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \CONTROL.addrstack_1_cry_1_c_RNIFGKK_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__32554),
            .in2(N__60734),
            .in3(N__26765),
            .lcout(\CONTROL.addrstack_1_2 ),
            .ltout(),
            .carryin(\CONTROL.addrstack_1_cry_1 ),
            .carryout(\CONTROL.addrstack_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_2_c_RNIHJLK_LC_9_25_3 .C_ON=1'b1;
    defparam \CONTROL.addrstack_1_cry_2_c_RNIHJLK_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_2_c_RNIHJLK_LC_9_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \CONTROL.addrstack_1_cry_2_c_RNIHJLK_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(N__34768),
            .in2(N__32568),
            .in3(N__26762),
            .lcout(\CONTROL.addrstack_1_3 ),
            .ltout(),
            .carryin(\CONTROL.addrstack_1_cry_2 ),
            .carryout(\CONTROL.addrstack_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_3_c_RNIJMMK_LC_9_25_4 .C_ON=1'b1;
    defparam \CONTROL.addrstack_1_cry_3_c_RNIJMMK_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_3_c_RNIJMMK_LC_9_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \CONTROL.addrstack_1_cry_3_c_RNIJMMK_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__32558),
            .in2(N__60812),
            .in3(N__26759),
            .lcout(\CONTROL.addrstack_1_4 ),
            .ltout(),
            .carryin(\CONTROL.addrstack_1_cry_3 ),
            .carryout(\CONTROL.addrstack_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_4_c_RNILPNK_LC_9_25_5 .C_ON=1'b1;
    defparam \CONTROL.addrstack_1_cry_4_c_RNILPNK_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_4_c_RNILPNK_LC_9_25_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \CONTROL.addrstack_1_cry_4_c_RNILPNK_LC_9_25_5  (
            .in0(_gnd_net_),
            .in1(N__27500),
            .in2(N__32569),
            .in3(N__26756),
            .lcout(\CONTROL.addrstack_1_5 ),
            .ltout(),
            .carryin(\CONTROL.addrstack_1_cry_4 ),
            .carryout(\CONTROL.addrstack_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_5_c_RNINSOK_LC_9_25_6 .C_ON=1'b1;
    defparam \CONTROL.addrstack_1_cry_5_c_RNINSOK_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_5_c_RNINSOK_LC_9_25_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \CONTROL.addrstack_1_cry_5_c_RNINSOK_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__32562),
            .in2(N__26752),
            .in3(N__26705),
            .lcout(\CONTROL.addrstack_1_6 ),
            .ltout(),
            .carryin(\CONTROL.addrstack_1_cry_5 ),
            .carryout(\CONTROL.addrstack_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_1_cry_6_c_RNIPVPK_LC_9_25_7 .C_ON=1'b0;
    defparam \CONTROL.addrstack_1_cry_6_c_RNIPVPK_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_1_cry_6_c_RNIPVPK_LC_9_25_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \CONTROL.addrstack_1_cry_6_c_RNIPVPK_LC_9_25_7  (
            .in0(_gnd_net_),
            .in1(N__42287),
            .in2(_gnd_net_),
            .in3(N__26702),
            .lcout(\CONTROL.addrstack_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI69B31_5_LC_10_10_0 .C_ON=1'b0;
    defparam \ALU.e_RNI69B31_5_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI69B31_5_LC_10_10_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNI69B31_5_LC_10_10_0  (
            .in0(N__40036),
            .in1(N__34568),
            .in2(N__40070),
            .in3(N__43931),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIE8D02_5_LC_10_10_1 .C_ON=1'b0;
    defparam \ALU.c_RNIE8D02_5_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIE8D02_5_LC_10_10_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNIE8D02_5_LC_10_10_1  (
            .in0(N__40144),
            .in1(N__40097),
            .in2(N__26699),
            .in3(N__47212),
            .lcout(\ALU.N_1090 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI8FH51_5_LC_10_10_2 .C_ON=1'b0;
    defparam \ALU.b_RNI8FH51_5_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI8FH51_5_LC_10_10_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI8FH51_5_LC_10_10_2  (
            .in0(N__39932),
            .in1(N__34567),
            .in2(N__39972),
            .in3(N__43930),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIKPK1_5_LC_10_10_3 .C_ON=1'b0;
    defparam \ALU.d_RNIIKPK1_5_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIKPK1_5_LC_10_10_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIIKPK1_5_LC_10_10_3  (
            .in0(N__40239),
            .in1(N__40220),
            .in2(N__26795),
            .in3(N__47213),
            .lcout(),
            .ltout(\ALU.N_1138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI31LU3_5_LC_10_10_4 .C_ON=1'b0;
    defparam \ALU.d_RNI31LU3_5_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI31LU3_5_LC_10_10_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNI31LU3_5_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__54143),
            .in2(N__26792),
            .in3(N__26789),
            .lcout(aluOut_5),
            .ltout(aluOut_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJRM75_5_LC_10_10_5 .C_ON=1'b0;
    defparam \ALU.d_RNIJRM75_5_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJRM75_5_LC_10_10_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.d_RNIJRM75_5_LC_10_10_5  (
            .in0(N__53289),
            .in1(N__49607),
            .in2(N__26783),
            .in3(N__50220),
            .lcout(\ALU.d_RNIJRM75Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILKJ1I_5_LC_10_11_0 .C_ON=1'b0;
    defparam \ALU.d_RNILKJ1I_5_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILKJ1I_5_LC_10_11_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNILKJ1I_5_LC_10_11_0  (
            .in0(N__59486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56077),
            .lcout(\ALU.d_RNILKJ1IZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIK31N31_10_LC_10_11_1 .C_ON=1'b0;
    defparam \ALU.c_RNIK31N31_10_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIK31N31_10_LC_10_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.c_RNIK31N31_10_LC_10_11_1  (
            .in0(N__61427),
            .in1(N__56377),
            .in2(N__68517),
            .in3(N__61667),
            .lcout(\ALU.c_RNIK31N31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7BDMH_7_LC_10_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNI7BDMH_7_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7BDMH_7_LC_10_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI7BDMH_7_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__62185),
            .in2(_gnd_net_),
            .in3(N__56078),
            .lcout(\ALU.d_RNI7BDMHZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILEAFE_5_LC_10_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNILEAFE_5_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILEAFE_5_LC_10_11_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \ALU.d_RNILEAFE_5_LC_10_11_3  (
            .in0(N__40585),
            .in1(N__28933),
            .in2(N__28921),
            .in3(N__28876),
            .lcout(\ALU.status_19_4 ),
            .ltout(\ALU.status_19_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI07V431_2_LC_10_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNI07V431_2_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI07V431_2_LC_10_11_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNI07V431_2_LC_10_11_4  (
            .in0(N__56378),
            .in1(N__60245),
            .in2(N__26780),
            .in3(N__66296),
            .lcout(\ALU.d_RNI07V431Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_15_c_RNO_LC_10_11_5 .C_ON=1'b0;
    defparam \ALU.status_17_I_15_c_RNO_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_15_c_RNO_LC_10_11_5 .LUT_INIT=16'b1110101111010111;
    LogicCell40 \ALU.status_17_I_15_c_RNO_LC_10_11_5  (
            .in0(N__34012),
            .in1(N__59881),
            .in2(N__26857),
            .in3(N__59487),
            .lcout(\ALU.status_17_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIUEFBI_1_LC_10_11_6 .C_ON=1'b0;
    defparam \ALU.d_RNIUEFBI_1_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIUEFBI_1_LC_10_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIUEFBI_1_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__65558),
            .in2(_gnd_net_),
            .in3(N__56196),
            .lcout(\ALU.d_RNIUEFBIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIALE3I_6_LC_10_12_0 .C_ON=1'b0;
    defparam \ALU.d_RNIALE3I_6_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIALE3I_6_LC_10_12_0 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \ALU.d_RNIALE3I_6_LC_10_12_0  (
            .in0(N__26812),
            .in1(_gnd_net_),
            .in2(N__63292),
            .in3(N__62506),
            .lcout(\ALU.d_RNIALE3IZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIJU2E_0_6_LC_10_12_1 .C_ON=1'b0;
    defparam \ALU.d_RNIIJU2E_0_6_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIJU2E_0_6_LC_10_12_1 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \ALU.d_RNIIJU2E_0_6_LC_10_12_1  (
            .in0(N__26933),
            .in1(N__27345),
            .in2(N__32693),
            .in3(N__40581),
            .lcout(\ALU.combOperand2_0_6 ),
            .ltout(\ALU.combOperand2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA9P4I_6_LC_10_12_2 .C_ON=1'b0;
    defparam \ALU.d_RNIA9P4I_6_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA9P4I_6_LC_10_12_2 .LUT_INIT=16'b1110001110000110;
    LogicCell40 \ALU.d_RNIA9P4I_6_LC_10_12_2  (
            .in0(N__63265),
            .in1(N__74890),
            .in2(N__26801),
            .in3(N__62505),
            .lcout(\ALU.N_22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI67HQ21_0_LC_10_12_3 .C_ON=1'b0;
    defparam \ALU.d_RNI67HQ21_0_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI67HQ21_0_LC_10_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI67HQ21_0_LC_10_12_3  (
            .in0(N__65545),
            .in1(N__60593),
            .in2(N__68506),
            .in3(N__56328),
            .lcout(\ALU.d_RNI67HQ21Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIJU2E_6_LC_10_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNIIJU2E_6_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIJU2E_6_LC_10_12_4 .LUT_INIT=16'b1110110011111111;
    LogicCell40 \ALU.d_RNIIJU2E_6_LC_10_12_4  (
            .in0(N__40580),
            .in1(N__32689),
            .in2(N__27347),
            .in3(N__26932),
            .lcout(\ALU.status_19_5 ),
            .ltout(\ALU.status_19_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5NE641_0_LC_10_12_5 .C_ON=1'b0;
    defparam \ALU.d_RNI5NE641_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5NE641_0_LC_10_12_5 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.d_RNI5NE641_0_LC_10_12_5  (
            .in0(N__65544),
            .in1(N__60594),
            .in2(N__26798),
            .in3(N__56223),
            .lcout(\ALU.d_RNI5NE641Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBLU321_6_LC_10_12_6 .C_ON=1'b0;
    defparam \ALU.d_RNIBLU321_6_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBLU321_6_LC_10_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIBLU321_6_LC_10_12_6  (
            .in0(N__55989),
            .in1(N__62504),
            .in2(N__62324),
            .in3(N__55801),
            .lcout(\ALU.d_RNIBLU321Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI73D441_6_LC_10_12_7 .C_ON=1'b0;
    defparam \ALU.d_RNI73D441_6_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI73D441_6_LC_10_12_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNI73D441_6_LC_10_12_7  (
            .in0(N__62503),
            .in1(N__56076),
            .in2(N__62316),
            .in3(N__56224),
            .lcout(\ALU.d_RNI73D441Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVPV6E_0_4_LC_10_13_0 .C_ON=1'b0;
    defparam \ALU.d_RNIVPV6E_0_4_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVPV6E_0_4_LC_10_13_0 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \ALU.d_RNIVPV6E_0_4_LC_10_13_0  (
            .in0(N__27755),
            .in1(N__26870),
            .in2(N__40592),
            .in3(N__28013),
            .lcout(\ALU.combOperand2_0_4 ),
            .ltout(\ALU.combOperand2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7BF7I_4_LC_10_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNI7BF7I_4_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7BF7I_4_LC_10_13_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \ALU.d_RNI7BF7I_4_LC_10_13_1  (
            .in0(N__59802),
            .in1(_gnd_net_),
            .in2(N__26876),
            .in3(N__63260),
            .lcout(\ALU.d_RNI7BF7IZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un14_log_a0_2_15_LC_10_13_2 .C_ON=1'b0;
    defparam \ALU.un14_log_a0_2_15_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un14_log_a0_2_15_LC_10_13_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ALU.un14_log_a0_2_15_LC_10_13_2  (
            .in0(N__50216),
            .in1(N__53232),
            .in2(N__49606),
            .in3(N__50327),
            .lcout(\ALU.un14_log_a0_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIU83C1_2_LC_10_13_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIU83C1_2_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIU83C1_2_LC_10_13_3 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \CONTROL.busState_1_RNIU83C1_2_LC_10_13_3  (
            .in0(N__37994),
            .in1(N__49600),
            .in2(N__33143),
            .in3(N__50217),
            .lcout(),
            .ltout(N_181_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVKK66_4_LC_10_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNIVKK66_4_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVKK66_4_LC_10_13_4 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \ALU.d_RNIVKK66_4_LC_10_13_4  (
            .in0(N__53233),
            .in1(N__71440),
            .in2(N__26873),
            .in3(N__27797),
            .lcout(\ALU.d_RNIVKK66Z0Z_4 ),
            .ltout(\ALU.d_RNIVKK66Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVPV6E_4_LC_10_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNIVPV6E_4_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVPV6E_4_LC_10_13_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \ALU.d_RNIVPV6E_4_LC_10_13_5  (
            .in0(N__28012),
            .in1(N__40576),
            .in2(N__26864),
            .in3(N__27754),
            .lcout(\ALU.status_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7VP8I_4_LC_10_13_6 .C_ON=1'b0;
    defparam \ALU.d_RNI7VP8I_4_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7VP8I_4_LC_10_13_6 .LUT_INIT=16'b1100101110010010;
    LogicCell40 \ALU.d_RNI7VP8I_4_LC_10_13_6  (
            .in0(N__63261),
            .in1(N__26844),
            .in2(N__74903),
            .in3(N__59801),
            .lcout(\ALU.log_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8JFO21_6_LC_10_14_0 .C_ON=1'b0;
    defparam \ALU.d_RNI8JFO21_6_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8JFO21_6_LC_10_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI8JFO21_6_LC_10_14_0  (
            .in0(N__68438),
            .in1(N__62502),
            .in2(N__62302),
            .in3(N__56345),
            .lcout(\ALU.d_RNI8JFO21Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_33_c_RNO_LC_10_14_1 .C_ON=1'b0;
    defparam \ALU.status_17_I_33_c_RNO_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_33_c_RNO_LC_10_14_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \ALU.status_17_I_33_c_RNO_LC_10_14_1  (
            .in0(N__57033),
            .in1(N__61463),
            .in2(N__61718),
            .in3(N__55549),
            .lcout(\ALU.status_17_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI1QK5K_10_LC_10_14_2 .C_ON=1'b0;
    defparam \ALU.c_RNI1QK5K_10_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI1QK5K_10_LC_10_14_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \ALU.c_RNI1QK5K_10_LC_10_14_2  (
            .in0(N__55548),
            .in1(_gnd_net_),
            .in2(N__63293),
            .in3(N__61714),
            .lcout(\ALU.c_RNI1QK5KZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIRRB4I_11_LC_10_14_3 .C_ON=1'b0;
    defparam \ALU.c_RNIRRB4I_11_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIRRB4I_11_LC_10_14_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ALU.c_RNIRRB4I_11_LC_10_14_3  (
            .in0(N__57032),
            .in1(N__63269),
            .in2(_gnd_net_),
            .in3(N__61464),
            .lcout(\ALU.c_RNIRRB4IZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC0VE6_5_LC_10_14_4 .C_ON=1'b0;
    defparam \ALU.d_RNIC0VE6_5_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC0VE6_5_LC_10_14_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.d_RNIC0VE6_5_LC_10_14_4  (
            .in0(N__71441),
            .in1(N__26939),
            .in2(N__53291),
            .in3(N__40001),
            .lcout(\ALU.d_RNIC0VE6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI18J1J_3_LC_10_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNI18J1J_3_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI18J1J_3_LC_10_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI18J1J_3_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__60219),
            .in2(_gnd_net_),
            .in3(N__55547),
            .lcout(\ALU.d_RNI18J1JZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKHEQH_7_LC_10_14_6 .C_ON=1'b0;
    defparam \ALU.d_RNIKHEQH_7_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKHEQH_7_LC_10_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIKHEQH_7_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__62274),
            .in2(_gnd_net_),
            .in3(N__56346),
            .lcout(\ALU.d_RNIKHEQHZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMCVI41_2_LC_10_14_7 .C_ON=1'b0;
    defparam \ALU.d_RNIMCVI41_2_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMCVI41_2_LC_10_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIMCVI41_2_LC_10_14_7  (
            .in0(N__60220),
            .in1(N__55546),
            .in2(N__55670),
            .in3(N__66299),
            .lcout(\ALU.d_RNIMCVI41Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4BCT_10_LC_10_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNI4BCT_10_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4BCT_10_LC_10_15_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNI4BCT_10_LC_10_15_1  (
            .in0(N__43304),
            .in1(_gnd_net_),
            .in2(N__36034),
            .in3(N__58234),
            .lcout(\ALU.d_RNI4BCTZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0SI26_6_LC_10_15_2 .C_ON=1'b0;
    defparam \ALU.d_RNI0SI26_6_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0SI26_6_LC_10_15_2 .LUT_INIT=16'b1011000010111111;
    LogicCell40 \ALU.d_RNI0SI26_6_LC_10_15_2  (
            .in0(N__49798),
            .in1(N__27572),
            .in2(N__71448),
            .in3(N__27818),
            .lcout(\ALU.combOperand2_0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI4VJC1_12_LC_10_15_3 .C_ON=1'b0;
    defparam \ALU.b_RNI4VJC1_12_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI4VJC1_12_LC_10_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_RNI4VJC1_12_LC_10_15_3  (
            .in0(N__43306),
            .in1(N__57685),
            .in2(_gnd_net_),
            .in3(N__39818),
            .lcout(\ALU.b_RNI4VJC1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI0RJC1_10_LC_10_15_4 .C_ON=1'b0;
    defparam \ALU.b_RNI0RJC1_10_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI0RJC1_10_LC_10_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.b_RNI0RJC1_10_LC_10_15_4  (
            .in0(N__36003),
            .in1(N__39137),
            .in2(_gnd_net_),
            .in3(N__43305),
            .lcout(),
            .ltout(\ALU.b_RNI0RJC1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHRVC5_10_LC_10_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNIHRVC5_10_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHRVC5_10_LC_10_15_5 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \ALU.d_RNIHRVC5_10_LC_10_15_5  (
            .in0(N__26915),
            .in1(N__27857),
            .in2(N__26909),
            .in3(N__53965),
            .lcout(\ALU.operand2_10 ),
            .ltout(\ALU.operand2_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINK8QF_10_LC_10_15_6 .C_ON=1'b0;
    defparam \ALU.d_RNINK8QF_10_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINK8QF_10_LC_10_15_6 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \ALU.d_RNINK8QF_10_LC_10_15_6  (
            .in0(N__71410),
            .in1(_gnd_net_),
            .in2(N__26981),
            .in3(N__37112),
            .lcout(\ALU.status_19_9 ),
            .ltout(\ALU.status_19_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0LDMJ_1_LC_10_15_7 .C_ON=1'b0;
    defparam \ALU.d_RNI0LDMJ_1_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0LDMJ_1_LC_10_15_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNI0LDMJ_1_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26978),
            .in3(N__65562),
            .lcout(\ALU.d_RNI0LDMJZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIBHMN_8_LC_10_16_0 .C_ON=1'b0;
    defparam \ALU.e_RNIBHMN_8_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIBHMN_8_LC_10_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.e_RNIBHMN_8_LC_10_16_0  (
            .in0(N__46280),
            .in1(N__48745),
            .in2(_gnd_net_),
            .in3(N__46944),
            .lcout(),
            .ltout(\ALU.e_RNIBHMNZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI34KF2_8_LC_10_16_1 .C_ON=1'b0;
    defparam \ALU.e_RNI34KF2_8_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI34KF2_8_LC_10_16_1 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.e_RNI34KF2_8_LC_10_16_1  (
            .in0(N__27968),
            .in1(N__53909),
            .in2(N__26975),
            .in3(N__46840),
            .lcout(\ALU.operand2_7_ns_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIINJ_8_LC_10_16_2 .C_ON=1'b0;
    defparam \ALU.d_RNIIINJ_8_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIINJ_8_LC_10_16_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIIINJ_8_LC_10_16_2  (
            .in0(N__48141),
            .in1(N__51580),
            .in2(_gnd_net_),
            .in3(N__43277),
            .lcout(\ALU.d_RNIIINJZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIE6BV_8_LC_10_16_4 .C_ON=1'b0;
    defparam \ALU.b_RNIE6BV_8_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIE6BV_8_LC_10_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.b_RNIE6BV_8_LC_10_16_4  (
            .in0(N__49045),
            .in1(N__48326),
            .in2(_gnd_net_),
            .in3(N__43279),
            .lcout(),
            .ltout(\ALU.b_RNIE6BVZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI77KG4_8_LC_10_16_5 .C_ON=1'b0;
    defparam \ALU.d_RNI77KG4_8_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI77KG4_8_LC_10_16_5 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \ALU.d_RNI77KG4_8_LC_10_16_5  (
            .in0(N__26972),
            .in1(N__26966),
            .in2(N__26960),
            .in3(N__53910),
            .lcout(\ALU.operand2_8 ),
            .ltout(\ALU.operand2_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI844QD_8_LC_10_16_6 .C_ON=1'b0;
    defparam \ALU.d_RNI844QD_8_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI844QD_8_LC_10_16_6 .LUT_INIT=16'b0111010011111100;
    LogicCell40 \ALU.d_RNI844QD_8_LC_10_16_6  (
            .in0(N__26948),
            .in1(N__71423),
            .in2(N__26942),
            .in3(N__27835),
            .lcout(\ALU.status_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI230L_10_LC_10_16_7 .C_ON=1'b0;
    defparam \ALU.c_RNI230L_10_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI230L_10_LC_10_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNI230L_10_LC_10_16_7  (
            .in0(N__43278),
            .in1(N__35722),
            .in2(_gnd_net_),
            .in3(N__36136),
            .lcout(\ALU.c_RNI230LZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_3_c_RNO_LC_10_17_0 .C_ON=1'b0;
    defparam \ALU.status_18_cry_3_c_RNO_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_3_c_RNO_LC_10_17_0 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \ALU.status_18_cry_3_c_RNO_LC_10_17_0  (
            .in0(N__38058),
            .in1(N__60218),
            .in2(N__33057),
            .in3(N__53238),
            .lcout(\ALU.status_18_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIUV6T5_2_LC_10_17_1 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIUV6T5_2_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIUV6T5_2_LC_10_17_1 .LUT_INIT=16'b0101010101000101;
    LogicCell40 \CONTROL.busState_1_RNIUV6T5_2_LC_10_17_1  (
            .in0(N__28576),
            .in1(N__49524),
            .in2(N__60247),
            .in3(N__50203),
            .lcout(N_228_0),
            .ltout(N_228_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHMDUU_3_LC_10_17_2 .C_ON=1'b0;
    defparam \ALU.d_RNIHMDUU_3_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHMDUU_3_LC_10_17_2 .LUT_INIT=16'b0000000011010001;
    LogicCell40 \ALU.d_RNIHMDUU_3_LC_10_17_2  (
            .in0(N__38057),
            .in1(N__53237),
            .in2(N__27029),
            .in3(N__68939),
            .lcout(\ALU.lshift62_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_3_LC_10_17_3 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_3_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_3_LC_10_17_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_3_LC_10_17_3  (
            .in0(N__27020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C_net ),
            .ce(N__32299),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI9NJL_3_LC_10_17_4 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI9NJL_3_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI9NJL_3_LC_10_17_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI9NJL_3_LC_10_17_4  (
            .in0(N__27026),
            .in1(N__32295),
            .in2(_gnd_net_),
            .in3(N__27019),
            .lcout(),
            .ltout(DROM_ROMDATA_dintern_3ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIDU0U1_2_LC_10_17_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIDU0U1_2_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIDU0U1_2_LC_10_17_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \CONTROL.busState_1_RNIDU0U1_2_LC_10_17_5  (
            .in0(N__49561),
            .in1(N__50280),
            .in2(N__27008),
            .in3(N__50202),
            .lcout(busState_1_RNIDU0U1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_adflt_LC_10_17_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_adflt_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_adflt_LC_10_17_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DROM.ROMDATA.dintern_adflt_LC_10_17_6  (
            .in0(N__27936),
            .in1(N__27898),
            .in2(_gnd_net_),
            .in3(N__27119),
            .lcout(DROM_ROMDATA_dintern_adflt),
            .ltout(DROM_ROMDATA_dintern_adflt_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIBS0U1_2_LC_10_17_7 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIBS0U1_2_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIBS0U1_2_LC_10_17_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \CONTROL.busState_1_RNIBS0U1_2_LC_10_17_7  (
            .in0(N__27005),
            .in1(N__49523),
            .in2(N__26999),
            .in3(N__50201),
            .lcout(busState_1_RNIBS0U1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_adflt_3_LC_10_18_0 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_adflt_3_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_adflt_3_LC_10_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DROM.ROMDATA.dintern_adflt_3_LC_10_18_0  (
            .in0(N__27113),
            .in1(N__27088),
            .in2(N__27938),
            .in3(N__27101),
            .lcout(\DROM.ROMDATA.dintern_adfltZ0Z_3 ),
            .ltout(\DROM.ROMDATA.dintern_adfltZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI5NIF1_0_LC_10_18_1 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI5NIF1_0_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI5NIF1_0_LC_10_18_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI5NIF1_0_LC_10_18_1  (
            .in0(N__27897),
            .in1(N__28003),
            .in2(N__27122),
            .in3(N__27955),
            .lcout(romOut_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_RNIDE6K_12_LC_10_18_2 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_RNIDE6K_12_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_RNIDE6K_12_LC_10_18_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \CONTROL.romAddReg_RNIDE6K_12_LC_10_18_2  (
            .in0(N__27954),
            .in1(N__27896),
            .in2(N__27937),
            .in3(N__50127),
            .lcout(\CONTROL.bus_6_a0_sx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_adflt_sx_LC_10_18_3 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_adflt_sx_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_adflt_sx_LC_10_18_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DROM.ROMDATA.dintern_adflt_sx_LC_10_18_3  (
            .in0(N__27099),
            .in1(N__27111),
            .in2(N__27089),
            .in3(N__27953),
            .lcout(\DROM.ROMDATA.dintern_adflt_sxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_adflt_3_x_LC_10_18_4 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_adflt_3_x_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_adflt_3_x_LC_10_18_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DROM.ROMDATA.dintern_adflt_3_x_LC_10_18_4  (
            .in0(N__27112),
            .in1(N__27087),
            .in2(_gnd_net_),
            .in3(N__27100),
            .lcout(dintern_adflt_3_x),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_13_LC_10_18_5 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_13_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.romAddReg_13_LC_10_18_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.romAddReg_13_LC_10_18_5  (
            .in0(N__27989),
            .in1(N__72102),
            .in2(N__52357),
            .in3(N__71870),
            .lcout(dataRomAddress_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.romAddReg_13C_net ),
            .ce(N__28111),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_14_LC_10_18_6 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_14_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.romAddReg_14_LC_10_18_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \CONTROL.romAddReg_14_LC_10_18_6  (
            .in0(N__71869),
            .in1(N__52304),
            .in2(N__31412),
            .in3(N__72104),
            .lcout(dataRomAddress_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.romAddReg_13C_net ),
            .ce(N__28111),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_15_LC_10_18_7 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_15_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.romAddReg_15_LC_10_18_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.romAddReg_15_LC_10_18_7  (
            .in0(N__45009),
            .in1(N__72103),
            .in2(N__50405),
            .in3(N__71871),
            .lcout(dataRomAddress_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.romAddReg_13C_net ),
            .ce(N__28111),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_ne_0_LC_10_19_0 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_ne_0_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_ne_0_LC_10_19_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \CONTROL.aluOperation_ne_0_LC_10_19_0  (
            .in0(N__41432),
            .in1(N__71872),
            .in2(_gnd_net_),
            .in3(N__54689),
            .lcout(aluOperation_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluOperation_ne_0C_net ),
            .ce(N__38144),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIDJR11_1_LC_10_19_1 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIDJR11_1_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIDJR11_1_LC_10_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIDJR11_1_LC_10_19_1  (
            .in0(N__27074),
            .in1(N__27067),
            .in2(_gnd_net_),
            .in3(N__32264),
            .lcout(DROM_ROMDATA_dintern_13ro),
            .ltout(DROM_ROMDATA_dintern_13ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIN5MIA_0_0_LC_10_19_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIN5MIA_0_0_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIN5MIA_0_0_LC_10_19_2 .LUT_INIT=16'b0000110011001100;
    LogicCell40 \CONTROL.busState_1_RNIN5MIA_0_0_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__34456),
            .in2(N__27293),
            .in3(N__27286),
            .lcout(bus_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIN5MIA_0_LC_10_19_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIN5MIA_0_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIN5MIA_0_LC_10_19_3 .LUT_INIT=16'b1111010101010101;
    LogicCell40 \CONTROL.busState_1_RNIN5MIA_0_LC_10_19_3  (
            .in0(N__34457),
            .in1(_gnd_net_),
            .in2(N__27290),
            .in3(N__27248),
            .lcout(bus_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNICAEO_2_LC_10_19_4 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNICAEO_2_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNICAEO_2_LC_10_19_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_RNICAEO_2_LC_10_19_4  (
            .in0(N__32263),
            .in1(N__27410),
            .in2(_gnd_net_),
            .in3(N__27433),
            .lcout(DROM_ROMDATA_dintern_10ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI9V0V_1_LC_10_19_5 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI9V0V_1_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI9V0V_1_LC_10_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI9V0V_1_LC_10_19_5  (
            .in0(N__27155),
            .in1(N__27178),
            .in2(_gnd_net_),
            .in3(N__32260),
            .lcout(DROM_ROMDATA_dintern_5ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIA01V_2_LC_10_19_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIA01V_2_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIA01V_2_LC_10_19_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIA01V_2_LC_10_19_6  (
            .in0(N__32261),
            .in1(N__27128),
            .in2(_gnd_net_),
            .in3(N__27145),
            .lcout(DROM_ROMDATA_dintern_6ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIB9EO_1_LC_10_19_7 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIB9EO_1_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIB9EO_1_LC_10_19_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIB9EO_1_LC_10_19_7  (
            .in0(N__27443),
            .in1(N__27466),
            .in2(_gnd_net_),
            .in3(N__32262),
            .lcout(DROM_ROMDATA_dintern_9ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_0_LC_10_20_0 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_0_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_0_LC_10_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_0_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28033),
            .lcout(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_1_LC_10_20_1 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_1_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_1_LC_10_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_1_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27179),
            .lcout(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_2_LC_10_20_2 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_2_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_2_LC_10_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_2_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27149),
            .lcout(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_3_LC_10_20_3 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_3_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_3_LC_10_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_3_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28061),
            .lcout(\DROM.ROMDATA.dintern_0_1_OLDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_1_LC_10_20_4 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_1_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_1_LC_10_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_1_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27467),
            .lcout(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_2_LC_10_20_5 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_2_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_2_LC_10_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_2_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27434),
            .lcout(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_3_LC_10_20_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_3_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_2_OLD_ne_3_LC_10_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_2_OLD_ne_3_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27404),
            .lcout(\DROM.ROMDATA.dintern_0_2_OLDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_0_LC_10_20_7 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_0_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_3_OLD_ne_0_LC_10_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DROM.ROMDATA.dintern_0_3_OLD_ne_0_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27377),
            .lcout(\DROM.ROMDATA.dintern_0_3_OLDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net ),
            .ce(N__32320),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_6_LC_10_21_0 .C_ON=1'b0;
    defparam \CONTROL.dout_6_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_6_LC_10_21_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \CONTROL.dout_6_LC_10_21_0  (
            .in0(N__40892),
            .in1(N__43744),
            .in2(N__79531),
            .in3(N__71579),
            .lcout(\CONTROL.ctrlOut_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_6C_net ),
            .ce(N__44457),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI5P5Q5_1_LC_10_21_1 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI5P5Q5_1_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI5P5Q5_1_LC_10_21_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \CONTROL.busState_1_RNI5P5Q5_1_LC_10_21_1  (
            .in0(N__62556),
            .in1(N__50324),
            .in2(N__27346),
            .in3(N__50113),
            .lcout(),
            .ltout(\CONTROL.N_199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIF3TV7_0_LC_10_21_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIF3TV7_0_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIF3TV7_0_LC_10_21_2 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \CONTROL.busState_1_RNIF3TV7_0_LC_10_21_2  (
            .in0(N__49786),
            .in1(N__27571),
            .in2(N__27314),
            .in3(N__49553),
            .lcout(bus_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI8OOJ_6_LC_10_21_3 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI8OOJ_6_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI8OOJ_6_LC_10_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNI8OOJ_6_LC_10_21_3  (
            .in0(N__27311),
            .in1(N__45583),
            .in2(_gnd_net_),
            .in3(N__50111),
            .lcout(),
            .ltout(\CONTROL.N_167_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI4TRD1_2_LC_10_21_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI4TRD1_2_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI4TRD1_2_LC_10_21_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \CONTROL.busState_1_RNI4TRD1_2_LC_10_21_4  (
            .in0(N__50112),
            .in1(N__27596),
            .in2(N__27575),
            .in3(N__49552),
            .lcout(N_183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_22dflt_LC_10_21_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_22dflt_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_22dflt_LC_10_21_5 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_22dflt_LC_10_21_5  (
            .in0(N__71578),
            .in1(N__79514),
            .in2(N__43745),
            .in3(N__40889),
            .lcout(controlWord_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_4_LC_10_21_6 .C_ON=1'b0;
    defparam \CONTROL.dout_4_LC_10_21_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_4_LC_10_21_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \CONTROL.dout_4_LC_10_21_6  (
            .in0(N__40891),
            .in1(N__65236),
            .in2(N__79530),
            .in3(N__74213),
            .lcout(\CONTROL.ctrlOut_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_6C_net ),
            .ce(N__44457),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_20dflt_LC_10_21_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_20dflt_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_20dflt_LC_10_21_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_20dflt_LC_10_21_7  (
            .in0(N__74212),
            .in1(N__79515),
            .in2(N__65237),
            .in3(N__40890),
            .lcout(controlWord_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI37DAN91_3_LC_10_22_0 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI37DAN91_3_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI37DAN91_3_LC_10_22_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI37DAN91_3_LC_10_22_0  (
            .in0(N__34771),
            .in1(N__57821),
            .in2(N__27659),
            .in3(N__41982),
            .lcout(\CONTROL.addrstackptr_N_8_mux_1_0 ),
            .ltout(\CONTROL.addrstackptr_N_8_mux_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNIAEEIH92_5_LC_10_22_1 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNIAEEIH92_5_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNIAEEIH92_5_LC_10_22_1 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \CONTROL.addrstackptr_RNIAEEIH92_5_LC_10_22_1  (
            .in0(N__27493),
            .in1(N__27529),
            .in2(N__27557),
            .in3(N__27536),
            .lcout(\CONTROL.addrstackptr_N_6_0_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_0_7_LC_10_22_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_0_7_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_0_7_LC_10_22_2 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIO2O5VB_0_7_LC_10_22_2  (
            .in0(N__54681),
            .in1(N__41488),
            .in2(N__71876),
            .in3(N__44696),
            .lcout(),
            .ltout(\CONTROL.g0_3_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIFRI6PV_0_7_LC_10_22_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIFRI6PV_0_7_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIFRI6PV_0_7_LC_10_22_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIFRI6PV_0_7_LC_10_22_3  (
            .in0(N__27665),
            .in1(N__38185),
            .in2(N__27539),
            .in3(N__27671),
            .lcout(\CONTROL.N_4_0 ),
            .ltout(\CONTROL.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_5_LC_10_22_4 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_5_LC_10_22_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_5_LC_10_22_4 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \CONTROL.addrstackptr_5_LC_10_22_4  (
            .in0(N__27530),
            .in1(N__27494),
            .in2(N__27509),
            .in3(N__27506),
            .lcout(\CONTROL.addrstackptrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.addrstackptr_5C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_1_LC_10_22_5 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_1_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_1_LC_10_22_5 .LUT_INIT=16'b1011111101111111;
    LogicCell40 \CONTROL.g0_3_i_1_LC_10_22_5  (
            .in0(N__42265),
            .in1(N__55470),
            .in2(N__72284),
            .in3(N__54680),
            .lcout(\CONTROL.g0_3_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_a7_2_LC_10_22_6 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_a7_2_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_a7_2_LC_10_22_6 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \CONTROL.g0_3_i_a7_2_LC_10_22_6  (
            .in0(N__54679),
            .in1(N__40676),
            .in2(N__63485),
            .in3(N__38272),
            .lcout(\CONTROL.g0_3_i_a7Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI1E361_4_LC_10_23_0 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI1E361_4_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI1E361_4_LC_10_23_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI1E361_4_LC_10_23_0  (
            .in0(N__38441),
            .in1(_gnd_net_),
            .in2(N__60814),
            .in3(N__60723),
            .lcout(\CONTROL.g0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_12_LC_10_23_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_12_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_12_LC_10_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_12_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27647),
            .lcout(\CONTROL.addrstack_reto_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73269),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_11_LC_10_23_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_11_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_11_LC_10_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_11_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27632),
            .lcout(CONTROL_addrstack_reto_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73269),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_13_LC_10_23_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_13_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_13_LC_10_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_13_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43676),
            .lcout(\CONTROL.dout_reto_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73269),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_7_LC_10_23_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_7_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_7_LC_10_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_7_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27620),
            .lcout(\CONTROL.addrstack_reto_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73269),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_14_LC_10_23_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_14_LC_10_23_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_14_LC_10_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_14_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27608),
            .lcout(\CONTROL.addrstack_reto_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73269),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIJDJ31_3_LC_10_23_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIJDJ31_3_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIJDJ31_3_LC_10_23_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIJDJ31_3_LC_10_23_6  (
            .in0(N__73668),
            .in1(N__64532),
            .in2(_gnd_net_),
            .in3(N__64487),
            .lcout(\CONTROL.programCounter_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_11_LC_10_24_1 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_11_LC_10_24_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_11_LC_10_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_11_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29726),
            .lcout(\CONTROL.tempCounterZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_11C_net ),
            .ce(N__34966),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_15_LC_10_24_5 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_15_LC_10_24_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_15_LC_10_24_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.tempCounter_15_LC_10_24_5  (
            .in0(N__33457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.tempCounterZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_11C_net ),
            .ce(N__34966),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_14_LC_10_24_7 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_14_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_14_LC_10_24_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.tempCounter_14_LC_10_24_7  (
            .in0(N__29648),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.tempCounterZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_11C_net ),
            .ce(N__34966),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_8_LC_10_25_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_8_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_8_LC_10_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_8_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27701),
            .lcout(CONTROL_addrstack_reto_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73278),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_9_LC_10_25_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_9_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_9_LC_10_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_9_LC_10_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27692),
            .lcout(\CONTROL.addrstack_reto_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73278),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHJSI82_4_LC_11_8_6 .C_ON=1'b0;
    defparam \ALU.d_RNIHJSI82_4_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHJSI82_4_LC_11_8_6 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.d_RNIHJSI82_4_LC_11_8_6  (
            .in0(N__59842),
            .in1(N__59585),
            .in2(N__28472),
            .in3(N__65953),
            .lcout(\ALU.N_860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFGGBO_0_6_LC_11_9_1 .C_ON=1'b0;
    defparam \ALU.d_RNIFGGBO_0_6_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFGGBO_0_6_LC_11_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIFGGBO_0_6_LC_11_9_1  (
            .in0(N__62570),
            .in1(N__62307),
            .in2(_gnd_net_),
            .in3(N__66735),
            .lcout(\ALU.N_609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_9_c_RNO_LC_11_9_2 .C_ON=1'b0;
    defparam \ALU.status_17_I_9_c_RNO_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_9_c_RNO_LC_11_9_2 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ALU.status_17_I_9_c_RNO_LC_11_9_2  (
            .in0(N__68270),
            .in1(N__66298),
            .in2(N__60262),
            .in3(N__68825),
            .lcout(\ALU.status_17_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI0QV651_10_LC_11_9_3 .C_ON=1'b0;
    defparam \ALU.c_RNI0QV651_10_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI0QV651_10_LC_11_9_3 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.c_RNI0QV651_10_LC_11_9_3  (
            .in0(N__56240),
            .in1(N__61426),
            .in2(N__61668),
            .in3(N__56394),
            .lcout(\ALU.c_RNI0QV651Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIOFVDI_5_LC_11_9_4 .C_ON=1'b0;
    defparam \ALU.d_RNIOFVDI_5_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIOFVDI_5_LC_11_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIOFVDI_5_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__59483),
            .in2(_gnd_net_),
            .in3(N__56239),
            .lcout(\ALU.d_RNIOFVDIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPNF141_4_LC_11_9_6 .C_ON=1'b0;
    defparam \ALU.d_RNIPNF141_4_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPNF141_4_LC_11_9_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNIPNF141_4_LC_11_9_6  (
            .in0(N__59840),
            .in1(N__55681),
            .in2(N__55816),
            .in3(N__59485),
            .lcout(\ALU.d_RNIPNF141Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI88K161_4_LC_11_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNI88K161_4_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI88K161_4_LC_11_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI88K161_4_LC_11_9_7  (
            .in0(N__59484),
            .in1(N__59841),
            .in2(N__55688),
            .in3(N__55585),
            .lcout(\ALU.d_RNI88K161Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_2_LC_11_10_0 .C_ON=1'b0;
    defparam \ALU.h_2_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_2_LC_11_10_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.h_2_LC_11_10_0  (
            .in0(N__39479),
            .in1(N__39611),
            .in2(_gnd_net_),
            .in3(N__39539),
            .lcout(h_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73148),
            .ce(N__69458),
            .sr(_gnd_net_));
    defparam \ALU.h_4_LC_11_10_1 .C_ON=1'b0;
    defparam \ALU.h_4_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \ALU.h_4_LC_11_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.h_4_LC_11_10_1  (
            .in0(N__57421),
            .in1(N__42549),
            .in2(_gnd_net_),
            .in3(N__39377),
            .lcout(h_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73148),
            .ce(N__69458),
            .sr(_gnd_net_));
    defparam \ALU.h_5_LC_11_10_2 .C_ON=1'b0;
    defparam \ALU.h_5_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.h_5_LC_11_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.h_5_LC_11_10_2  (
            .in0(N__57422),
            .in1(N__39319),
            .in2(_gnd_net_),
            .in3(N__52635),
            .lcout(h_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73148),
            .ce(N__69458),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITPMMO_0_6_LC_11_10_3 .C_ON=1'b0;
    defparam \ALU.d_RNITPMMO_0_6_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITPMMO_0_6_LC_11_10_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNITPMMO_0_6_LC_11_10_3  (
            .in0(N__62551),
            .in1(N__59479),
            .in2(_gnd_net_),
            .in3(N__66733),
            .lcout(\ALU.N_608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITPMMO_6_LC_11_10_4 .C_ON=1'b0;
    defparam \ALU.d_RNITPMMO_6_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITPMMO_6_LC_11_10_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNITPMMO_6_LC_11_10_4  (
            .in0(N__66734),
            .in1(_gnd_net_),
            .in2(N__59540),
            .in3(N__62552),
            .lcout(\ALU.N_833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2RK5I_5_LC_11_10_5 .C_ON=1'b0;
    defparam \ALU.d_RNI2RK5I_5_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2RK5I_5_LC_11_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI2RK5I_5_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__59476),
            .in2(_gnd_net_),
            .in3(N__56360),
            .lcout(\ALU.d_RNI2RK5IZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6HBMG_5_LC_11_10_6 .C_ON=1'b0;
    defparam \ALU.d_RNI6HBMG_5_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6HBMG_5_LC_11_10_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI6HBMG_5_LC_11_10_6  (
            .in0(N__59477),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55985),
            .lcout(\ALU.d_RNI6HBMGZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIB5POH_5_LC_11_10_7 .C_ON=1'b0;
    defparam \ALU.d_RNIB5POH_5_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIB5POH_5_LC_11_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIB5POH_5_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__59478),
            .in2(_gnd_net_),
            .in3(N__55768),
            .lcout(\ALU.d_RNIB5POHZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMQM8I_5_LC_11_11_0 .C_ON=1'b0;
    defparam \ALU.d_RNIMQM8I_5_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMQM8I_5_LC_11_11_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIMQM8I_5_LC_11_11_0  (
            .in0(N__55661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59549),
            .lcout(\ALU.d_RNIMQM8IZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISSV4I_9_LC_11_11_1 .C_ON=1'b0;
    defparam \ALU.d_RNISSV4I_9_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISSV4I_9_LC_11_11_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNISSV4I_9_LC_11_11_1  (
            .in0(N__56202),
            .in1(N__62829),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ALU.d_RNISSV4IZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIK9E841_6_LC_11_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNIK9E841_6_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIK9E841_6_LC_11_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIK9E841_6_LC_11_11_2  (
            .in0(N__56359),
            .in1(N__62518),
            .in2(N__62315),
            .in3(N__56201),
            .lcout(\ALU.d_RNIK9E841Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJ0U031_2_LC_11_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIJ0U031_2_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJ0U031_2_LC_11_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIJ0U031_2_LC_11_11_3  (
            .in0(N__56068),
            .in1(N__60190),
            .in2(N__56229),
            .in3(N__66297),
            .lcout(\ALU.d_RNIJ0U031Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIV1LMH_3_LC_11_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNIV1LMH_3_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIV1LMH_3_LC_11_11_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIV1LMH_3_LC_11_11_4  (
            .in0(N__60189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56200),
            .lcout(\ALU.d_RNIV1LMHZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9DAEH_3_LC_11_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNI9DAEH_3_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9DAEH_3_LC_11_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI9DAEH_3_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__60188),
            .in2(_gnd_net_),
            .in3(N__56357),
            .lcout(\ALU.d_RNI9DAEHZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIITFA41_0_LC_11_11_7 .C_ON=1'b0;
    defparam \ALU.d_RNIITFA41_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIITFA41_0_LC_11_11_7 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.d_RNIITFA41_0_LC_11_11_7  (
            .in0(N__65539),
            .in1(N__60589),
            .in2(N__56228),
            .in3(N__56358),
            .lcout(\ALU.d_RNIITFA41Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISP66I_1_LC_11_12_0 .C_ON=1'b0;
    defparam \ALU.d_RNISP66I_1_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISP66I_1_LC_11_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNISP66I_1_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__55660),
            .in2(_gnd_net_),
            .in3(N__65541),
            .lcout(\ALU.d_RNISP66IZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKRBVN_4_LC_11_12_1 .C_ON=1'b0;
    defparam \ALU.d_RNIKRBVN_4_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKRBVN_4_LC_11_12_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.d_RNIKRBVN_4_LC_11_12_1  (
            .in0(N__60192),
            .in1(_gnd_net_),
            .in2(N__59866),
            .in3(N__66662),
            .lcout(\ALU.N_831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKG0L11_2_LC_11_12_2 .C_ON=1'b0;
    defparam \ALU.d_RNIKG0L11_2_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKG0L11_2_LC_11_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIKG0L11_2_LC_11_12_2  (
            .in0(N__56327),
            .in1(N__60196),
            .in2(N__68505),
            .in3(N__66269),
            .lcout(\ALU.d_RNIKG0L11Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI12A911_2_LC_11_12_3 .C_ON=1'b0;
    defparam \ALU.d_RNI12A911_2_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI12A911_2_LC_11_12_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNI12A911_2_LC_11_12_3  (
            .in0(N__66270),
            .in1(N__55959),
            .in2(N__60241),
            .in3(N__56082),
            .lcout(\ALU.d_RNI12A911Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINIF011_2_LC_11_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNINIF011_2_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINIF011_2_LC_11_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNINIF011_2_LC_11_12_4  (
            .in0(N__60227),
            .in1(N__55767),
            .in2(N__55984),
            .in3(N__66271),
            .lcout(\ALU.d_RNINIF011Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJTUN21_4_LC_11_12_5 .C_ON=1'b0;
    defparam \ALU.d_RNIJTUN21_4_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJTUN21_4_LC_11_12_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNIJTUN21_4_LC_11_12_5  (
            .in0(N__59817),
            .in1(N__55960),
            .in2(N__56096),
            .in3(N__59550),
            .lcout(\ALU.d_RNIJTUN21Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIS69AH_3_LC_11_12_6 .C_ON=1'b0;
    defparam \ALU.d_RNIS69AH_3_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIS69AH_3_LC_11_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIS69AH_3_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__60191),
            .in2(_gnd_net_),
            .in3(N__56069),
            .lcout(\ALU.d_RNIS69AHZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8Q43I_1_LC_11_12_7 .C_ON=1'b0;
    defparam \ALU.d_RNI8Q43I_1_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8Q43I_1_LC_11_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI8Q43I_1_LC_11_12_7  (
            .in0(N__65540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56326),
            .lcout(\ALU.d_RNI8Q43IZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_3_c_RNIGCKVJ5_LC_11_13_0 .C_ON=1'b0;
    defparam \ALU.addsub_cry_3_c_RNIGCKVJ5_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_3_c_RNIGCKVJ5_LC_11_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.addsub_cry_3_c_RNIGCKVJ5_LC_11_13_0  (
            .in0(N__59672),
            .in1(N__66976),
            .in2(_gnd_net_),
            .in3(N__35282),
            .lcout(),
            .ltout(\ALU.addsub_cry_3_c_RNIGCKVJZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_3_c_RNIM4CUT9_LC_11_13_1 .C_ON=1'b0;
    defparam \ALU.addsub_cry_3_c_RNIM4CUT9_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_3_c_RNIM4CUT9_LC_11_13_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \ALU.addsub_cry_3_c_RNIM4CUT9_LC_11_13_1  (
            .in0(N__34178),
            .in1(N__48554),
            .in2(N__27746),
            .in3(N__68431),
            .lcout(\ALU.addsub_cry_3_c_RNIM4CUTZ0Z9 ),
            .ltout(\ALU.addsub_cry_3_c_RNIM4CUTZ0Z9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_4_LC_11_13_2 .C_ON=1'b0;
    defparam \ALU.a_4_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.a_4_LC_11_13_2 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \ALU.a_4_LC_11_13_2  (
            .in0(N__42550),
            .in1(N__57406),
            .in2(N__27743),
            .in3(_gnd_net_),
            .lcout(\ALU.aZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73168),
            .ce(N__71212),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI26JM_4_LC_11_13_3 .C_ON=1'b0;
    defparam \ALU.e_RNI26JM_4_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI26JM_4_LC_11_13_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.e_RNI26JM_4_LC_11_13_3  (
            .in0(N__44000),
            .in1(_gnd_net_),
            .in2(N__32663),
            .in3(N__27782),
            .lcout(),
            .ltout(\ALU.e_RNI26JMZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIFKVD2_4_LC_11_13_4 .C_ON=1'b0;
    defparam \ALU.e_RNIFKVD2_4_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIFKVD2_4_LC_11_13_4 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.e_RNIFKVD2_4_LC_11_13_4  (
            .in0(N__53956),
            .in1(N__53435),
            .in2(N__27740),
            .in3(N__27791),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI19244_4_LC_11_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNI19244_4_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI19244_4_LC_11_13_5 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNI19244_4_LC_11_13_5  (
            .in0(N__43325),
            .in1(N__53957),
            .in2(N__27800),
            .in3(N__43430),
            .lcout(\ALU.operand2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI6IVQ_4_LC_11_13_6 .C_ON=1'b0;
    defparam \ALU.c_RNI6IVQ_4_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI6IVQ_4_LC_11_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNI6IVQ_4_LC_11_13_6  (
            .in0(N__35796),
            .in1(N__35852),
            .in2(_gnd_net_),
            .in3(N__43999),
            .lcout(\ALU.c_RNI6IVQZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI6DH51_4_LC_11_14_0 .C_ON=1'b0;
    defparam \ALU.b_RNI6DH51_4_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI6DH51_4_LC_11_14_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI6DH51_4_LC_11_14_0  (
            .in0(N__43448),
            .in1(N__34560),
            .in2(N__44155),
            .in3(N__43920),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEGPK1_4_LC_11_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNIEGPK1_4_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEGPK1_4_LC_11_14_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.d_RNIEGPK1_4_LC_11_14_1  (
            .in0(N__43348),
            .in1(N__43386),
            .in2(N__27785),
            .in3(N__47203),
            .lcout(\ALU.N_1137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI47B31_4_LC_11_14_2 .C_ON=1'b0;
    defparam \ALU.e_RNI47B31_4_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI47B31_4_LC_11_14_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNI47B31_4_LC_11_14_2  (
            .in0(N__27781),
            .in1(N__34561),
            .in2(N__32662),
            .in3(N__43921),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIA4D02_4_LC_11_14_3 .C_ON=1'b0;
    defparam \ALU.c_RNIA4D02_4_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIA4D02_4_LC_11_14_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNIA4D02_4_LC_11_14_3  (
            .in0(N__35797),
            .in1(N__35851),
            .in2(N__27770),
            .in3(N__47204),
            .lcout(),
            .ltout(\ALU.N_1089_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIROKU3_4_LC_11_14_4 .C_ON=1'b0;
    defparam \ALU.d_RNIROKU3_4_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIROKU3_4_LC_11_14_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIROKU3_4_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__54138),
            .in2(N__27767),
            .in3(N__27764),
            .lcout(aluOut_4),
            .ltout(aluOut_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBJM75_4_LC_11_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNIBJM75_4_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBJM75_4_LC_11_14_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.d_RNIBJM75_4_LC_11_14_5  (
            .in0(N__53245),
            .in1(N__49583),
            .in2(N__27758),
            .in3(N__50199),
            .lcout(\ALU.d_RNIBJM75Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI990621_0_LC_11_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNI990621_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI990621_0_LC_11_15_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNI990621_0_LC_11_15_0  (
            .in0(N__55994),
            .in1(N__65538),
            .in2(N__60609),
            .in3(N__55724),
            .lcout(\ALU.d_RNI990621Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRU9M31_6_LC_11_15_2 .C_ON=1'b0;
    defparam \ALU.d_RNIRU9M31_6_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRU9M31_6_LC_11_15_2 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.d_RNIRU9M31_6_LC_11_15_2  (
            .in0(N__62265),
            .in1(N__55647),
            .in2(N__62572),
            .in3(N__55726),
            .lcout(\ALU.d_RNIRU9M31Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIINE1H_3_LC_11_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNIINE1H_3_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIINE1H_3_LC_11_15_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIINE1H_3_LC_11_15_4  (
            .in0(N__60157),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55725),
            .lcout(\ALU.d_RNIINE1HZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKDVI51_4_LC_11_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNIKDVI51_4_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKDVI51_4_LC_11_15_5 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.d_RNIKDVI51_4_LC_11_15_5  (
            .in0(N__59800),
            .in1(N__59595),
            .in2(N__57024),
            .in3(N__55558),
            .lcout(\ALU.d_RNIKDVI51Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJP1AE_9_LC_11_15_6 .C_ON=1'b0;
    defparam \ALU.d_RNIJP1AE_9_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJP1AE_9_LC_11_15_6 .LUT_INIT=16'b1110110011111111;
    LogicCell40 \ALU.d_RNIJP1AE_9_LC_11_15_6  (
            .in0(N__40593),
            .in1(N__40540),
            .in2(N__40494),
            .in3(N__40520),
            .lcout(\ALU.status_19_8 ),
            .ltout(\ALU.status_19_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITCCHH_3_LC_11_15_7 .C_ON=1'b0;
    defparam \ALU.d_RNITCCHH_3_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITCCHH_3_LC_11_15_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNITCCHH_3_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27824),
            .in3(N__60158),
            .lcout(\ALU.d_RNITCCHHZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIPLDD2_6_LC_11_16_0 .C_ON=1'b0;
    defparam \ALU.e_RNIPLDD2_6_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIPLDD2_6_LC_11_16_0 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \ALU.e_RNIPLDD2_6_LC_11_16_0  (
            .in0(N__27806),
            .in1(N__27878),
            .in2(N__53969),
            .in3(N__46831),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJIG34_6_LC_11_16_1 .C_ON=1'b0;
    defparam \ALU.d_RNIJIG34_6_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJIG34_6_LC_11_16_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIJIG34_6_LC_11_16_1  (
            .in0(N__27872),
            .in1(N__27812),
            .in2(N__27821),
            .in3(N__53961),
            .lcout(\ALU.operand2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI9JSP_6_LC_11_16_2 .C_ON=1'b0;
    defparam \ALU.b_RNI9JSP_6_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI9JSP_6_LC_11_16_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.b_RNI9JSP_6_LC_11_16_2  (
            .in0(N__39899),
            .in1(N__70585),
            .in2(_gnd_net_),
            .in3(N__46943),
            .lcout(\ALU.b_RNI9JSPZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI6AJM_6_LC_11_16_3 .C_ON=1'b0;
    defparam \ALU.e_RNI6AJM_6_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI6AJM_6_LC_11_16_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_RNI6AJM_6_LC_11_16_3  (
            .in0(N__43998),
            .in1(N__32732),
            .in2(_gnd_net_),
            .in3(N__42937),
            .lcout(\ALU.e_RNI6AJMZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIAMVQ_6_LC_11_16_4 .C_ON=1'b0;
    defparam \ALU.c_RNIAMVQ_6_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIAMVQ_6_LC_11_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIAMVQ_6_LC_11_16_4  (
            .in0(N__35768),
            .in1(N__35834),
            .in2(_gnd_net_),
            .in3(N__43997),
            .lcout(\ALU.c_RNIAMVQZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDV8E_6_LC_11_16_5 .C_ON=1'b0;
    defparam \ALU.d_RNIDV8E_6_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDV8E_6_LC_11_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIDV8E_6_LC_11_16_5  (
            .in0(N__46942),
            .in1(N__37438),
            .in2(_gnd_net_),
            .in3(N__36062),
            .lcout(\ALU.d_RNIDV8EZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIUI741_10_LC_11_16_6 .C_ON=1'b0;
    defparam \ALU.a_RNIUI741_10_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIUI741_10_LC_11_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.a_RNIUI741_10_LC_11_16_6  (
            .in0(N__32635),
            .in1(N__37076),
            .in2(_gnd_net_),
            .in3(N__43287),
            .lcout(),
            .ltout(\ALU.a_RNIUI741Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI9B2L2_10_LC_11_16_7 .C_ON=1'b0;
    defparam \ALU.c_RNI9B2L2_10_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI9B2L2_10_LC_11_16_7 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.c_RNI9B2L2_10_LC_11_16_7  (
            .in0(N__46832),
            .in1(N__27866),
            .in2(N__27860),
            .in3(N__53962),
            .lcout(\ALU.operand2_7_ns_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNISTG51_8_LC_11_17_0 .C_ON=1'b0;
    defparam \ALU.b_RNISTG51_8_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNISTG51_8_LC_11_17_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNISTG51_8_LC_11_17_0  (
            .in0(N__48325),
            .in1(N__32825),
            .in2(N__49044),
            .in3(N__36341),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBFGH1_8_LC_11_17_1 .C_ON=1'b0;
    defparam \ALU.d_RNIBFGH1_8_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBFGH1_8_LC_11_17_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIBFGH1_8_LC_11_17_1  (
            .in0(N__48142),
            .in1(N__51587),
            .in2(N__27851),
            .in3(N__54297),
            .lcout(ALU_N_1141),
            .ltout(ALU_N_1141_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_RNIEQRR4_0_LC_11_17_2 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_RNIEQRR4_0_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_ne_RNIEQRR4_0_LC_11_17_2 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \CONTROL.operand1_ne_RNIEQRR4_0_LC_11_17_2  (
            .in0(N__34481),
            .in1(N__54141),
            .in2(N__27848),
            .in3(N__29026),
            .lcout(),
            .ltout(\CONTROL.bus_0_sx_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIA1EN6_0_0_LC_11_17_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIA1EN6_0_0_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIA1EN6_0_0_LC_11_17_3 .LUT_INIT=16'b0000110000001111;
    LogicCell40 \CONTROL.busState_1_RNIA1EN6_0_0_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__49758),
            .in2(N__27845),
            .in3(N__33166),
            .lcout(CONTROL_bus_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIQNA31_8_LC_11_17_4 .C_ON=1'b0;
    defparam \ALU.e_RNIQNA31_8_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIQNA31_8_LC_11_17_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNIQNA31_8_LC_11_17_4  (
            .in0(N__48752),
            .in1(N__32824),
            .in2(N__46279),
            .in3(N__36340),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI734T1_8_LC_11_17_5 .C_ON=1'b0;
    defparam \ALU.c_RNI734T1_8_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI734T1_8_LC_11_17_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNI734T1_8_LC_11_17_5  (
            .in0(N__50431),
            .in1(N__46378),
            .in2(N__27971),
            .in3(N__54296),
            .lcout(ALU_N_1093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFT2S_8_LC_11_17_6 .C_ON=1'b0;
    defparam \ALU.c_RNIFT2S_8_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFT2S_8_LC_11_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.c_RNIFT2S_8_LC_11_17_6  (
            .in0(N__46379),
            .in1(N__50430),
            .in2(_gnd_net_),
            .in3(N__46946),
            .lcout(\ALU.c_RNIFT2SZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_10_LC_11_18_0 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_10_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.romAddReg_10_LC_11_18_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.romAddReg_10_LC_11_18_0  (
            .in0(N__31277),
            .in1(N__72008),
            .in2(N__35723),
            .in3(N__71867),
            .lcout(dataRomAddress_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.romAddReg_10C_net ),
            .ce(N__28110),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_12_LC_11_18_1 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_12_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.romAddReg_12_LC_11_18_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \CONTROL.romAddReg_12_LC_11_18_1  (
            .in0(N__71866),
            .in1(N__28228),
            .in2(N__72140),
            .in3(N__52412),
            .lcout(dataRomAddress_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.romAddReg_10C_net ),
            .ce(N__28110),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_adflt_4_LC_11_18_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_adflt_4_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_adflt_4_LC_11_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PROM.ROMDATA.dintern_adflt_4_LC_11_18_2  (
            .in0(N__28310),
            .in1(N__28286),
            .in2(N__29747),
            .in3(N__28418),
            .lcout(\PROM.ROMDATA.dintern_adfltZ0Z_4 ),
            .ltout(\PROM.ROMDATA.dintern_adfltZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_adflt_LC_11_18_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_adflt_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_adflt_LC_11_18_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_adflt_LC_11_18_3  (
            .in0(N__28442),
            .in1(N__30346),
            .in2(N__27917),
            .in3(N__28519),
            .lcout(PROM_ROMDATA_dintern_adflt),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_12dflt_0_1_LC_11_18_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_12dflt_0_1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_12dflt_0_1_LC_11_18_4 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \PROM.ROMDATA.dintern_12dflt_0_1_LC_11_18_4  (
            .in0(N__30373),
            .in1(N__64663),
            .in2(N__30407),
            .in3(N__28441),
            .lcout(),
            .ltout(\PROM.ROMDATA.dintern_12dflt_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_12dflt_0_LC_11_18_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_12dflt_0_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_12dflt_0_LC_11_18_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_12dflt_0_LC_11_18_5  (
            .in0(N__72712),
            .in1(N__28520),
            .in2(N__27914),
            .in3(N__27911),
            .lcout(\PROM.ROMDATA.dintern_12dfltZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_11_LC_11_18_6 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_11_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.romAddReg_11_LC_11_18_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.romAddReg_11_LC_11_18_6  (
            .in0(N__35678),
            .in1(N__72009),
            .in2(N__31233),
            .in3(N__71868),
            .lcout(dataRomAddress_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.romAddReg_10C_net ),
            .ce(N__28110),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNO_0_0_LC_11_19_0 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNO_0_0_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNO_0_0_LC_11_19_0 .LUT_INIT=16'b0000000101010001;
    LogicCell40 \CONTROL.busState_1_RNO_0_0_LC_11_19_0  (
            .in0(N__35141),
            .in1(N__35189),
            .in2(N__41702),
            .in3(N__30794),
            .lcout(),
            .ltout(\CONTROL.busState_1_e_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_0_LC_11_19_1 .C_ON=1'b0;
    defparam \CONTROL.busState_1_0_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.busState_1_0_LC_11_19_1 .LUT_INIT=16'b1110111100100011;
    LogicCell40 \CONTROL.busState_1_0_LC_11_19_1  (
            .in0(N__28079),
            .in1(N__40636),
            .in2(N__28130),
            .in3(N__49742),
            .lcout(busState_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.busState_1_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState_1_sqmuxa_i_0_LC_11_19_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_0_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_0_LC_11_19_2 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \CONTROL.un1_busState_1_sqmuxa_i_0_LC_11_19_2  (
            .in0(N__38713),
            .in1(N__31466),
            .in2(N__29539),
            .in3(N__30793),
            .lcout(\CONTROL.un1_busState_1_sqmuxa_iZ0Z_0 ),
            .ltout(\CONTROL.un1_busState_1_sqmuxa_iZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState_1_sqmuxa_i_i_LC_11_19_3 .C_ON=1'b0;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_i_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_i_LC_11_19_3 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \CONTROL.un1_busState_1_sqmuxa_i_i_LC_11_19_3  (
            .in0(N__36621),
            .in1(N__38715),
            .in2(N__28127),
            .in3(N__54750),
            .lcout(N_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_1_LC_11_19_4 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_1_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_1_LC_11_19_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \CONTROL.busState_cnst_2_0__m11_0_a2_1_LC_11_19_4  (
            .in0(N__38714),
            .in1(N__41260),
            .in2(N__29540),
            .in3(N__41431),
            .lcout(\CONTROL.N_352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_sr_en_LC_11_19_5 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_sr_en_LC_11_19_5 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_0_sr_en_LC_11_19_5 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_sr_en_LC_11_19_5  (
            .in0(N__38716),
            .in1(N__54751),
            .in2(N__36626),
            .in3(N__28073),
            .lcout(\DROM.ROMDATA.dintern_0_0_sr_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.busState_1_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIB11V_3_LC_11_19_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIB11V_3_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIB11V_3_LC_11_19_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIB11V_3_LC_11_19_6  (
            .in0(N__28067),
            .in1(N__28057),
            .in2(_gnd_net_),
            .in3(N__32246),
            .lcout(DROM_ROMDATA_dintern_7ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI8U0V_0_LC_11_19_7 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI8U0V_0_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI8U0V_0_LC_11_19_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI8U0V_0_LC_11_19_7  (
            .in0(N__32247),
            .in1(N__28040),
            .in2(_gnd_net_),
            .in3(N__28034),
            .lcout(DROM_ROMDATA_dintern_4ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_29dflt_LC_11_20_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_29dflt_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_29dflt_LC_11_20_0 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \PROM.ROMDATA.dintern_29dflt_LC_11_20_0  (
            .in0(N__76637),
            .in1(N__43690),
            .in2(N__44324),
            .in3(N__43721),
            .lcout(controlWord_29),
            .ltout(controlWord_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_13_LC_11_20_1 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_13_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_13_LC_11_20_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \CONTROL.ramAddReg_13_LC_11_20_1  (
            .in0(N__70462),
            .in1(N__57621),
            .in2(N__28232),
            .in3(N__70763),
            .lcout(A13_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_13C_net ),
            .ce(N__70340),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_28dflt_LC_11_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_28dflt_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_28dflt_LC_11_20_2 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_28dflt_LC_11_20_2  (
            .in0(N__72741),
            .in1(N__47477),
            .in2(N__65149),
            .in3(N__72133),
            .lcout(controlWord_28),
            .ltout(controlWord_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_12_LC_11_20_3 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_12_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_12_LC_11_20_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \CONTROL.ramAddReg_12_LC_11_20_3  (
            .in0(N__70461),
            .in1(N__57675),
            .in2(N__28208),
            .in3(N__70762),
            .lcout(A12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_13C_net ),
            .ce(N__70340),
            .sr(_gnd_net_));
    defparam \RAM.un1_WR_105_0_10_LC_11_20_4 .C_ON=1'b0;
    defparam \RAM.un1_WR_105_0_10_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \RAM.un1_WR_105_0_10_LC_11_20_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \RAM.un1_WR_105_0_10_LC_11_20_4  (
            .in0(N__28186),
            .in1(N__44021),
            .in2(_gnd_net_),
            .in3(N__28159),
            .lcout(\RAM.un1_WR_105_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m520_LC_11_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m520_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m520_LC_11_20_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m520_LC_11_20_5  (
            .in0(N__79871),
            .in1(N__44320),
            .in2(N__79529),
            .in3(N__76636),
            .lcout(\PROM.ROMDATA.m520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_29dflt_1_LC_11_20_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_29dflt_1_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_29dflt_1_LC_11_20_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \PROM.ROMDATA.dintern_29dflt_1_LC_11_20_6  (
            .in0(N__79522),
            .in1(N__79872),
            .in2(N__72772),
            .in3(N__72132),
            .lcout(\PROM.ROMDATA.dintern_29dfltZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m514_ns_1_LC_11_20_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m514_ns_1_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m514_ns_1_LC_11_20_7 .LUT_INIT=16'b0000000010000100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m514_ns_1_LC_11_20_7  (
            .in0(N__79870),
            .in1(N__76635),
            .in2(N__79528),
            .in3(N__75985),
            .lcout(\PROM.ROMDATA.m514_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_0_c_LC_11_21_0 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_0_c_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_0_c_LC_11_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \CONTROL.programCounter_1_cry_0_c_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__36728),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\CONTROL.programCounter_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_0_c_RNI26EE1_LC_11_21_1 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_0_c_RNI26EE1_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_0_c_RNI26EE1_LC_11_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_0_c_RNI26EE1_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__29789),
            .in2(_gnd_net_),
            .in3(N__28136),
            .lcout(\CONTROL.programCounter_1_1 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_0 ),
            .carryout(\CONTROL.programCounter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_1_c_RNIRV7S1_LC_11_21_2 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_1_c_RNIRV7S1_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_1_c_RNIRV7S1_LC_11_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_1_c_RNIRV7S1_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__78065),
            .in2(_gnd_net_),
            .in3(N__28133),
            .lcout(\CONTROL.programCounter_1_2 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_1 ),
            .carryout(\CONTROL.programCounter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_2_c_RNIAGGE1_LC_11_21_3 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_2_c_RNIAGGE1_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_2_c_RNIAGGE1_LC_11_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_2_c_RNIAGGE1_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__28271),
            .in2(_gnd_net_),
            .in3(N__28259),
            .lcout(\CONTROL.programCounter_1_3 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_2 ),
            .carryout(\CONTROL.programCounter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_3_c_RNIELHE1_LC_11_21_4 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_3_c_RNIELHE1_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_3_c_RNIELHE1_LC_11_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_3_c_RNIELHE1_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__47330),
            .in2(_gnd_net_),
            .in3(N__28256),
            .lcout(\CONTROL.programCounter_1_4 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_3 ),
            .carryout(\CONTROL.programCounter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_4_c_RNI5AT91_LC_11_21_5 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_4_c_RNI5AT91_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_4_c_RNI5AT91_LC_11_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_4_c_RNI5AT91_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__36743),
            .in2(_gnd_net_),
            .in3(N__28253),
            .lcout(\CONTROL.programCounter_1_5 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_4 ),
            .carryout(\CONTROL.programCounter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_5_c_RNIOM9I1_LC_11_21_6 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_5_c_RNIOM9I1_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_5_c_RNIOM9I1_LC_11_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_5_c_RNIOM9I1_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__79486),
            .in2(_gnd_net_),
            .in3(N__28250),
            .lcout(\CONTROL.programCounter_1_6 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_5 ),
            .carryout(\CONTROL.programCounter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_6_c_RNIDKV91_LC_11_21_7 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_6_c_RNIDKV91_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_6_c_RNIDKV91_LC_11_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_6_c_RNIDKV91_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__72737),
            .in2(_gnd_net_),
            .in3(N__28247),
            .lcout(\CONTROL.programCounter_1_7 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_6 ),
            .carryout(\CONTROL.programCounter_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_7_c_RNIHP0A1_LC_11_22_0 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_7_c_RNIHP0A1_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_7_c_RNIHP0A1_LC_11_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_7_c_RNIHP0A1_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__28376),
            .in2(_gnd_net_),
            .in3(N__28244),
            .lcout(\CONTROL.programCounter_1_8 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\CONTROL.programCounter_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_8_c_RNI39V71_LC_11_22_1 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_8_c_RNI39V71_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_8_c_RNI39V71_LC_11_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_8_c_RNI39V71_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__28547),
            .in2(_gnd_net_),
            .in3(N__28241),
            .lcout(\CONTROL.programCounter_1_9 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_8 ),
            .carryout(\CONTROL.programCounter_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_9_c_RNI67I81_LC_11_22_2 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_9_c_RNI67I81_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_9_c_RNI67I81_LC_11_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_9_c_RNI67I81_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__28440),
            .in2(_gnd_net_),
            .in3(N__28238),
            .lcout(\CONTROL.programCounter_1_10 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_9 ),
            .carryout(\CONTROL.programCounter_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_10_c_RNIHFO21_LC_11_22_3 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_10_c_RNIHFO21_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_10_c_RNIHFO21_LC_11_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_10_c_RNIHFO21_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__30350),
            .in2(_gnd_net_),
            .in3(N__28235),
            .lcout(\CONTROL.programCounter_1_11 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_10 ),
            .carryout(\CONTROL.programCounter_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_11_c_RNIBCO41_LC_11_22_4 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_11_c_RNIBCO41_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_11_c_RNIBCO41_LC_11_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_11_c_RNIBCO41_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__28417),
            .in2(_gnd_net_),
            .in3(N__28355),
            .lcout(\CONTROL.programCounter_1_12 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_11 ),
            .carryout(\CONTROL.programCounter_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_12_c_RNIFHP41_LC_11_22_5 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_12_c_RNIFHP41_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_12_c_RNIFHP41_LC_11_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_12_c_RNIFHP41_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__28309),
            .in2(_gnd_net_),
            .in3(N__28352),
            .lcout(\CONTROL.programCounter_1_13 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_12 ),
            .carryout(\CONTROL.programCounter_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_13_c_RNIJMQ41_LC_11_22_6 .C_ON=1'b1;
    defparam \CONTROL.programCounter_1_cry_13_c_RNIJMQ41_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_13_c_RNIJMQ41_LC_11_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \CONTROL.programCounter_1_cry_13_c_RNIJMQ41_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__28285),
            .in2(_gnd_net_),
            .in3(N__28349),
            .lcout(\CONTROL.programCounter_1_14 ),
            .ltout(),
            .carryin(\CONTROL.programCounter_1_cry_13 ),
            .carryout(\CONTROL.programCounter_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_14_c_RNINRR41_LC_11_22_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_1_cry_14_c_RNINRR41_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_14_c_RNINRR41_LC_11_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CONTROL.programCounter_1_cry_14_c_RNINRR41_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__29740),
            .in2(_gnd_net_),
            .in3(N__28346),
            .lcout(\CONTROL.programCounter_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_13_LC_11_23_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_13_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_13_LC_11_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_1_13_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28342),
            .lcout(\CONTROL.programCounter_1_reto_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73263),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI3EMQ_13_LC_11_23_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI3EMQ_13_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI3EMQ_13_LC_11_23_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI3EMQ_13_LC_11_23_1  (
            .in0(N__28325),
            .in1(N__28319),
            .in2(_gnd_net_),
            .in3(N__42080),
            .lcout(),
            .ltout(\CONTROL.N_428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI7NCV_13_LC_11_23_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI7NCV_13_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI7NCV_13_LC_11_23_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI7NCV_13_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__29822),
            .in2(N__28313),
            .in3(N__28448),
            .lcout(progRomAddress_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIAQCV_14_LC_11_23_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIAQCV_14_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIAQCV_14_LC_11_23_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIAQCV_14_LC_11_23_3  (
            .in0(N__29823),
            .in1(_gnd_net_),
            .in2(N__28295),
            .in3(N__29510),
            .lcout(progRomAddress_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_13_LC_11_23_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_13_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_13_LC_11_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_13_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28463),
            .lcout(\CONTROL.addrstack_reto_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73263),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI8MDT_10_LC_11_23_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI8MDT_10_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI8MDT_10_LC_11_23_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI8MDT_10_LC_11_23_5  (
            .in0(N__28391),
            .in1(N__64619),
            .in2(_gnd_net_),
            .in3(N__29795),
            .lcout(progRomAddress_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI4KCV_12_LC_11_23_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI4KCV_12_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI4KCV_12_LC_11_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI4KCV_12_LC_11_23_6  (
            .in0(N__28424),
            .in1(N__36701),
            .in2(_gnd_net_),
            .in3(N__29821),
            .lcout(progRomAddress_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_10_LC_11_23_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_10_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_10_LC_11_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_10_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28403),
            .lcout(\CONTROL.addrstack_reto_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73263),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_8_LC_11_24_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_8_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_8_LC_11_24_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_8_LC_11_24_0  (
            .in0(N__33586),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73270),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIK8GE_8_LC_11_24_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIK8GE_8_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIK8GE_8_LC_11_24_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIK8GE_8_LC_11_24_1  (
            .in0(N__28385),
            .in1(N__29504),
            .in2(_gnd_net_),
            .in3(N__45121),
            .lcout(N_423),
            .ltout(N_423_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNILCUU_8_LC_11_24_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNILCUU_8_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNILCUU_8_LC_11_24_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNILCUU_8_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__73687),
            .in2(N__28379),
            .in3(N__28538),
            .lcout(\CONTROL.programCounter_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_9_LC_11_24_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_9_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_9_LC_11_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_1_9_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28496),
            .lcout(\CONTROL.programCounter_1_reto_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73270),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_addrstack_0_0_RNO_0_LC_11_24_4 .C_ON=1'b0;
    defparam \CONTROL.addrstack_addrstack_0_0_RNO_0_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_addrstack_0_0_RNO_0_LC_11_24_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \CONTROL.addrstack_addrstack_0_0_RNO_0_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(N__50836),
            .in2(_gnd_net_),
            .in3(N__50903),
            .lcout(\CONTROL.programCounter10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNID2FG_9_LC_11_24_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNID2FG_9_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNID2FG_9_LC_11_24_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CONTROL.programCounter_ret_1_RNID2FG_9_LC_11_24_5  (
            .in0(N__29753),
            .in1(N__28562),
            .in2(_gnd_net_),
            .in3(N__42086),
            .lcout(),
            .ltout(\CONTROL.N_424_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI6QRS_9_LC_11_24_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI6QRS_9_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI6QRS_9_LC_11_24_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI6QRS_9_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__28556),
            .in2(N__28550),
            .in3(N__29824),
            .lcout(progRomAddress_9),
            .ltout(progRomAddress_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_adflt_3_LC_11_24_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_adflt_3_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_adflt_3_LC_11_24_7 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \PROM.ROMDATA.dintern_adflt_3_LC_11_24_7  (
            .in0(N__28537),
            .in1(N__28529),
            .in2(N__28523),
            .in3(N__64655),
            .lcout(\PROM.ROMDATA.dintern_adfltZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_10_LC_11_25_0 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_10_LC_11_25_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_10_LC_11_25_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \CONTROL.tempCounter_10_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(N__29842),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.tempCounterZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_10C_net ),
            .ce(N__34964),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_9_LC_11_25_3 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_9_LC_11_25_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_9_LC_11_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_9_LC_11_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28495),
            .lcout(\CONTROL.tempCounterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_10C_net ),
            .ce(N__34964),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_0_LC_12_7_0 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_0_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_0_LC_12_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CONTROL.addrstackptr_0_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__57728),
            .in2(_gnd_net_),
            .in3(N__41990),
            .lcout(\CONTROL.addrstack_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.addrstackptr_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNINS3U7_0_LC_12_8_0 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNINS3U7_0_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNINS3U7_0_LC_12_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.busState_1_RNINS3U7_0_LC_12_8_0  (
            .in0(N__33101),
            .in1(N__28640),
            .in2(_gnd_net_),
            .in3(N__49817),
            .lcout(bus_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN3QUB1_0_2_LC_12_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNIN3QUB1_0_2_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN3QUB1_0_2_LC_12_8_1 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.d_RNIN3QUB1_0_2_LC_12_8_1  (
            .in0(N__66602),
            .in1(N__66312),
            .in2(N__60263),
            .in3(N__65951),
            .lcout(\ALU.rshift_3_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5SIF41_4_LC_12_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNI5SIF41_4_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5SIF41_4_LC_12_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI5SIF41_4_LC_12_8_2  (
            .in0(N__59586),
            .in1(N__59874),
            .in2(N__56268),
            .in3(N__56115),
            .lcout(\ALU.d_RNI5SIF41Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_1_c_RNO_LC_12_8_4 .C_ON=1'b0;
    defparam \ALU.status_17_I_1_c_RNO_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_1_c_RNO_LC_12_8_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \ALU.status_17_I_1_c_RNO_LC_12_8_4  (
            .in0(N__65952),
            .in1(N__65570),
            .in2(N__60629),
            .in3(N__66603),
            .lcout(\ALU.status_17_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0PI3E1_8_LC_12_9_0 .C_ON=1'b0;
    defparam \ALU.d_RNI0PI3E1_8_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0PI3E1_8_LC_12_9_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNI0PI3E1_8_LC_12_9_0  (
            .in0(N__65965),
            .in1(N__62874),
            .in2(N__61976),
            .in3(N__68823),
            .lcout(\ALU.d_RNI0PI3E1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFGGBO_6_LC_12_9_1 .C_ON=1'b0;
    defparam \ALU.d_RNIFGGBO_6_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFGGBO_6_LC_12_9_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ALU.d_RNIFGGBO_6_LC_12_9_1  (
            .in0(N__62273),
            .in1(_gnd_net_),
            .in2(N__62585),
            .in3(N__66601),
            .lcout(),
            .ltout(\ALU.N_834_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMQD952_6_LC_12_9_2 .C_ON=1'b0;
    defparam \ALU.d_RNIMQD952_6_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMQD952_6_LC_12_9_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNIMQD952_6_LC_12_9_2  (
            .in0(N__65963),
            .in1(_gnd_net_),
            .in2(N__28586),
            .in3(N__42772),
            .lcout(\ALU.N_864 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIUFQIG_7_LC_12_9_3 .C_ON=1'b0;
    defparam \ALU.d_RNIUFQIG_7_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIUFQIG_7_LC_12_9_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIUFQIG_7_LC_12_9_3  (
            .in0(N__62271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68256),
            .lcout(\ALU.d_RNIUFQIGZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC6EBM2_2_LC_12_9_5 .C_ON=1'b0;
    defparam \ALU.d_RNIC6EBM2_2_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC6EBM2_2_LC_12_9_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \ALU.d_RNIC6EBM2_2_LC_12_9_5  (
            .in0(N__68824),
            .in1(N__47985),
            .in2(N__45723),
            .in3(N__65964),
            .lcout(\ALU.d_RNIC6EBM2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITLGIL_7_LC_12_9_6 .C_ON=1'b0;
    defparam \ALU.d_RNITLGIL_7_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITLGIL_7_LC_12_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNITLGIL_7_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__62270),
            .in2(_gnd_net_),
            .in3(N__68822),
            .lcout(\ALU.d_RNITLGILZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIB692D1_6_LC_12_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNIB692D1_6_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIB692D1_6_LC_12_9_7 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.d_RNIB692D1_6_LC_12_9_7  (
            .in0(N__62272),
            .in1(N__65962),
            .in2(N__62584),
            .in3(N__66600),
            .lcout(\ALU.mult_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISRIE42_2_LC_12_10_0 .C_ON=1'b0;
    defparam \ALU.d_RNISRIE42_2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISRIE42_2_LC_12_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALU.d_RNISRIE42_2_LC_12_10_0  (
            .in0(N__66653),
            .in1(N__68940),
            .in2(N__68280),
            .in3(N__66010),
            .lcout(\ALU.lshift62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9OBVC_3_LC_12_10_1 .C_ON=1'b0;
    defparam \ALU.d_RNI9OBVC_3_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9OBVC_3_LC_12_10_1 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \ALU.d_RNI9OBVC_3_LC_12_10_1  (
            .in0(N__38065),
            .in1(N__28583),
            .in2(N__53288),
            .in3(N__34586),
            .lcout(\ALU.status_19_2 ),
            .ltout(\ALU.status_19_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJBM6G_3_LC_12_10_2 .C_ON=1'b0;
    defparam \ALU.d_RNIJBM6G_3_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJBM6G_3_LC_12_10_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNIJBM6G_3_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28661),
            .in3(N__60197),
            .lcout(\ALU.d_RNIJBM6GZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFBJI61_0_LC_12_10_3 .C_ON=1'b0;
    defparam \ALU.d_RNIFBJI61_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFBJI61_0_LC_12_10_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNIFBJI61_0_LC_12_10_3  (
            .in0(N__68941),
            .in1(N__65550),
            .in2(N__60628),
            .in3(N__68231),
            .lcout(\ALU.d_RNIFBJI61Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITK2D51_2_LC_12_10_4 .C_ON=1'b0;
    defparam \ALU.d_RNITK2D51_2_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITK2D51_2_LC_12_10_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNITK2D51_2_LC_12_10_4  (
            .in0(N__68232),
            .in1(N__66288),
            .in2(N__60264),
            .in3(N__68942),
            .lcout(\ALU.d_RNITK2D51Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI04H8G_3_LC_12_10_5 .C_ON=1'b0;
    defparam \ALU.d_RNI04H8G_3_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI04H8G_3_LC_12_10_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.d_RNI04H8G_3_LC_12_10_5  (
            .in0(N__60198),
            .in1(N__63289),
            .in2(_gnd_net_),
            .in3(N__68233),
            .lcout(\ALU.d_RNI04H8GZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI7U266_2_LC_12_10_7 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI7U266_2_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI7U266_2_LC_12_10_7 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \CONTROL.busState_1_RNI7U266_2_LC_12_10_7  (
            .in0(N__59865),
            .in1(N__49605),
            .in2(N__28658),
            .in3(N__50221),
            .lcout(\CONTROL.busState_1_RNI7U266Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_95_c_LC_12_11_0 .C_ON=1'b1;
    defparam \ALU.mult_95_c_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_95_c_LC_12_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_95_c_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__34046),
            .in2(N__28847),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\ALU.mult_3_c3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_95_c_RNINLQ452_LC_12_11_1 .C_ON=1'b1;
    defparam \ALU.mult_95_c_RNINLQ452_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_95_c_RNINLQ452_LC_12_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_95_c_RNINLQ452_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__30206),
            .in2(N__28859),
            .in3(N__28631),
            .lcout(\ALU.mult_3_4 ),
            .ltout(),
            .carryin(\ALU.mult_3_c3 ),
            .carryout(\ALU.mult_3_c4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_101_c_RNIKJVKQ1_LC_12_11_2 .C_ON=1'b1;
    defparam \ALU.mult_101_c_RNIKJVKQ1_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_101_c_RNIKJVKQ1_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_101_c_RNIKJVKQ1_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__30245),
            .in2(N__28628),
            .in3(N__28619),
            .lcout(\ALU.mult_3_5 ),
            .ltout(),
            .carryin(\ALU.mult_3_c4 ),
            .carryout(\ALU.mult_3_c5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_107_c_RNIILDTH1_LC_12_11_3 .C_ON=1'b1;
    defparam \ALU.mult_107_c_RNIILDTH1_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_107_c_RNIILDTH1_LC_12_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_107_c_RNIILDTH1_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__28616),
            .in2(N__28610),
            .in3(N__28601),
            .lcout(\ALU.mult_3_6 ),
            .ltout(),
            .carryin(\ALU.mult_3_c5 ),
            .carryout(\ALU.mult_3_c6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_113_c_RNIH8VLK1_LC_12_11_4 .C_ON=1'b1;
    defparam \ALU.mult_113_c_RNIH8VLK1_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_113_c_RNIH8VLK1_LC_12_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_113_c_RNIH8VLK1_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__28790),
            .in2(N__28784),
            .in3(N__28772),
            .lcout(\ALU.mult_3_7 ),
            .ltout(),
            .carryin(\ALU.mult_3_c6 ),
            .carryout(\ALU.mult_3_c7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_119_c_RNI03FQK1_LC_12_11_5 .C_ON=1'b1;
    defparam \ALU.mult_119_c_RNI03FQK1_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_119_c_RNI03FQK1_LC_12_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_119_c_RNI03FQK1_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__28769),
            .in2(N__28763),
            .in3(N__28754),
            .lcout(\ALU.mult_3_8 ),
            .ltout(),
            .carryin(\ALU.mult_3_c7 ),
            .carryout(\ALU.mult_3_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_125_c_RNI84ENI1_LC_12_11_6 .C_ON=1'b1;
    defparam \ALU.mult_125_c_RNI84ENI1_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_125_c_RNI84ENI1_LC_12_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_125_c_RNI84ENI1_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__28751),
            .in2(N__28745),
            .in3(N__28736),
            .lcout(\ALU.mult_3_9 ),
            .ltout(),
            .carryin(\ALU.mult_3_c8 ),
            .carryout(\ALU.mult_3_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_131_c_RNICCA4H1_LC_12_11_7 .C_ON=1'b1;
    defparam \ALU.mult_131_c_RNICCA4H1_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_131_c_RNICCA4H1_LC_12_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_131_c_RNICCA4H1_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__28733),
            .in2(N__28808),
            .in3(N__28727),
            .lcout(\ALU.mult_3_10 ),
            .ltout(),
            .carryin(\ALU.mult_3_c9 ),
            .carryout(\ALU.mult_3_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_137_c_RNI7M9PJ1_LC_12_12_0 .C_ON=1'b1;
    defparam \ALU.mult_137_c_RNI7M9PJ1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_137_c_RNI7M9PJ1_LC_12_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_137_c_RNI7M9PJ1_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__28724),
            .in2(N__28820),
            .in3(N__28715),
            .lcout(\ALU.mult_3_11 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\ALU.mult_3_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_143_c_RNIUMAAM1_LC_12_12_1 .C_ON=1'b1;
    defparam \ALU.mult_143_c_RNIUMAAM1_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_143_c_RNIUMAAM1_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_143_c_RNIUMAAM1_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__28712),
            .in2(N__28700),
            .in3(N__28685),
            .lcout(\ALU.mult_3_12 ),
            .ltout(),
            .carryin(\ALU.mult_3_c11 ),
            .carryout(\ALU.mult_3_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_149_c_RNIK33CN1_LC_12_12_2 .C_ON=1'b1;
    defparam \ALU.mult_149_c_RNIK33CN1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_149_c_RNIK33CN1_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_149_c_RNIK33CN1_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__28682),
            .in2(N__28829),
            .in3(N__28667),
            .lcout(\ALU.mult_3_13 ),
            .ltout(),
            .carryin(\ALU.mult_3_c12 ),
            .carryout(\ALU.mult_3_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_155_c_RNI2IBOL1_LC_12_12_3 .C_ON=1'b1;
    defparam \ALU.mult_155_c_RNI2IBOL1_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_155_c_RNI2IBOL1_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_155_c_RNI2IBOL1_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__28796),
            .in2(N__28964),
            .in3(N__28664),
            .lcout(\ALU.mult_3_14 ),
            .ltout(),
            .carryin(\ALU.mult_3_c13 ),
            .carryout(\ALU.mult_3_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_3_c14_THRU_LUT4_0_LC_12_12_4 .C_ON=1'b0;
    defparam \ALU.mult_3_c14_THRU_LUT4_0_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_3_c14_THRU_LUT4_0_LC_12_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.mult_3_c14_THRU_LUT4_0_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28832),
            .lcout(\ALU.mult_3_c14_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9E4F21_4_LC_12_12_5 .C_ON=1'b0;
    defparam \ALU.d_RNI9E4F21_4_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9E4F21_4_LC_12_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI9E4F21_4_LC_12_12_5  (
            .in0(N__55800),
            .in1(N__59588),
            .in2(N__55990),
            .in3(N__59833),
            .lcout(\ALU.d_RNI9E4F21Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIH49MH_1_LC_12_12_6 .C_ON=1'b0;
    defparam \ALU.d_RNIH49MH_1_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIH49MH_1_LC_12_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIH49MH_1_LC_12_12_6  (
            .in0(N__65543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55799),
            .lcout(\ALU.d_RNIH49MHZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRJ3VH_1_LC_12_12_7 .C_ON=1'b0;
    defparam \ALU.d_RNIRJ3VH_1_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRJ3VH_1_LC_12_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIRJ3VH_1_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__65542),
            .in2(_gnd_net_),
            .in3(N__56086),
            .lcout(\ALU.d_RNIRJ3VHZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI371041_8_LC_12_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNI371041_8_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI371041_8_LC_12_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI371041_8_LC_12_13_1  (
            .in0(N__62845),
            .in1(N__56116),
            .in2(N__56272),
            .in3(N__61901),
            .lcout(\ALU.d_RNI371041Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2IA441_2_LC_12_13_3 .C_ON=1'b0;
    defparam \ALU.d_RNI2IA441_2_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2IA441_2_LC_12_13_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.d_RNI2IA441_2_LC_12_13_3  (
            .in0(N__66249),
            .in1(N__60213),
            .in2(N__57029),
            .in3(N__55577),
            .lcout(\ALU.d_RNI2IA441Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7SQI21_2_LC_12_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNI7SQI21_2_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7SQI21_2_LC_12_13_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI7SQI21_2_LC_12_13_4  (
            .in0(N__55674),
            .in1(N__60209),
            .in2(N__55823),
            .in3(N__66248),
            .lcout(\ALU.d_RNI7SQI21Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIK8R951_0_LC_12_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNIK8R951_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIK8R951_0_LC_12_13_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.d_RNIK8R951_0_LC_12_13_5  (
            .in0(N__60598),
            .in1(N__65493),
            .in2(N__57028),
            .in3(N__55578),
            .lcout(\ALU.d_RNIK8R951Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID31VF_3_LC_12_13_6 .C_ON=1'b0;
    defparam \ALU.d_RNID31VF_3_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID31VF_3_LC_12_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNID31VF_3_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__60208),
            .in2(_gnd_net_),
            .in3(N__55957),
            .lcout(\ALU.d_RNID31VFZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBRFE41_2_LC_12_13_7 .C_ON=1'b0;
    defparam \ALU.d_RNIBRFE41_2_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBRFE41_2_LC_12_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIBRFE41_2_LC_12_13_7  (
            .in0(N__66250),
            .in1(N__60214),
            .in2(N__57030),
            .in3(N__56905),
            .lcout(\ALU.d_RNIBRFE41Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN3H0D_3_LC_12_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNIN3H0D_3_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN3H0D_3_LC_12_14_1 .LUT_INIT=16'b1000000010110000;
    LogicCell40 \ALU.d_RNIN3H0D_3_LC_12_14_1  (
            .in0(N__33058),
            .in1(N__53165),
            .in2(N__70012),
            .in3(N__38066),
            .lcout(\ALU.d_RNIN3H0DZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9IN2H_3_LC_12_14_2 .C_ON=1'b0;
    defparam \ALU.d_RNI9IN2H_3_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9IN2H_3_LC_12_14_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI9IN2H_3_LC_12_14_2  (
            .in0(N__60101),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57015),
            .lcout(\ALU.d_RNI9IN2HZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRD18N_2_LC_12_14_3 .C_ON=1'b0;
    defparam \ALU.d_RNIRD18N_2_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRD18N_2_LC_12_14_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNIRD18N_2_LC_12_14_3  (
            .in0(N__60118),
            .in1(N__66251),
            .in2(_gnd_net_),
            .in3(N__66377),
            .lcout(\ALU.N_767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI2N741_12_LC_12_14_4 .C_ON=1'b0;
    defparam \ALU.a_RNI2N741_12_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI2N741_12_LC_12_14_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.a_RNI2N741_12_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__48269),
            .in2(N__51421),
            .in3(N__43309),
            .lcout(\ALU.a_RNI2N741Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILEAFE_0_5_LC_12_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNILEAFE_0_5_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILEAFE_0_5_LC_12_14_5 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \ALU.d_RNILEAFE_0_5_LC_12_14_5  (
            .in0(N__40594),
            .in1(N__28940),
            .in2(N__28922),
            .in3(N__28877),
            .lcout(\ALU.combOperand2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI693UN_3_LC_12_14_6 .C_ON=1'b0;
    defparam \ALU.d_RNI693UN_3_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI693UN_3_LC_12_14_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI693UN_3_LC_12_14_6  (
            .in0(N__60100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65929),
            .lcout(\ALU.d_RNI693UNZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_95_c_RNO_0_LC_12_14_7 .C_ON=1'b0;
    defparam \ALU.mult_95_c_RNO_0_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_95_c_RNO_0_LC_12_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_95_c_RNO_0_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__60099),
            .in2(_gnd_net_),
            .in3(N__66376),
            .lcout(\ALU.mult_95_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI42AE1_11_LC_12_15_0 .C_ON=1'b0;
    defparam \ALU.b_RNI42AE1_11_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI42AE1_11_LC_12_15_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI42AE1_11_LC_12_15_0  (
            .in0(N__39841),
            .in1(N__47284),
            .in2(N__35968),
            .in3(N__54304),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI88772_11_LC_12_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNI88772_11_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI88772_11_LC_12_15_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNI88772_11_LC_12_15_1  (
            .in0(N__57981),
            .in1(N__36188),
            .in2(N__28835),
            .in3(N__47210),
            .lcout(\ALU.N_1144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI2TJC1_11_LC_12_15_2 .C_ON=1'b0;
    defparam \ALU.b_RNI2TJC1_11_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI2TJC1_11_LC_12_15_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.b_RNI2TJC1_11_LC_12_15_2  (
            .in0(N__39842),
            .in1(_gnd_net_),
            .in2(N__35969),
            .in3(N__43310),
            .lcout(\ALU.b_RNI2TJC1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI4OEM1_11_LC_12_15_3 .C_ON=1'b0;
    defparam \ALU.c_RNI4OEM1_11_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI4OEM1_11_LC_12_15_3 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \ALU.c_RNI4OEM1_11_LC_12_15_3  (
            .in0(N__36104),
            .in1(N__29081),
            .in2(N__35671),
            .in3(N__47211),
            .lcout(),
            .ltout(\ALU.N_1096_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIF4474_11_LC_12_15_4 .C_ON=1'b0;
    defparam \ALU.c_RNIF4474_11_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIF4474_11_LC_12_15_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.c_RNIF4474_11_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__29015),
            .in2(N__29009),
            .in3(N__54142),
            .lcout(aluOut_11),
            .ltout(aluOut_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNICV1S5_1_LC_12_15_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNICV1S5_1_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNICV1S5_1_LC_12_15_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \CONTROL.busState_1_RNICV1S5_1_LC_12_15_5  (
            .in0(N__29006),
            .in1(N__50341),
            .in2(N__28994),
            .in3(N__50219),
            .lcout(N_204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBH5A2_11_LC_12_16_0 .C_ON=1'b0;
    defparam \ALU.c_RNIBH5A2_11_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBH5A2_11_LC_12_16_0 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.c_RNIBH5A2_11_LC_12_16_0  (
            .in0(N__29087),
            .in1(N__53936),
            .in2(N__28973),
            .in3(N__46836),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN5325_11_LC_12_16_1 .C_ON=1'b0;
    defparam \ALU.d_RNIN5325_11_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN5325_11_LC_12_16_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIN5325_11_LC_12_16_1  (
            .in0(N__53937),
            .in1(N__36170),
            .in2(N__28991),
            .in3(N__28988),
            .lcout(),
            .ltout(\ALU.operand2_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMR627_11_LC_12_16_2 .C_ON=1'b0;
    defparam \ALU.d_RNIMR627_11_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMR627_11_LC_12_16_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.d_RNIMR627_11_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__30677),
            .in2(N__28979),
            .in3(N__71399),
            .lcout(),
            .ltout(\ALU.d_RNIMR627Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVUCRD_11_LC_12_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNIVUCRD_11_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVUCRD_11_LC_12_16_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ALU.d_RNIVUCRD_11_LC_12_16_3  (
            .in0(N__30664),
            .in1(N__53161),
            .in2(N__28976),
            .in3(N__49588),
            .lcout(\ALU.status_19_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIV5PU_11_LC_12_16_4 .C_ON=1'b0;
    defparam \ALU.a_RNIV5PU_11_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIV5PU_11_LC_12_16_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.a_RNIV5PU_11_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__46935),
            .in2(N__37265),
            .in3(N__32599),
            .lcout(\ALU.a_RNIV5PUZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3MHF_11_LC_12_16_5 .C_ON=1'b0;
    defparam \ALU.c_RNI3MHF_11_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3MHF_11_LC_12_16_5 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \ALU.c_RNI3MHF_11_LC_12_16_5  (
            .in0(N__35664),
            .in1(N__36103),
            .in2(N__46945),
            .in3(_gnd_net_),
            .lcout(\ALU.c_RNI3MHFZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI2QT51_11_LC_12_16_6 .C_ON=1'b0;
    defparam \ALU.a_RNI2QT51_11_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI2QT51_11_LC_12_16_6 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.a_RNI2QT51_11_LC_12_16_6  (
            .in0(N__37261),
            .in1(N__47285),
            .in2(N__32606),
            .in3(N__54303),
            .lcout(\ALU.dout_3_ns_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNICADA1_10_LC_12_17_0 .C_ON=1'b0;
    defparam \ALU.a_RNICADA1_10_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNICADA1_10_LC_12_17_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.a_RNICADA1_10_LC_12_17_0  (
            .in0(N__37075),
            .in1(N__36338),
            .in2(N__32636),
            .in3(N__32822),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBCLN1_10_LC_12_17_1 .C_ON=1'b0;
    defparam \ALU.c_RNIBCLN1_10_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBCLN1_10_LC_12_17_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNIBCLN1_10_LC_12_17_1  (
            .in0(N__35712),
            .in1(N__36137),
            .in2(N__29075),
            .in3(N__54292),
            .lcout(\ALU.N_1095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIEIPI1_10_LC_12_17_2 .C_ON=1'b0;
    defparam \ALU.b_RNIEIPI1_10_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIEIPI1_10_LC_12_17_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.b_RNIEIPI1_10_LC_12_17_2  (
            .in0(N__39133),
            .in1(N__36339),
            .in2(N__36004),
            .in3(N__32823),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFSD82_10_LC_12_17_3 .C_ON=1'b0;
    defparam \ALU.d_RNIFSD82_10_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFSD82_10_LC_12_17_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIFSD82_10_LC_12_17_3  (
            .in0(N__58227),
            .in1(N__36035),
            .in2(N__29072),
            .in3(N__54293),
            .lcout(),
            .ltout(\ALU.N_1143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNITCH94_10_LC_12_17_4 .C_ON=1'b0;
    defparam \ALU.c_RNITCH94_10_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNITCH94_10_LC_12_17_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.c_RNITCH94_10_LC_12_17_4  (
            .in0(N__54128),
            .in1(_gnd_net_),
            .in2(N__29069),
            .in3(N__29066),
            .lcout(aluOut_10),
            .ltout(aluOut_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIDR6R7_0_LC_12_17_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIDR6R7_0_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIDR6R7_0_LC_12_17_5 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \CONTROL.busState_1_RNIDR6R7_0_LC_12_17_5  (
            .in0(N__30833),
            .in1(N__34482),
            .in2(N__29060),
            .in3(N__49785),
            .lcout(\CONTROL.bus_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILM2O3_8_LC_12_17_7 .C_ON=1'b0;
    defparam \ALU.d_RNILM2O3_8_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILM2O3_8_LC_12_17_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNILM2O3_8_LC_12_17_7  (
            .in0(N__29033),
            .in1(N__54129),
            .in2(_gnd_net_),
            .in3(N__29027),
            .lcout(aluOut_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.combOperand2_d_bm_7_LC_12_18_0 .C_ON=1'b0;
    defparam \ALU.combOperand2_d_bm_7_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \ALU.combOperand2_d_bm_7_LC_12_18_0 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \ALU.combOperand2_d_bm_7_LC_12_18_0  (
            .in0(N__29183),
            .in1(N__49532),
            .in2(N__29174),
            .in3(N__50124),
            .lcout(\ALU.combOperand2_d_bmZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_7_LC_12_18_1 .C_ON=1'b0;
    defparam \CONTROL.dout_7_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_7_LC_12_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \CONTROL.dout_7_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__29141),
            .in2(_gnd_net_),
            .in3(N__72101),
            .lcout(\CONTROL.ctrlOut_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_7C_net ),
            .ce(N__44452),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNIAQOJ_7_LC_12_18_2 .C_ON=1'b0;
    defparam \CONTROL.dout_RNIAQOJ_7_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNIAQOJ_7_LC_12_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNIAQOJ_7_LC_12_18_2  (
            .in0(N__29204),
            .in1(N__33391),
            .in2(_gnd_net_),
            .in3(N__50123),
            .lcout(N_168),
            .ltout(N_168_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI77OM1_2_LC_12_18_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI77OM1_2_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI77OM1_2_LC_12_18_3 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \CONTROL.busState_1_RNI77OM1_2_LC_12_18_3  (
            .in0(N__50126),
            .in1(N__49544),
            .in2(N__29177),
            .in3(N__29173),
            .lcout(),
            .ltout(\CONTROL.bus_7_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNITSIT7_0_LC_12_18_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNITSIT7_0_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNITSIT7_0_LC_12_18_4 .LUT_INIT=16'b0010011100000101;
    LogicCell40 \CONTROL.busState_1_RNITSIT7_0_LC_12_18_4  (
            .in0(N__49711),
            .in1(N__49534),
            .in2(N__29144),
            .in3(N__43769),
            .lcout(bus_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_23dflt_LC_12_18_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_23dflt_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_23dflt_LC_12_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PROM.ROMDATA.dintern_23dflt_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__29140),
            .in2(_gnd_net_),
            .in3(N__72100),
            .lcout(controlWord_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIP3P31_0_LC_12_18_6 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIP3P31_0_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIP3P31_0_LC_12_18_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \CONTROL.busState_1_RNIP3P31_0_LC_12_18_6  (
            .in0(N__49709),
            .in1(N__49533),
            .in2(_gnd_net_),
            .in3(N__50125),
            .lcout(\CONTROL.bus_7_a1_1_8 ),
            .ltout(\CONTROL.bus_7_a1_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIA1EN6_0_LC_12_18_7 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIA1EN6_0_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIA1EN6_0_LC_12_18_7 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \CONTROL.busState_1_RNIA1EN6_0_LC_12_18_7  (
            .in0(N__33167),
            .in1(N__61836),
            .in2(N__29123),
            .in3(N__49710),
            .lcout(\CONTROL.bus_sx_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_2_LC_12_19_0 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_2_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_2_LC_12_19_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.gpuAddReg_2_LC_12_19_0  (
            .in0(N__29597),
            .in1(N__70708),
            .in2(N__34399),
            .in3(N__70458),
            .lcout(gpuAddress_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_2C_net ),
            .ce(N__30759),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_3_LC_12_19_1 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_3_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_3_LC_12_19_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \CONTROL.gpuAddReg_3_LC_12_19_1  (
            .in0(N__70455),
            .in1(N__58610),
            .in2(N__70764),
            .in3(N__44255),
            .lcout(gpuAddress_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_2C_net ),
            .ce(N__30759),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_4_LC_12_19_2 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_4_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_4_LC_12_19_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \CONTROL.gpuAddReg_4_LC_12_19_2  (
            .in0(N__70514),
            .in1(N__70709),
            .in2(N__43403),
            .in3(N__44188),
            .lcout(gpuAddress_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_2C_net ),
            .ce(N__30759),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_5_LC_12_19_3 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_5_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_5_LC_12_19_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \CONTROL.gpuAddReg_5_LC_12_19_3  (
            .in0(N__70456),
            .in1(N__29455),
            .in2(N__70765),
            .in3(N__40268),
            .lcout(gpuAddress_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_2C_net ),
            .ce(N__30759),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_6_LC_12_19_4 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_6_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_6_LC_12_19_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.gpuAddReg_6_LC_12_19_4  (
            .in0(N__70828),
            .in1(N__70710),
            .in2(N__37445),
            .in3(N__70459),
            .lcout(gpuAddress_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_2C_net ),
            .ce(N__30759),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_7_LC_12_19_5 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_7_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_7_LC_12_19_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \CONTROL.gpuAddReg_7_LC_12_19_5  (
            .in0(N__70457),
            .in1(N__43835),
            .in2(N__70766),
            .in3(N__29368),
            .lcout(gpuAddress_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_2C_net ),
            .ce(N__30759),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuAddReg_8_LC_12_19_6 .C_ON=1'b0;
    defparam \CONTROL.gpuAddReg_8_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuAddReg_8_LC_12_19_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.gpuAddReg_8_LC_12_19_6  (
            .in0(N__31084),
            .in1(N__70711),
            .in2(N__48146),
            .in3(N__70460),
            .lcout(gpuAddress_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuAddReg_2C_net ),
            .ce(N__30759),
            .sr(_gnd_net_));
    defparam \CONTROL.ramWrite_5_m9_0_a2_0_LC_12_20_0 .C_ON=1'b0;
    defparam \CONTROL.ramWrite_5_m9_0_a2_0_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.ramWrite_5_m9_0_a2_0_LC_12_20_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \CONTROL.ramWrite_5_m9_0_a2_0_LC_12_20_0  (
            .in0(N__38597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30790),
            .lcout(\CONTROL.N_346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuWrite_RNO_3_LC_12_20_1 .C_ON=1'b0;
    defparam \CONTROL.gpuWrite_RNO_3_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.gpuWrite_RNO_3_LC_12_20_1 .LUT_INIT=16'b1000100011000100;
    LogicCell40 \CONTROL.gpuWrite_RNO_3_LC_12_20_1  (
            .in0(N__41430),
            .in1(N__41241),
            .in2(N__36404),
            .in3(N__54688),
            .lcout(),
            .ltout(\CONTROL.un1_busState119_1_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuWrite_RNO_1_LC_12_20_2 .C_ON=1'b0;
    defparam \CONTROL.gpuWrite_RNO_1_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.gpuWrite_RNO_1_LC_12_20_2 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \CONTROL.gpuWrite_RNO_1_LC_12_20_2  (
            .in0(N__41596),
            .in1(_gnd_net_),
            .in2(N__29207),
            .in3(N__54746),
            .lcout(\CONTROL.N_66_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuWrite_RNO_2_LC_12_20_3 .C_ON=1'b0;
    defparam \CONTROL.gpuWrite_RNO_2_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.gpuWrite_RNO_2_LC_12_20_3 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \CONTROL.gpuWrite_RNO_2_LC_12_20_3  (
            .in0(N__31462),
            .in1(N__38595),
            .in2(N__41698),
            .in3(N__41595),
            .lcout(),
            .ltout(\CONTROL.gpuWrite_RNOZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuWrite_RNO_0_LC_12_20_4 .C_ON=1'b0;
    defparam \CONTROL.gpuWrite_RNO_0_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.gpuWrite_RNO_0_LC_12_20_4 .LUT_INIT=16'b0010000000110000;
    LogicCell40 \CONTROL.gpuWrite_RNO_0_LC_12_20_4  (
            .in0(N__38596),
            .in1(N__38324),
            .in2(N__29498),
            .in3(N__30789),
            .lcout(\CONTROL.gpuWrite_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState101_3_0_a2_1_LC_12_20_5 .C_ON=1'b0;
    defparam \CONTROL.un1_busState101_3_0_a2_1_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState101_3_0_a2_1_LC_12_20_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \CONTROL.un1_busState101_3_0_a2_1_LC_12_20_5  (
            .in0(N__54687),
            .in1(N__44899),
            .in2(N__44773),
            .in3(N__44714),
            .lcout(\CONTROL.busState96 ),
            .ltout(\CONTROL.busState96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState101_3_0_1_LC_12_20_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState101_3_0_1_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState101_3_0_1_LC_12_20_6 .LUT_INIT=16'b0000010100001111;
    LogicCell40 \CONTROL.un1_busState101_3_0_1_LC_12_20_6  (
            .in0(N__36605),
            .in1(_gnd_net_),
            .in2(N__29495),
            .in3(N__36494),
            .lcout(\CONTROL.un1_busState101_3_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.gpuWrite_LC_12_20_7 .C_ON=1'b0;
    defparam \CONTROL.gpuWrite_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.gpuWrite_LC_12_20_7 .LUT_INIT=16'b0100000001010001;
    LogicCell40 \CONTROL.gpuWrite_LC_12_20_7  (
            .in0(N__29492),
            .in1(N__29486),
            .in2(N__29473),
            .in3(N__29480),
            .lcout(gpuWrite),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.gpuWriteC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_5_LC_12_21_1 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_5_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_5_LC_12_21_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.ramAddReg_5_LC_12_21_1  (
            .in0(N__39986),
            .in1(N__70722),
            .in2(N__29456),
            .in3(N__70467),
            .lcout(A5_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_5C_net ),
            .ce(N__70317),
            .sr(_gnd_net_));
    defparam \RAM.un1_WR_105_0_3_LC_12_21_2 .C_ON=1'b0;
    defparam \RAM.un1_WR_105_0_3_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \RAM.un1_WR_105_0_3_LC_12_21_2 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \RAM.un1_WR_105_0_3_LC_12_21_2  (
            .in0(N__29557),
            .in1(N__29344),
            .in2(_gnd_net_),
            .in3(N__31294),
            .lcout(),
            .ltout(\RAM.un1_WR_105_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RAM.un1_WR_105_0_11_LC_12_21_3 .C_ON=1'b0;
    defparam \RAM.un1_WR_105_0_11_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \RAM.un1_WR_105_0_11_LC_12_21_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \RAM.un1_WR_105_0_11_LC_12_21_3  (
            .in0(N__70369),
            .in1(N__31151),
            .in2(N__29417),
            .in3(N__29398),
            .lcout(\RAM.un1_WR_105_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_7_LC_12_21_5 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_7_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_7_LC_12_21_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.ramAddReg_7_LC_12_21_5  (
            .in0(N__29369),
            .in1(N__70723),
            .in2(N__49091),
            .in3(N__70468),
            .lcout(A7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_5C_net ),
            .ce(N__70317),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_18dflt_LC_12_21_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_18dflt_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_18dflt_LC_12_21_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_18dflt_LC_12_21_6  (
            .in0(N__45767),
            .in1(N__72775),
            .in2(N__41012),
            .in3(N__72131),
            .lcout(controlWord_18),
            .ltout(controlWord_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_2_LC_12_21_7 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_2_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_2_LC_12_21_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.ramAddReg_2_LC_12_21_7  (
            .in0(N__35636),
            .in1(N__70721),
            .in2(N__29579),
            .in3(N__70466),
            .lcout(A2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_5C_net ),
            .ce(N__70317),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_4_LC_12_22_0 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_4_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_4_LC_12_22_0 .LUT_INIT=16'b1001111111111111;
    LogicCell40 \CONTROL.g0_3_i_4_LC_12_22_0  (
            .in0(N__42266),
            .in1(N__54659),
            .in2(N__72315),
            .in3(N__55471),
            .lcout(),
            .ltout(\CONTROL.g0_3_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIFRI6PV_7_LC_12_22_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIFRI6PV_7_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIFRI6PV_7_LC_12_22_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIFRI6PV_7_LC_12_22_1  (
            .in0(N__29516),
            .in1(N__38501),
            .in2(N__29546),
            .in3(N__38186),
            .lcout(\CONTROL.N_4_1 ),
            .ltout(\CONTROL.N_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_4_LC_12_22_2 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_4_LC_12_22_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_4_LC_12_22_2 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \CONTROL.addrstackptr_4_LC_12_22_2  (
            .in0(N__29708),
            .in1(N__60780),
            .in2(N__29543),
            .in3(N__29675),
            .lcout(\CONTROL.addrstackptrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.addrstackptr_4C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI1MMTM91_3_LC_12_22_3 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI1MMTM91_3_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI1MMTM91_3_LC_12_22_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI1MMTM91_3_LC_12_22_3  (
            .in0(N__41977),
            .in1(N__34772),
            .in2(N__31481),
            .in3(N__60730),
            .lcout(\CONTROL.un1_addrstackptr_c4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_7_174_i_i_o2_LC_12_22_4 .C_ON=1'b0;
    defparam \CONTROL.aluParams_7_174_i_i_o2_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluParams_7_174_i_i_o2_LC_12_22_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \CONTROL.aluParams_7_174_i_i_o2_LC_12_22_4  (
            .in0(N__44701),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54657),
            .lcout(\CONTROL.N_81_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_a7_LC_12_22_6 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_a7_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_a7_LC_12_22_6 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \CONTROL.g0_3_i_a7_LC_12_22_6  (
            .in0(N__45221),
            .in1(N__54658),
            .in2(N__63481),
            .in3(N__38273),
            .lcout(\CONTROL.g0_3_i_a7_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI5GMQ_14_LC_12_23_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI5GMQ_14_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI5GMQ_14_LC_12_23_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI5GMQ_14_LC_12_23_0  (
            .in0(N__29603),
            .in1(N__29633),
            .in2(_gnd_net_),
            .in3(N__42081),
            .lcout(\CONTROL.N_429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_8_LC_12_23_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_8_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_8_LC_12_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_8_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31346),
            .lcout(\CONTROL.dout_reto_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73253),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIDTCV_15_LC_12_23_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIDTCV_15_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIDTCV_15_LC_12_23_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIDTCV_15_LC_12_23_2  (
            .in0(N__33482),
            .in1(_gnd_net_),
            .in2(N__31424),
            .in3(N__29825),
            .lcout(progRomAddress_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_11_LC_12_23_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_11_LC_12_23_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_11_LC_12_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_11_LC_12_23_3  (
            .in0(N__29722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73253),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI5PM5H92_4_LC_12_23_4 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI5PM5H92_4_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI5PM5H92_4_LC_12_23_4 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \CONTROL.addrstackptr_RNI5PM5H92_4_LC_12_23_4  (
            .in0(N__29707),
            .in1(N__29681),
            .in2(N__60805),
            .in3(N__29674),
            .lcout(\CONTROL.addrstackptr_8_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_14_LC_12_23_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_14_LC_12_23_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_14_LC_12_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_14_LC_12_23_5  (
            .in0(N__29647),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73253),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI8INO_11_LC_12_23_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI8INO_11_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI8INO_11_LC_12_23_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI8INO_11_LC_12_23_6  (
            .in0(N__29627),
            .in1(N__29621),
            .in2(_gnd_net_),
            .in3(N__45120),
            .lcout(N_426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_11_LC_12_23_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_11_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_11_LC_12_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_11_LC_12_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30650),
            .lcout(\CONTROL.dout_reto_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73253),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m470_am_LC_12_24_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m470_am_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m470_am_LC_12_24_0 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m470_am_LC_12_24_0  (
            .in0(N__76624),
            .in1(N__75908),
            .in2(N__64265),
            .in3(N__64973),
            .lcout(\PROM.ROMDATA.m470_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_14_LC_12_24_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_14_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_14_LC_12_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_14_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30452),
            .lcout(\CONTROL.dout_reto_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73264),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_LC_12_24_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_LC_12_24_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_18_LC_12_24_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CONTROL.programCounter_ret_18_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__50837),
            .in2(_gnd_net_),
            .in3(N__50904),
            .lcout(\CONTROL.un1_programCounter9_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73264),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_10_LC_12_24_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_10_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_10_LC_12_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_1_10_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29846),
            .lcout(\CONTROL.programCounter_1_reto_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73264),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_35_rep1_LC_12_24_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_35_rep1_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_35_rep1_LC_12_24_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \CONTROL.programCounter_ret_35_rep1_LC_12_24_5  (
            .in0(N__50905),
            .in1(_gnd_net_),
            .in2(N__50843),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter11_reto_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73264),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI6GNO_10_LC_12_24_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI6GNO_10_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI6GNO_10_LC_12_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI6GNO_10_LC_12_24_6  (
            .in0(N__45119),
            .in1(N__34895),
            .in2(_gnd_net_),
            .in3(N__29801),
            .lcout(\CONTROL.N_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNID7J31_1_LC_12_24_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNID7J31_1_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNID7J31_1_LC_12_24_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.programCounter_ret_36_RNID7J31_1_LC_12_24_7  (
            .in0(N__73686),
            .in1(N__73574),
            .in2(_gnd_net_),
            .in3(N__73820),
            .lcout(\CONTROL.programCounter_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI45TU352_1_LC_12_25_0 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI45TU352_1_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI45TU352_1_LC_12_25_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \CONTROL.addrstackptr_RNI45TU352_1_LC_12_25_0  (
            .in0(N__31492),
            .in1(N__31444),
            .in2(N__31531),
            .in3(N__31541),
            .lcout(\CONTROL.addrstackptr_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI19JNL91_0_LC_12_25_2 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI19JNL91_0_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI19JNL91_0_LC_12_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CONTROL.addrstackptr_RNI19JNL91_0_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(N__57761),
            .in2(_gnd_net_),
            .in3(N__41981),
            .lcout(\CONTROL.addrstackptr_RNI19JNL91Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_9_LC_12_25_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_9_LC_12_25_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_9_LC_12_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_9_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40322),
            .lcout(\CONTROL.dout_reto_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73271),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_5_LC_13_7_0 .C_ON=1'b0;
    defparam \ALU.a_5_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \ALU.a_5_LC_13_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_5_LC_13_7_0  (
            .in0(N__57321),
            .in1(N__52637),
            .in2(_gnd_net_),
            .in3(N__39323),
            .lcout(\ALU.aZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73138),
            .ce(N__71215),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIET09P_0_12_LC_13_8_1 .C_ON=1'b0;
    defparam \ALU.c_RNIET09P_0_12_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIET09P_0_12_LC_13_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.c_RNIET09P_0_12_LC_13_8_1  (
            .in0(N__61195),
            .in1(N__61462),
            .in2(_gnd_net_),
            .in3(N__66598),
            .lcout(\ALU.N_614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICP0UG_5_LC_13_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNICP0UG_5_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICP0UG_5_LC_13_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNICP0UG_5_LC_13_8_2  (
            .in0(N__59583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68281),
            .lcout(\ALU.d_RNICP0UGZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBK47O_8_LC_13_8_3 .C_ON=1'b0;
    defparam \ALU.d_RNIBK47O_8_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBK47O_8_LC_13_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNIBK47O_8_LC_13_8_3  (
            .in0(N__61977),
            .in1(N__62872),
            .in2(_gnd_net_),
            .in3(N__66597),
            .lcout(\ALU.N_836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6CL331_4_LC_13_8_4 .C_ON=1'b0;
    defparam \ALU.d_RNI6CL331_4_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6CL331_4_LC_13_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI6CL331_4_LC_13_8_4  (
            .in0(N__59584),
            .in1(N__59894),
            .in2(N__68394),
            .in3(N__56401),
            .lcout(\ALU.d_RNI6CL331Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_173_c_RNO_0_LC_13_8_5 .C_ON=1'b0;
    defparam \ALU.mult_173_c_RNO_0_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_173_c_RNO_0_LC_13_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_173_c_RNO_0_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__59582),
            .in2(_gnd_net_),
            .in3(N__66596),
            .lcout(\ALU.mult_173_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILJMRC1_8_LC_13_8_6 .C_ON=1'b0;
    defparam \ALU.d_RNILJMRC1_8_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILJMRC1_8_LC_13_8_6 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \ALU.d_RNILJMRC1_8_LC_13_8_6  (
            .in0(N__66599),
            .in1(N__61978),
            .in2(N__62320),
            .in3(N__65954),
            .lcout(),
            .ltout(\ALU.d_RNILJMRC1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITH0GI3_8_LC_13_8_7 .C_ON=1'b0;
    defparam \ALU.d_RNITH0GI3_8_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITH0GI3_8_LC_13_8_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.d_RNITH0GI3_8_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__30326),
            .in2(N__29861),
            .in3(N__48232),
            .lcout(\ALU.N_642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_239_c_LC_13_9_0 .C_ON=1'b1;
    defparam \ALU.mult_239_c_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_239_c_LC_13_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_239_c_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__31721),
            .in2(N__31730),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\ALU.mult_7_c7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_239_c_RNI6DER62_LC_13_9_1 .C_ON=1'b1;
    defparam \ALU.mult_239_c_RNI6DER62_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_239_c_RNI6DER62_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_239_c_RNI6DER62_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__32864),
            .in2(N__29870),
            .in3(N__29858),
            .lcout(\ALU.mult_7_8 ),
            .ltout(),
            .carryin(\ALU.mult_7_c7 ),
            .carryout(\ALU.mult_7_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_245_c_RNISI9DS1_LC_13_9_2 .C_ON=1'b1;
    defparam \ALU.mult_245_c_RNISI9DS1_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_245_c_RNISI9DS1_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_245_c_RNISI9DS1_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__29855),
            .in2(N__29879),
            .in3(N__29849),
            .lcout(\ALU.mult_7_9 ),
            .ltout(),
            .carryin(\ALU.mult_7_c8 ),
            .carryout(\ALU.mult_7_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_251_c_RNIH3GMJ1_LC_13_9_3 .C_ON=1'b1;
    defparam \ALU.mult_251_c_RNIH3GMJ1_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_251_c_RNIH3GMJ1_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_251_c_RNIH3GMJ1_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__29993),
            .in2(N__29987),
            .in3(N__29969),
            .lcout(\ALU.mult_7_10 ),
            .ltout(),
            .carryin(\ALU.mult_7_c9 ),
            .carryout(\ALU.mult_7_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_257_c_RNIP79EM1_LC_13_9_4 .C_ON=1'b1;
    defparam \ALU.mult_257_c_RNIP79EM1_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_257_c_RNIP79EM1_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_257_c_RNIP79EM1_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__29966),
            .in2(N__29951),
            .in3(N__29933),
            .lcout(\ALU.mult_7_11 ),
            .ltout(),
            .carryin(\ALU.mult_7_c10 ),
            .carryout(\ALU.mult_7_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_263_c_RNIVGHJM1_LC_13_9_5 .C_ON=1'b1;
    defparam \ALU.mult_263_c_RNIVGHJM1_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_263_c_RNIVGHJM1_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_263_c_RNIVGHJM1_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__29930),
            .in2(N__30098),
            .in3(N__29915),
            .lcout(\ALU.mult_7_12 ),
            .ltout(),
            .carryin(\ALU.mult_7_c11 ),
            .carryout(\ALU.mult_7_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_269_c_RNIG3OFK1_LC_13_9_6 .C_ON=1'b1;
    defparam \ALU.mult_269_c_RNIG3OFK1_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_269_c_RNIG3OFK1_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_269_c_RNIG3OFK1_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__29912),
            .in2(N__37001),
            .in3(N__29900),
            .lcout(\ALU.mult_7_13 ),
            .ltout(),
            .carryin(\ALU.mult_7_c12 ),
            .carryout(\ALU.mult_7_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_275_c_RNIKBKSI1_LC_13_9_7 .C_ON=1'b1;
    defparam \ALU.mult_275_c_RNIKBKSI1_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_275_c_RNIKBKSI1_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_275_c_RNIKBKSI1_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__29897),
            .in2(N__46586),
            .in3(N__29885),
            .lcout(\ALU.mult_7_14 ),
            .ltout(),
            .carryin(\ALU.mult_7_c13 ),
            .carryout(\ALU.mult_7_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_7_c14_THRU_LUT4_0_LC_13_10_0 .C_ON=1'b0;
    defparam \ALU.mult_7_c14_THRU_LUT4_0_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_7_c14_THRU_LUT4_0_LC_13_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.mult_7_c14_THRU_LUT4_0_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29882),
            .lcout(\ALU.mult_7_c14_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFGNR61_4_LC_13_10_1 .C_ON=1'b0;
    defparam \ALU.d_RNIFGNR61_4_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFGNR61_4_LC_13_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIFGNR61_4_LC_13_10_1  (
            .in0(N__68745),
            .in1(N__59864),
            .in2(N__59599),
            .in3(N__68229),
            .lcout(\ALU.d_RNIFGNR61Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHNHG61_6_LC_13_10_2 .C_ON=1'b0;
    defparam \ALU.d_RNIHNHG61_6_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHNHG61_6_LC_13_10_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.d_RNIHNHG61_6_LC_13_10_2  (
            .in0(N__68230),
            .in1(N__62285),
            .in2(N__62557),
            .in3(N__68746),
            .lcout(\ALU.d_RNIHNHG61Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4LU7E1_6_LC_13_10_3 .C_ON=1'b0;
    defparam \ALU.d_RNI4LU7E1_6_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4LU7E1_6_LC_13_10_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNI4LU7E1_6_LC_13_10_3  (
            .in0(N__68744),
            .in1(N__62519),
            .in2(N__62306),
            .in3(N__66011),
            .lcout(\ALU.d_RNI4LU7E1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJAJOO_0_10_LC_13_10_4 .C_ON=1'b0;
    defparam \ALU.c_RNIJAJOO_0_10_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJAJOO_0_10_LC_13_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIJAJOO_0_10_LC_13_10_4  (
            .in0(N__62873),
            .in1(N__61666),
            .in2(_gnd_net_),
            .in3(N__66652),
            .lcout(\ALU.N_612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA6P2I_7_LC_13_10_6 .C_ON=1'b0;
    defparam \ALU.d_RNIA6P2I_7_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA6P2I_7_LC_13_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIA6P2I_7_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__62281),
            .in2(_gnd_net_),
            .in3(N__56267),
            .lcout(\ALU.d_RNIA6P2IZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIOGRG_1_LC_13_10_7 .C_ON=1'b0;
    defparam \ALU.d_RNIIOGRG_1_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIOGRG_1_LC_13_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIIOGRG_1_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__65520),
            .in2(_gnd_net_),
            .in3(N__68228),
            .lcout(\ALU.d_RNIIOGRGZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_5_c_LC_13_11_0 .C_ON=1'b1;
    defparam \ALU.mult_5_c_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_5_c_LC_13_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_5_c_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__32063),
            .in2(N__30503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\ALU.mult_1_c1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_5_c_RNIFR9072_LC_13_11_1 .C_ON=1'b1;
    defparam \ALU.mult_5_c_RNIFR9072_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_5_c_RNIFR9072_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_5_c_RNIFR9072_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__32402),
            .in2(N__32411),
            .in3(N__30086),
            .lcout(\ALU.mult_1_2 ),
            .ltout(),
            .carryin(\ALU.mult_1_c1 ),
            .carryout(\ALU.mult_1_c2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_11_c_RNIL35NS1_LC_13_11_2 .C_ON=1'b1;
    defparam \ALU.mult_11_c_RNIL35NS1_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_11_c_RNIL35NS1_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_11_c_RNIL35NS1_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__32099),
            .in2(N__30083),
            .in3(N__30074),
            .lcout(\ALU.mult_1_3 ),
            .ltout(),
            .carryin(\ALU.mult_1_c2 ),
            .carryout(\ALU.mult_1_c3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_17_c_RNIJ5JVJ1_LC_13_11_3 .C_ON=1'b1;
    defparam \ALU.mult_17_c_RNIJ5JVJ1_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_17_c_RNIJ5JVJ1_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_17_c_RNIJ5JVJ1_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__30071),
            .in2(N__30065),
            .in3(N__30050),
            .lcout(\ALU.mult_1_4 ),
            .ltout(),
            .carryin(\ALU.mult_1_c3 ),
            .carryout(\ALU.mult_1_c4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_23_c_RNIIO4OM1_LC_13_11_4 .C_ON=1'b1;
    defparam \ALU.mult_23_c_RNIIO4OM1_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_23_c_RNIIO4OM1_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_23_c_RNIIO4OM1_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__30047),
            .in2(N__30035),
            .in3(N__30023),
            .lcout(\ALU.mult_1_5 ),
            .ltout(),
            .carryin(\ALU.mult_1_c4 ),
            .carryout(\ALU.mult_1_c5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_29_c_RNI1JKSM1_LC_13_11_5 .C_ON=1'b1;
    defparam \ALU.mult_29_c_RNI1JKSM1_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_29_c_RNI1JKSM1_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_29_c_RNI1JKSM1_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__30020),
            .in2(N__30008),
            .in3(N__29996),
            .lcout(\ALU.mult_1_6 ),
            .ltout(),
            .carryin(\ALU.mult_1_c5 ),
            .carryout(\ALU.mult_1_c6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_35_c_RNI9KJPK1_LC_13_11_6 .C_ON=1'b1;
    defparam \ALU.mult_35_c_RNI9KJPK1_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_35_c_RNI9KJPK1_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_35_c_RNI9KJPK1_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__40163),
            .in2(N__30197),
            .in3(N__30185),
            .lcout(\ALU.mult_1_7 ),
            .ltout(),
            .carryin(\ALU.mult_1_c6 ),
            .carryout(\ALU.mult_1_c7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_41_c_RNIDSF6J1_LC_13_11_7 .C_ON=1'b1;
    defparam \ALU.mult_41_c_RNIDSF6J1_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_41_c_RNIDSF6J1_LC_13_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_41_c_RNIDSF6J1_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__30182),
            .in2(N__33977),
            .in3(N__30170),
            .lcout(\ALU.mult_1_8 ),
            .ltout(),
            .carryin(\ALU.mult_1_c7 ),
            .carryout(\ALU.mult_1_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_47_c_RNI86FRL1_LC_13_12_0 .C_ON=1'b1;
    defparam \ALU.mult_47_c_RNI86FRL1_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_47_c_RNI86FRL1_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_47_c_RNI86FRL1_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__30167),
            .in2(N__30254),
            .in3(N__30161),
            .lcout(\ALU.mult_1_9 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\ALU.mult_1_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_53_c_RNIV6GCO1_LC_13_12_1 .C_ON=1'b1;
    defparam \ALU.mult_53_c_RNIV6GCO1_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_53_c_RNIV6GCO1_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_53_c_RNIV6GCO1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__30260),
            .in2(N__30158),
            .in3(N__30146),
            .lcout(\ALU.mult_1_10 ),
            .ltout(),
            .carryin(\ALU.mult_1_c9 ),
            .carryout(\ALU.mult_1_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_59_c_RNILJ8EP1_LC_13_12_2 .C_ON=1'b1;
    defparam \ALU.mult_59_c_RNILJ8EP1_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_59_c_RNILJ8EP1_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_59_c_RNILJ8EP1_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__30143),
            .in2(N__30131),
            .in3(N__30122),
            .lcout(\ALU.mult_1_11 ),
            .ltout(),
            .carryin(\ALU.mult_1_c10 ),
            .carryout(\ALU.mult_1_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_65_c_RNI32HQN1_LC_13_12_3 .C_ON=1'b1;
    defparam \ALU.mult_65_c_RNI32HQN1_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_65_c_RNI32HQN1_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_65_c_RNI32HQN1_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__30236),
            .in2(N__30575),
            .in3(N__30119),
            .lcout(\ALU.mult_1_12 ),
            .ltout(),
            .carryin(\ALU.mult_1_c11 ),
            .carryout(\ALU.mult_1_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_71_c_RNIPD3ES1_LC_13_12_4 .C_ON=1'b1;
    defparam \ALU.mult_71_c_RNIPD3ES1_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_71_c_RNIPD3ES1_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_71_c_RNIPD3ES1_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__30116),
            .in2(N__37205),
            .in3(N__30104),
            .lcout(\ALU.mult_1_13 ),
            .ltout(),
            .carryin(\ALU.mult_1_c12 ),
            .carryout(\ALU.mult_1_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_77_c_RNIF6U9Q1_LC_13_12_5 .C_ON=1'b1;
    defparam \ALU.mult_77_c_RNIF6U9Q1_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_77_c_RNIF6U9Q1_LC_13_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_77_c_RNIF6U9Q1_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__30230),
            .in2(N__30221),
            .in3(N__30101),
            .lcout(\ALU.mult_1_14 ),
            .ltout(),
            .carryin(\ALU.mult_1_c13 ),
            .carryout(\ALU.mult_1_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_83_c_RNIKEU6B2_LC_13_12_6 .C_ON=1'b0;
    defparam \ALU.mult_83_c_RNIKEU6B2_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_83_c_RNIKEU6B2_LC_13_12_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_83_c_RNIKEU6B2_LC_13_12_6  (
            .in0(N__30212),
            .in1(N__30284),
            .in2(N__30278),
            .in3(N__30263),
            .lcout(\ALU.mult_83_c_RNIKEU6BZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI83GO51_0_LC_13_13_0 .C_ON=1'b0;
    defparam \ALU.d_RNI83GO51_0_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI83GO51_0_LC_13_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI83GO51_0_LC_13_13_0  (
            .in0(N__60542),
            .in1(N__65481),
            .in2(N__55686),
            .in3(N__55576),
            .lcout(\ALU.d_RNI83GO51Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPIBO31_0_LC_13_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIPIBO31_0_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPIBO31_0_LC_13_13_1 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.d_RNIPIBO31_0_LC_13_13_1  (
            .in0(N__65483),
            .in1(N__60541),
            .in2(N__55685),
            .in3(N__55821),
            .lcout(\ALU.d_RNIPIBO31Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIHC6L_3_LC_13_13_2 .C_ON=1'b0;
    defparam \ALU.d_RNIIHC6L_3_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIHC6L_3_LC_13_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIIHC6L_3_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__68658),
            .in2(_gnd_net_),
            .in3(N__60206),
            .lcout(\ALU.d_RNIIHC6LZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITH0K51_0_LC_13_13_3 .C_ON=1'b0;
    defparam \ALU.d_RNITH0K51_0_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITH0K51_0_LC_13_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNITH0K51_0_LC_13_13_3  (
            .in0(N__57039),
            .in1(N__56904),
            .in2(N__65546),
            .in3(N__60543),
            .lcout(\ALU.d_RNITH0K51Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0H41K_1_LC_13_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNI0H41K_1_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0H41K_1_LC_13_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI0H41K_1_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__56805),
            .in2(_gnd_net_),
            .in3(N__65479),
            .lcout(\ALU.d_RNI0H41KZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIETL861_0_LC_13_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNIETL861_0_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIETL861_0_LC_13_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIETL861_0_LC_13_13_5  (
            .in0(N__65482),
            .in1(N__56737),
            .in2(N__56823),
            .in3(N__60544),
            .lcout(\ALU.d_RNIETL861Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8FM541_0_LC_13_13_6 .C_ON=1'b0;
    defparam \ALU.d_RNI8FM541_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8FM541_0_LC_13_13_6 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.d_RNI8FM541_0_LC_13_13_6  (
            .in0(N__60545),
            .in1(N__74609),
            .in2(N__56748),
            .in3(N__65480),
            .lcout(\ALU.d_RNI8FM541Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGIF4D1_2_LC_13_13_7 .C_ON=1'b0;
    defparam \ALU.d_RNIGIF4D1_2_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGIF4D1_2_LC_13_13_7 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.d_RNIGIF4D1_2_LC_13_13_7  (
            .in0(N__60207),
            .in1(N__66241),
            .in2(N__68733),
            .in3(N__66012),
            .lcout(\ALU.d_RNIGIF4D1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINLH9L_2_LC_13_14_0 .C_ON=1'b0;
    defparam \ALU.d_RNINLH9L_2_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINLH9L_2_LC_13_14_0 .LUT_INIT=16'b0111011001101000;
    LogicCell40 \ALU.d_RNINLH9L_2_LC_13_14_0  (
            .in0(N__68720),
            .in1(N__74834),
            .in2(N__63290),
            .in3(N__66252),
            .lcout(\ALU.log_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN178L_2_LC_13_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNIN178L_2_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN178L_2_LC_13_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.d_RNIN178L_2_LC_13_14_1  (
            .in0(N__66253),
            .in1(N__63248),
            .in2(_gnd_net_),
            .in3(N__68719),
            .lcout(\ALU.d_RNIN178LZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIBPDT_11_LC_13_14_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIBPDT_11_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIBPDT_11_LC_13_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIBPDT_11_LC_13_14_3  (
            .in0(N__30406),
            .in1(N__30377),
            .in2(_gnd_net_),
            .in3(N__64664),
            .lcout(progRomAddress_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILJMRC1_0_8_LC_13_14_4 .C_ON=1'b0;
    defparam \ALU.d_RNILJMRC1_0_8_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILJMRC1_0_8_LC_13_14_4 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \ALU.d_RNILJMRC1_0_8_LC_13_14_4  (
            .in0(N__62261),
            .in1(N__66441),
            .in2(N__61975),
            .in3(N__65930),
            .lcout(\ALU.d_RNILJMRC1_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI58QFI_5_LC_13_14_7 .C_ON=1'b0;
    defparam \ALU.d_RNI58QFI_5_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI58QFI_5_LC_13_14_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.d_RNI58QFI_5_LC_13_14_7  (
            .in0(N__59625),
            .in1(N__63249),
            .in2(_gnd_net_),
            .in3(N__33993),
            .lcout(\ALU.d_RNI58QFIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.combOperand2_1_0_LC_13_15_0 .C_ON=1'b0;
    defparam \ALU.combOperand2_1_0_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.combOperand2_1_0_LC_13_15_0 .LUT_INIT=16'b0001000100011011;
    LogicCell40 \ALU.combOperand2_1_0_LC_13_15_0  (
            .in0(N__53145),
            .in1(N__36918),
            .in2(N__32846),
            .in3(N__38847),
            .lcout(),
            .ltout(\ALU.combOperand2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFFCPG_0_LC_13_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIFFCPG_0_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFFCPG_0_LC_13_15_1 .LUT_INIT=16'b0001111100001110;
    LogicCell40 \ALU.d_RNIFFCPG_0_LC_13_15_1  (
            .in0(N__71395),
            .in1(N__53146),
            .in2(N__30314),
            .in3(N__37870),
            .lcout(\ALU.status_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI6KJL_0_LC_13_15_2 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI6KJL_0_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI6KJL_0_LC_13_15_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI6KJL_0_LC_13_15_2  (
            .in0(N__32318),
            .in1(N__30473),
            .in2(_gnd_net_),
            .in3(N__30490),
            .lcout(),
            .ltout(DROM_ROMDATA_dintern_0ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIAR0U1_2_LC_13_15_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIAR0U1_2_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIAR0U1_2_LC_13_15_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \CONTROL.busState_1_RNIAR0U1_2_LC_13_15_3  (
            .in0(N__49562),
            .in1(N__30311),
            .in2(N__30299),
            .in3(N__30296),
            .lcout(busState_1_RNIAR0U1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.combOperand2_a0_0_6_LC_13_15_4 .C_ON=1'b0;
    defparam \ALU.combOperand2_a0_0_6_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.combOperand2_a0_0_6_LC_13_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.combOperand2_a0_0_6_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__71394),
            .in2(_gnd_net_),
            .in3(N__49793),
            .lcout(\ALU.combOperand2_a0_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIR8PGB_0_LC_13_15_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIR8PGB_0_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIR8PGB_0_LC_13_15_5 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \CONTROL.busState_1_RNIR8PGB_0_LC_13_15_5  (
            .in0(N__38848),
            .in1(N__49797),
            .in2(N__36925),
            .in3(N__32845),
            .lcout(bus_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_5_c_RNO_0_LC_13_15_6 .C_ON=1'b0;
    defparam \ALU.mult_5_c_RNO_0_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_5_c_RNO_0_LC_13_15_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_5_c_RNO_0_LC_13_15_6  (
            .in0(N__65351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66375),
            .lcout(\ALU.mult_5_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_0_LC_13_15_7 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_0_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_0_LC_13_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_0_LC_13_15_7  (
            .in0(N__30491),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C_net ),
            .ce(N__32319),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_14_LC_13_16_0 .C_ON=1'b0;
    defparam \CONTROL.dout_14_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_14_LC_13_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \CONTROL.dout_14_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__30994),
            .in2(_gnd_net_),
            .in3(N__40915),
            .lcout(\CONTROL.ctrlOut_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_14C_net ),
            .ce(N__44453),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI6ADU_14_LC_13_16_1 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI6ADU_14_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI6ADU_14_LC_13_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNI6ADU_14_LC_13_16_1  (
            .in0(N__30467),
            .in1(N__30445),
            .in2(_gnd_net_),
            .in3(N__50147),
            .lcout(),
            .ltout(\CONTROL.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIHTF52_2_LC_13_16_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIHTF52_2_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIHTF52_2_LC_13_16_2 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \CONTROL.busState_1_RNIHTF52_2_LC_13_16_2  (
            .in0(N__50148),
            .in1(N__30434),
            .in2(N__30413),
            .in3(N__49572),
            .lcout(N_191),
            .ltout(N_191_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNISBR29_0_LC_13_16_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNISBR29_0_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNISBR29_0_LC_13_16_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \CONTROL.busState_1_RNISBR29_0_LC_13_16_3  (
            .in0(N__49573),
            .in1(N__47072),
            .in2(N__30410),
            .in3(N__49815),
            .lcout(bus_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_30dflt_LC_13_16_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_30dflt_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_30dflt_LC_13_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PROM.ROMDATA.dintern_30dflt_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(N__30993),
            .in2(_gnd_net_),
            .in3(N__40914),
            .lcout(controlWord_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIRA1I6_2_LC_13_16_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIRA1I6_2_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIRA1I6_2_LC_13_16_5 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \CONTROL.busState_1_RNIRA1I6_2_LC_13_16_5  (
            .in0(N__49574),
            .in1(N__34099),
            .in2(N__50200),
            .in3(N__65408),
            .lcout(),
            .ltout(\CONTROL.busState_1_RNIRA1I6Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI2BDF8_0_LC_13_16_6 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI2BDF8_0_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI2BDF8_0_LC_13_16_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \CONTROL.busState_1_RNI2BDF8_0_LC_13_16_6  (
            .in0(N__49816),
            .in1(_gnd_net_),
            .in2(N__30578),
            .in3(N__33032),
            .lcout(bus_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8VHNH_1_LC_13_16_7 .C_ON=1'b0;
    defparam \ALU.d_RNI8VHNH_1_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8VHNH_1_LC_13_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNI8VHNH_1_LC_13_16_7  (
            .in0(N__56987),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65407),
            .lcout(\ALU.d_RNI8VHNHZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI13B91_12_LC_13_17_0 .C_ON=1'b0;
    defparam \ALU.a_RNI13B91_12_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI13B91_12_LC_13_17_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.a_RNI13B91_12_LC_13_17_0  (
            .in0(N__48265),
            .in1(N__43917),
            .in2(N__51422),
            .in3(N__32821),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI49JM1_12_LC_13_17_1 .C_ON=1'b0;
    defparam \ALU.c_RNI49JM1_12_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI49JM1_12_LC_13_17_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNI49JM1_12_LC_13_17_1  (
            .in0(N__52410),
            .in1(N__67549),
            .in2(N__30560),
            .in3(N__54294),
            .lcout(\ALU.N_1097 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI4EQI1_12_LC_13_17_2 .C_ON=1'b0;
    defparam \ALU.b_RNI4EQI1_12_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI4EQI1_12_LC_13_17_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI4EQI1_12_LC_13_17_2  (
            .in0(N__39817),
            .in1(N__34542),
            .in2(N__57686),
            .in3(N__43916),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9SE82_12_LC_13_17_3 .C_ON=1'b0;
    defparam \ALU.d_RNI9SE82_12_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9SE82_12_LC_13_17_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNI9SE82_12_LC_13_17_3  (
            .in0(N__57934),
            .in1(N__65089),
            .in2(N__30557),
            .in3(N__54295),
            .lcout(),
            .ltout(\ALU.N_1145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIG9G84_12_LC_13_17_4 .C_ON=1'b0;
    defparam \ALU.c_RNIG9G84_12_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIG9G84_12_LC_13_17_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.c_RNIG9G84_12_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__30554),
            .in2(N__30548),
            .in3(N__54130),
            .lcout(aluOut_12),
            .ltout(aluOut_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI6CUR7_0_LC_13_17_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI6CUR7_0_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI6CUR7_0_LC_13_17_5 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \CONTROL.busState_1_RNI6CUR7_0_LC_13_17_5  (
            .in0(N__30587),
            .in1(N__34483),
            .in2(N__30545),
            .in3(N__49810),
            .lcout(\CONTROL.bus_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI04DU_11_LC_13_18_0 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI04DU_11_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI04DU_11_LC_13_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.dout_RNI04DU_11_LC_13_18_0  (
            .in0(N__50106),
            .in1(N__30527),
            .in2(_gnd_net_),
            .in3(N__30643),
            .lcout(),
            .ltout(\CONTROL.N_172_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI8VQQ1_2_LC_13_18_1 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI8VQQ1_2_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI8VQQ1_2_LC_13_18_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \CONTROL.busState_1_RNI8VQQ1_2_LC_13_18_1  (
            .in0(N__49494),
            .in1(N__30701),
            .in2(N__30680),
            .in3(N__50107),
            .lcout(N_188),
            .ltout(N_188_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIQBOE8_0_LC_13_18_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIQBOE8_0_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIQBOE8_0_LC_13_18_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \CONTROL.busState_1_RNIQBOE8_0_LC_13_18_2  (
            .in0(N__30668),
            .in1(N__49811),
            .in2(N__30653),
            .in3(N__49495),
            .lcout(bus_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_11_LC_13_18_3 .C_ON=1'b0;
    defparam \CONTROL.dout_11_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_11_LC_13_18_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \CONTROL.dout_11_LC_13_18_3  (
            .in0(N__72129),
            .in1(N__47475),
            .in2(N__72768),
            .in3(N__36950),
            .lcout(\CONTROL.ctrlOut_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_11C_net ),
            .ce(N__44415),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_27dflt_LC_13_18_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_27dflt_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_27dflt_LC_13_18_4 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_27dflt_LC_13_18_4  (
            .in0(N__36949),
            .in1(N__72713),
            .in2(N__47488),
            .in3(N__72128),
            .lcout(controlWord_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_12_LC_13_18_5 .C_ON=1'b0;
    defparam \CONTROL.dout_12_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_12_LC_13_18_5 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \CONTROL.dout_12_LC_13_18_5  (
            .in0(N__72130),
            .in1(N__65150),
            .in2(N__72769),
            .in3(N__47476),
            .lcout(\CONTROL.ctrlOut_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_11C_net ),
            .ce(N__44415),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI26DU_12_LC_13_18_6 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI26DU_12_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI26DU_12_LC_13_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.dout_RNI26DU_12_LC_13_18_6  (
            .in0(N__50104),
            .in1(N__30632),
            .in2(_gnd_net_),
            .in3(N__38764),
            .lcout(),
            .ltout(\CONTROL.N_173_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIB9N32_2_LC_13_18_7 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIB9N32_2_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIB9N32_2_LC_13_18_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \CONTROL.busState_1_RNIB9N32_2_LC_13_18_7  (
            .in0(N__49493),
            .in1(N__30611),
            .in2(N__30590),
            .in3(N__50105),
            .lcout(\CONTROL.N_189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState14_1_i_o2_LC_13_19_0 .C_ON=1'b0;
    defparam \CONTROL.un1_busState14_1_i_o2_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState14_1_i_o2_LC_13_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \CONTROL.un1_busState14_1_i_o2_LC_13_19_0  (
            .in0(N__41245),
            .in1(N__41408),
            .in2(N__36883),
            .in3(N__54677),
            .lcout(\CONTROL.un1_busState14_1_i_o2_0 ),
            .ltout(\CONTROL.un1_busState14_1_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState12_2_i_a2_d_0_tz_LC_13_19_1 .C_ON=1'b0;
    defparam \CONTROL.un1_busState12_2_i_a2_d_0_tz_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState12_2_i_a2_d_0_tz_LC_13_19_1 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \CONTROL.un1_busState12_2_i_a2_d_0_tz_LC_13_19_1  (
            .in0(N__30880),
            .in1(N__36433),
            .in2(N__30581),
            .in3(N__41246),
            .lcout(),
            .ltout(\CONTROL.un1_busState12_2_i_a2_0_1_tz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState12_2_i_a2_0_i_LC_13_19_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState12_2_i_a2_0_i_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState12_2_i_a2_0_i_LC_13_19_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \CONTROL.un1_busState12_2_i_a2_0_i_LC_13_19_2  (
            .in0(N__36821),
            .in1(N__35171),
            .in2(N__30821),
            .in3(N__30791),
            .lcout(\CONTROL.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_LC_13_19_3 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_LC_13_19_3 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \CONTROL.aluReadBus_1_sqmuxa_0_a2_LC_13_19_3  (
            .in0(N__30881),
            .in1(N__38717),
            .in2(N__36448),
            .in3(N__41248),
            .lcout(\CONTROL.aluReadBus_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState119_i_i_a2_LC_13_19_4 .C_ON=1'b0;
    defparam \CONTROL.busState119_i_i_a2_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState119_i_i_a2_LC_13_19_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \CONTROL.busState119_i_i_a2_LC_13_19_4  (
            .in0(N__36684),
            .in1(N__54678),
            .in2(N__41259),
            .in3(N__44708),
            .lcout(\CONTROL.N_244 ),
            .ltout(\CONTROL.N_244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_LC_13_19_5 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluReadBus_LC_13_19_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \CONTROL.aluReadBus_LC_13_19_5  (
            .in0(N__36578),
            .in1(N__30809),
            .in2(N__30818),
            .in3(N__71314),
            .lcout(aluReadBus),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluReadBusC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState98_1_1_0_LC_13_19_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState98_1_1_0_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState98_1_1_0_LC_13_19_6 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \CONTROL.un1_busState98_1_1_0_LC_13_19_6  (
            .in0(N__41249),
            .in1(N__36443),
            .in2(_gnd_net_),
            .in3(N__33473),
            .lcout(\CONTROL.un1_busState98_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState14_1_i_a2_1_i_1_LC_13_19_7 .C_ON=1'b0;
    defparam \CONTROL.un1_busState14_1_i_a2_1_i_1_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState14_1_i_a2_1_i_1_LC_13_19_7 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \CONTROL.un1_busState14_1_i_a2_1_i_1_LC_13_19_7  (
            .in0(N__30879),
            .in1(N__30815),
            .in2(N__36447),
            .in3(N__41247),
            .lcout(\CONTROL.un1_busState14_1_i_a2_1_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_RNO_0_LC_13_20_0 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_RNO_0_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluReadBus_RNO_0_LC_13_20_0 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \CONTROL.aluReadBus_RNO_0_LC_13_20_0  (
            .in0(N__41429),
            .in1(N__30707),
            .in2(N__36609),
            .in3(N__44898),
            .lcout(\CONTROL.aluReadBus_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState14_1_i_a2_1_i_LC_13_20_1 .C_ON=1'b0;
    defparam \CONTROL.un1_busState14_1_i_a2_1_i_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState14_1_i_a2_1_i_LC_13_20_1 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \CONTROL.un1_busState14_1_i_a2_1_i_LC_13_20_1  (
            .in0(N__38323),
            .in1(N__30800),
            .in2(N__38657),
            .in3(N__30792),
            .lcout(\CONTROL.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState101_3_0_m2_LC_13_20_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState101_3_0_m2_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState101_3_0_m2_LC_13_20_2 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \CONTROL.un1_busState101_3_0_m2_LC_13_20_2  (
            .in0(N__41428),
            .in1(N__55474),
            .in2(N__36884),
            .in3(N__54670),
            .lcout(\CONTROL.N_89 ),
            .ltout(\CONTROL.N_89_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState101_3_0_0_LC_13_20_3 .C_ON=1'b0;
    defparam \CONTROL.un1_busState101_3_0_0_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState101_3_0_0_LC_13_20_3 .LUT_INIT=16'b0000001100001111;
    LogicCell40 \CONTROL.un1_busState101_3_0_0_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__41594),
            .in2(N__30887),
            .in3(N__36688),
            .lcout(\CONTROL.un1_busState101_3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState103_0_o2_0_LC_13_20_4 .C_ON=1'b0;
    defparam \CONTROL.un1_busState103_0_o2_0_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState103_0_o2_0_LC_13_20_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \CONTROL.un1_busState103_0_o2_0_LC_13_20_4  (
            .in0(N__44705),
            .in1(N__54668),
            .in2(N__41435),
            .in3(N__44897),
            .lcout(\CONTROL.N_101_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState97_1_0_o2_LC_13_20_5 .C_ON=1'b0;
    defparam \CONTROL.un1_busState97_1_0_o2_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState97_1_0_o2_LC_13_20_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \CONTROL.un1_busState97_1_0_o2_LC_13_20_5  (
            .in0(N__54669),
            .in1(N__55473),
            .in2(_gnd_net_),
            .in3(N__44707),
            .lcout(\CONTROL.N_87_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_0_0_LC_13_20_6 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_0_0_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_0_0_LC_13_20_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \CONTROL.aluReadBus_1_sqmuxa_0_a2_0_0_LC_13_20_6  (
            .in0(N__55472),
            .in1(N__42244),
            .in2(_gnd_net_),
            .in3(N__72181),
            .lcout(),
            .ltout(\CONTROL.aluReadBus_1_sqmuxa_0_a2_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_LC_13_20_7 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_LC_13_20_7 .LUT_INIT=16'b0001001100100111;
    LogicCell40 \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_LC_13_20_7  (
            .in0(N__44896),
            .in1(N__36506),
            .in2(N__30884),
            .in3(N__44706),
            .lcout(\CONTROL.aluReadBus_1_sqmuxa_0_o2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_10_LC_13_21_0 .C_ON=1'b0;
    defparam \CONTROL.dout_10_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_10_LC_13_21_0 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \CONTROL.dout_10_LC_13_21_0  (
            .in0(N__72191),
            .in1(N__73945),
            .in2(N__72790),
            .in3(N__62609),
            .lcout(\CONTROL.ctrlOut_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_10C_net ),
            .ce(N__44445),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNIU1DU_10_LC_13_21_1 .C_ON=1'b0;
    defparam \CONTROL.dout_RNIU1DU_10_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNIU1DU_10_LC_13_21_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNIU1DU_10_LC_13_21_1  (
            .in0(N__30869),
            .in1(N__34906),
            .in2(_gnd_net_),
            .in3(N__50019),
            .lcout(),
            .ltout(\CONTROL.N_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI5LU12_2_LC_13_21_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI5LU12_2_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI5LU12_2_LC_13_21_2 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \CONTROL.busState_1_RNI5LU12_2_LC_13_21_2  (
            .in0(N__50021),
            .in1(N__30854),
            .in2(N__30836),
            .in3(N__49391),
            .lcout(\CONTROL.N_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_26dflt_LC_13_21_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_26dflt_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_26dflt_LC_13_21_3 .LUT_INIT=16'b1101000100000000;
    LogicCell40 \PROM.ROMDATA.dintern_26dflt_LC_13_21_3  (
            .in0(N__62608),
            .in1(N__72777),
            .in2(N__73946),
            .in3(N__72189),
            .lcout(controlWord_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_0_LC_13_21_4 .C_ON=1'b0;
    defparam \CONTROL.dout_0_LC_13_21_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_0_LC_13_21_4 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \CONTROL.dout_0_LC_13_21_4  (
            .in0(N__72190),
            .in1(N__64057),
            .in2(N__72789),
            .in3(N__74330),
            .lcout(\CONTROL.ctrlOut_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_10C_net ),
            .ce(N__44445),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNISBOJ_0_LC_13_21_5 .C_ON=1'b0;
    defparam \CONTROL.dout_RNISBOJ_0_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNISBOJ_0_LC_13_21_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNISBOJ_0_LC_13_21_5  (
            .in0(N__31028),
            .in1(N__45076),
            .in2(_gnd_net_),
            .in3(N__50020),
            .lcout(),
            .ltout(\CONTROL.N_161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNII0IO1_2_LC_13_21_6 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNII0IO1_2_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNII0IO1_2_LC_13_21_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \CONTROL.busState_1_RNII0IO1_2_LC_13_21_6  (
            .in0(N__50022),
            .in1(N__31010),
            .in2(N__30998),
            .in3(N__49392),
            .lcout(N_177),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_16dflt_LC_13_21_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_16dflt_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_16dflt_LC_13_21_7 .LUT_INIT=16'b1101000100000000;
    LogicCell40 \PROM.ROMDATA.dintern_16dflt_LC_13_21_7  (
            .in0(N__74329),
            .in1(N__72776),
            .in2(N__64058),
            .in3(N__72188),
            .lcout(controlWord_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.combOperand2_d_bm_15_LC_13_22_0 .C_ON=1'b0;
    defparam \ALU.combOperand2_d_bm_15_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \ALU.combOperand2_d_bm_15_LC_13_22_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \ALU.combOperand2_d_bm_15_LC_13_22_0  (
            .in0(N__50005),
            .in1(N__30941),
            .in2(N__30935),
            .in3(N__49545),
            .lcout(\ALU.combOperand2_d_bmZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_15_LC_13_22_1 .C_ON=1'b0;
    defparam \CONTROL.dout_15_LC_13_22_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_15_LC_13_22_1 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \CONTROL.dout_15_LC_13_22_1  (
            .in0(N__72193),
            .in1(N__30992),
            .in2(N__72791),
            .in3(N__47490),
            .lcout(\CONTROL.ctrlOut_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_15C_net ),
            .ce(N__44435),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31dflt_LC_13_22_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31dflt_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31dflt_LC_13_22_2 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31dflt_LC_13_22_2  (
            .in0(N__47489),
            .in1(N__72784),
            .in2(N__30995),
            .in3(N__72192),
            .lcout(controlWord_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI8CDU_15_LC_13_22_3 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI8CDU_15_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI8CDU_15_LC_13_22_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNI8CDU_15_LC_13_22_3  (
            .in0(N__30962),
            .in1(N__33433),
            .in2(_gnd_net_),
            .in3(N__50004),
            .lcout(N_176),
            .ltout(N_176_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIK7CU1_2_LC_13_22_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIK7CU1_2_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIK7CU1_2_LC_13_22_4 .LUT_INIT=16'b0000111101110111;
    LogicCell40 \CONTROL.busState_1_RNIK7CU1_2_LC_13_22_4  (
            .in0(N__50006),
            .in1(N__30934),
            .in2(N__30890),
            .in3(N__49546),
            .lcout(\CONTROL.bus_7_ns_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_8_LC_13_22_6 .C_ON=1'b0;
    defparam \CONTROL.dout_8_LC_13_22_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_8_LC_13_22_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \CONTROL.dout_8_LC_13_22_6  (
            .in0(N__31376),
            .in1(N__72785),
            .in2(N__47495),
            .in3(N__72194),
            .lcout(\CONTROL.ctrlOut_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_15C_net ),
            .ce(N__44435),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNICSOJ_8_LC_13_22_7 .C_ON=1'b0;
    defparam \CONTROL.dout_RNICSOJ_8_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNICSOJ_8_LC_13_22_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNICSOJ_8_LC_13_22_7  (
            .in0(N__31367),
            .in1(N__31345),
            .in2(_gnd_net_),
            .in3(N__50003),
            .lcout(\CONTROL.N_169 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_0_LC_13_23_0 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_0_LC_13_23_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_0_LC_13_23_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.ramAddReg_0_LC_13_23_0  (
            .in0(N__33313),
            .in1(N__70754),
            .in2(N__49136),
            .in3(N__70525),
            .lcout(A0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_0C_net ),
            .ce(N__70318),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_1_LC_13_23_1 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_1_LC_13_23_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_1_LC_13_23_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \CONTROL.ramAddReg_1_LC_13_23_1  (
            .in0(N__70523),
            .in1(N__33247),
            .in2(N__49181),
            .in3(N__70759),
            .lcout(A1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_0C_net ),
            .ce(N__70318),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_10_LC_13_23_2 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_10_LC_13_23_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_10_LC_13_23_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.ramAddReg_10_LC_13_23_2  (
            .in0(N__31275),
            .in1(N__70755),
            .in2(N__36008),
            .in3(N__70526),
            .lcout(A10_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_0C_net ),
            .ce(N__70318),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_11_LC_13_23_3 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_11_LC_13_23_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_11_LC_13_23_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \CONTROL.ramAddReg_11_LC_13_23_3  (
            .in0(N__70522),
            .in1(N__35967),
            .in2(N__31238),
            .in3(N__70758),
            .lcout(A11_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_0C_net ),
            .ce(N__70318),
            .sr(_gnd_net_));
    defparam \RAM.un1_WR_105_0_9_LC_13_23_4 .C_ON=1'b0;
    defparam \RAM.un1_WR_105_0_9_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \RAM.un1_WR_105_0_9_LC_13_23_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RAM.un1_WR_105_0_9_LC_13_23_4  (
            .in0(N__31039),
            .in1(N__31192),
            .in2(N__31168),
            .in3(N__31096),
            .lcout(\RAM.un1_WR_105_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_9_LC_13_23_6 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_9_LC_13_23_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_9_LC_13_23_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \CONTROL.ramAddReg_9_LC_13_23_6  (
            .in0(N__48998),
            .in1(N__70756),
            .in2(N__31136),
            .in3(N__70527),
            .lcout(A9_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_0C_net ),
            .ce(N__70318),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_8_LC_13_23_7 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_8_LC_13_23_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_8_LC_13_23_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \CONTROL.ramAddReg_8_LC_13_23_7  (
            .in0(N__70524),
            .in1(N__49052),
            .in2(N__31085),
            .in3(N__70760),
            .lcout(A8_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_0C_net ),
            .ce(N__70318),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI0N94M91_1_LC_13_24_0 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI0N94M91_1_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI0N94M91_1_LC_13_24_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \CONTROL.addrstackptr_RNI0N94M91_1_LC_13_24_0  (
            .in0(N__38415),
            .in1(N__57809),
            .in2(_gnd_net_),
            .in3(N__41960),
            .lcout(\CONTROL.g1_0 ),
            .ltout(\CONTROL.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_1_LC_13_24_1 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_1_LC_13_24_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_1_LC_13_24_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \CONTROL.addrstackptr_1_LC_13_24_1  (
            .in0(N__31445),
            .in1(N__31535),
            .in2(N__31499),
            .in3(N__31493),
            .lcout(\CONTROL.addrstackptrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.addrstackptr_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_1_i_a6_4_LC_13_24_2 .C_ON=1'b0;
    defparam \CONTROL.g0_1_i_a6_4_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_1_i_a6_4_LC_13_24_2 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \CONTROL.g0_1_i_a6_4_LC_13_24_2  (
            .in0(N__42264),
            .in1(N__36281),
            .in2(N__48488),
            .in3(N__38216),
            .lcout(),
            .ltout(\CONTROL.g0_1_i_a6Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_1_i_a6_LC_13_24_3 .C_ON=1'b0;
    defparam \CONTROL.g0_1_i_a6_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_1_i_a6_LC_13_24_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \CONTROL.g0_1_i_a6_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__40709),
            .in2(N__31496),
            .in3(N__40691),
            .lcout(\CONTROL.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNITQCP_1_LC_13_24_4 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNITQCP_1_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNITQCP_1_LC_13_24_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \CONTROL.addrstackptr_RNITQCP_1_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__38411),
            .in2(_gnd_net_),
            .in3(N__57808),
            .lcout(\CONTROL.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState_1_sqmuxa_i_a2_2_LC_13_24_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_a2_2_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_a2_2_LC_13_24_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \CONTROL.un1_busState_1_sqmuxa_i_a2_2_LC_13_24_6  (
            .in0(N__42263),
            .in1(N__55399),
            .in2(N__72306),
            .in3(N__71854),
            .lcout(\CONTROL.N_366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI94D27G_7_LC_13_25_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI94D27G_7_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI94D27G_7_LC_13_25_5 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI94D27G_7_LC_13_25_5  (
            .in0(N__72271),
            .in1(N__55475),
            .in2(N__36650),
            .in3(N__41496),
            .lcout(\CONTROL.g0_1_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_15_LC_13_25_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_15_LC_13_25_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_15_LC_13_25_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_36_15_LC_13_25_7  (
            .in0(N__31433),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.addrstack_reto_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73265),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_14_LC_13_26_0 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_14_LC_13_26_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_14_LC_13_26_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.ramAddReg_14_LC_13_26_0  (
            .in0(N__31404),
            .in1(N__70757),
            .in2(N__57593),
            .in3(N__70521),
            .lcout(A14_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_14C_net ),
            .ce(N__70328),
            .sr(_gnd_net_));
    defparam \ALU.mult_173_c_LC_14_8_0 .C_ON=1'b1;
    defparam \ALU.mult_173_c_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_173_c_LC_14_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_173_c_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__33713),
            .in2(N__31688),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\ALU.mult_5_c5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_173_c_RNIFBQH72_LC_14_8_1 .C_ON=1'b1;
    defparam \ALU.mult_173_c_RNIFBQH72_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_173_c_RNIFBQH72_LC_14_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_173_c_RNIFBQH72_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__33947),
            .in2(N__32093),
            .in3(N__31679),
            .lcout(\ALU.mult_5_6 ),
            .ltout(),
            .carryin(\ALU.mult_5_c5 ),
            .carryout(\ALU.mult_5_c6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_179_c_RNIE2T2T1_LC_14_8_2 .C_ON=1'b1;
    defparam \ALU.mult_179_c_RNIE2T2T1_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_179_c_RNIE2T2T1_LC_14_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_179_c_RNIE2T2T1_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__31676),
            .in2(N__33959),
            .in3(N__31667),
            .lcout(\ALU.mult_5_7 ),
            .ltout(),
            .carryin(\ALU.mult_5_c6 ),
            .carryout(\ALU.mult_5_c7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_185_c_RNI3J3CK1_LC_14_8_3 .C_ON=1'b1;
    defparam \ALU.mult_185_c_RNI3J3CK1_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_185_c_RNI3J3CK1_LC_14_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_185_c_RNI3J3CK1_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__31664),
            .in2(N__31658),
            .in3(N__31649),
            .lcout(\ALU.mult_5_8 ),
            .ltout(),
            .carryin(\ALU.mult_5_c7 ),
            .carryout(\ALU.mult_5_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_191_c_RNI26L4N1_LC_14_8_4 .C_ON=1'b1;
    defparam \ALU.mult_191_c_RNI26L4N1_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_191_c_RNI26L4N1_LC_14_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_191_c_RNI26L4N1_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__31646),
            .in2(N__33773),
            .in3(N__31634),
            .lcout(\ALU.mult_5_9 ),
            .ltout(),
            .carryin(\ALU.mult_5_c8 ),
            .carryout(\ALU.mult_5_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_197_c_RNIH059N1_LC_14_8_5 .C_ON=1'b1;
    defparam \ALU.mult_197_c_RNIH059N1_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_197_c_RNIH059N1_LC_14_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_197_c_RNIH059N1_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__31631),
            .in2(N__31619),
            .in3(N__31607),
            .lcout(\ALU.mult_5_10 ),
            .ltout(),
            .carryin(\ALU.mult_5_c9 ),
            .carryout(\ALU.mult_5_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_203_c_RNIG7BVK1_LC_14_8_6 .C_ON=1'b1;
    defparam \ALU.mult_203_c_RNIG7BVK1_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_203_c_RNIG7BVK1_LC_14_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_203_c_RNIG7BVK1_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__31604),
            .in2(N__31589),
            .in3(N__31574),
            .lcout(\ALU.mult_5_11 ),
            .ltout(),
            .carryin(\ALU.mult_5_c10 ),
            .carryout(\ALU.mult_5_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_209_c_RNIT0FBJ1_LC_14_8_7 .C_ON=1'b1;
    defparam \ALU.mult_209_c_RNIT0FBJ1_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_209_c_RNIT0FBJ1_LC_14_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_209_c_RNIT0FBJ1_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__31571),
            .in2(N__31559),
            .in3(N__31544),
            .lcout(\ALU.mult_5_12 ),
            .ltout(),
            .carryin(\ALU.mult_5_c11 ),
            .carryout(\ALU.mult_5_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_215_c_RNIFP61M1_LC_14_9_0 .C_ON=1'b1;
    defparam \ALU.mult_215_c_RNIFP61M1_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_215_c_RNIFP61M1_LC_14_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_215_c_RNIFP61M1_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__31862),
            .in2(N__31850),
            .in3(N__31838),
            .lcout(\ALU.mult_5_13 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\ALU.mult_5_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_221_c_RNI6Q7IO1_LC_14_9_1 .C_ON=1'b1;
    defparam \ALU.mult_221_c_RNI6Q7IO1_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_221_c_RNI6Q7IO1_LC_14_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_221_c_RNI6Q7IO1_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__31835),
            .in2(N__31826),
            .in3(N__31811),
            .lcout(\ALU.mult_5_14 ),
            .ltout(),
            .carryin(\ALU.mult_5_c13 ),
            .carryout(\ALU.mult_5_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_227_c_RNIBPRV92_LC_14_9_2 .C_ON=1'b0;
    defparam \ALU.mult_227_c_RNIBPRV92_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_227_c_RNIBPRV92_LC_14_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_227_c_RNIBPRV92_LC_14_9_2  (
            .in0(N__31808),
            .in1(N__31802),
            .in2(N__31787),
            .in3(N__31769),
            .lcout(\ALU.mult_227_c_RNIBPRVZ0Z92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILTVJG3_3_LC_14_9_3 .C_ON=1'b0;
    defparam \ALU.d_RNILTVJG3_3_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILTVJG3_3_LC_14_9_3 .LUT_INIT=16'b1000000010001111;
    LogicCell40 \ALU.d_RNILTVJG3_3_LC_14_9_3  (
            .in0(N__57238),
            .in1(N__56465),
            .in2(N__70016),
            .in3(N__31766),
            .lcout(\ALU.d_RNILTVJG3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_239_c_RNO_0_LC_14_9_4 .C_ON=1'b0;
    defparam \ALU.mult_239_c_RNO_0_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_239_c_RNO_0_LC_14_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_239_c_RNO_0_LC_14_9_4  (
            .in0(N__62269),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66570),
            .lcout(\ALU.mult_239_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_239_c_RNO_LC_14_9_6 .C_ON=1'b0;
    defparam \ALU.mult_239_c_RNO_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_239_c_RNO_LC_14_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_239_c_RNO_LC_14_9_6  (
            .in0(N__65828),
            .in1(N__62314),
            .in2(N__66696),
            .in3(N__62523),
            .lcout(\ALU.mult_239_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_5_c_RNI6LDHN2_LC_14_10_0 .C_ON=1'b1;
    defparam \ALU.mult_5_c_RNI6LDHN2_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_5_c_RNI6LDHN2_LC_14_10_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ALU.mult_5_c_RNI6LDHN2_LC_14_10_0  (
            .in0(N__31714),
            .in1(N__33806),
            .in2(N__31715),
            .in3(_gnd_net_),
            .lcout(\ALU.mult_2 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\ALU.mult_17_c2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_388_c_RNI23SO83_LC_14_10_1 .C_ON=1'b1;
    defparam \ALU.mult_388_c_RNI23SO83_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_388_c_RNI23SO83_LC_14_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_388_c_RNI23SO83_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__34112),
            .in2(N__31700),
            .in3(N__31691),
            .lcout(\ALU.mult_3 ),
            .ltout(),
            .carryin(\ALU.mult_17_c2 ),
            .carryout(\ALU.mult_17_c3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_391_c_RNIQB68P3_LC_14_10_2 .C_ON=1'b1;
    defparam \ALU.mult_391_c_RNIQB68P3_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_391_c_RNIQB68P3_LC_14_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_391_c_RNIQB68P3_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__32057),
            .in2(N__32045),
            .in3(N__32036),
            .lcout(\ALU.mult_17_4 ),
            .ltout(),
            .carryin(\ALU.mult_17_c3 ),
            .carryout(\ALU.mult_17_c4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_394_c_RNIP20HH3_LC_14_10_3 .C_ON=1'b1;
    defparam \ALU.mult_394_c_RNIP20HH3_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_394_c_RNIP20HH3_LC_14_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_394_c_RNIP20HH3_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__32033),
            .in2(N__32027),
            .in3(N__32012),
            .lcout(\ALU.mult_17_5 ),
            .ltout(),
            .carryin(\ALU.mult_17_c4 ),
            .carryout(\ALU.mult_17_c5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_397_c_RNI951U83_LC_14_10_4 .C_ON=1'b1;
    defparam \ALU.mult_397_c_RNI951U83_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_397_c_RNI951U83_LC_14_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_397_c_RNI951U83_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(N__32009),
            .in2(N__32000),
            .in3(N__31985),
            .lcout(\ALU.mult_17_6 ),
            .ltout(),
            .carryin(\ALU.mult_17_c5 ),
            .carryout(\ALU.mult_17_c6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_400_c_RNI1KKT93_LC_14_10_5 .C_ON=1'b1;
    defparam \ALU.mult_400_c_RNI1KKT93_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_400_c_RNI1KKT93_LC_14_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_400_c_RNI1KKT93_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__31982),
            .in2(N__31976),
            .in3(N__31961),
            .lcout(\ALU.mult_17_7 ),
            .ltout(),
            .carryin(\ALU.mult_17_c6 ),
            .carryout(\ALU.mult_17_c7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_403_c_RNINS3F83_LC_14_10_6 .C_ON=1'b1;
    defparam \ALU.mult_403_c_RNINS3F83_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_403_c_RNINS3F83_LC_14_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_403_c_RNINS3F83_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__31958),
            .in2(N__31952),
            .in3(N__31937),
            .lcout(\ALU.mult_17_8 ),
            .ltout(),
            .carryin(\ALU.mult_17_c7 ),
            .carryout(\ALU.mult_17_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_406_c_RNITD5193_LC_14_10_7 .C_ON=1'b1;
    defparam \ALU.mult_406_c_RNITD5193_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_406_c_RNITD5193_LC_14_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_406_c_RNITD5193_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__31934),
            .in2(N__31925),
            .in3(N__31910),
            .lcout(\ALU.mult_17_9 ),
            .ltout(),
            .carryin(\ALU.mult_17_c8 ),
            .carryout(\ALU.mult_17_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_409_c_RNIRS5V93_LC_14_11_0 .C_ON=1'b1;
    defparam \ALU.mult_409_c_RNIRS5V93_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_409_c_RNIRS5V93_LC_14_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_409_c_RNIRS5V93_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__31907),
            .in2(N__31898),
            .in3(N__31889),
            .lcout(\ALU.mult_17_10 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\ALU.mult_17_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_412_c_RNI68PMD3_LC_14_11_1 .C_ON=1'b1;
    defparam \ALU.mult_412_c_RNI68PMD3_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_412_c_RNI68PMD3_LC_14_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_412_c_RNI68PMD3_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__31886),
            .in2(N__31880),
            .in3(N__31865),
            .lcout(\ALU.mult_17_11 ),
            .ltout(),
            .carryin(\ALU.mult_17_c10 ),
            .carryout(\ALU.mult_17_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_415_c_RNIET5KE3_LC_14_11_2 .C_ON=1'b1;
    defparam \ALU.mult_415_c_RNIET5KE3_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_415_c_RNIET5KE3_LC_14_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_415_c_RNIET5KE3_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(N__32189),
            .in2(N__32183),
            .in3(N__32168),
            .lcout(\ALU.mult_17_12 ),
            .ltout(),
            .carryin(\ALU.mult_17_c11 ),
            .carryout(\ALU.mult_17_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_418_c_RNITRJ9K3_LC_14_11_3 .C_ON=1'b1;
    defparam \ALU.mult_418_c_RNITRJ9K3_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_418_c_RNITRJ9K3_LC_14_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_418_c_RNITRJ9K3_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__32165),
            .in2(N__32159),
            .in3(N__32144),
            .lcout(\ALU.mult_17_13 ),
            .ltout(),
            .carryin(\ALU.mult_17_c12 ),
            .carryout(\ALU.mult_17_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_421_c_RNIRNI2G3_LC_14_11_4 .C_ON=1'b1;
    defparam \ALU.mult_421_c_RNIRNI2G3_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_421_c_RNIRNI2G3_LC_14_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_421_c_RNIRNI2G3_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__32141),
            .in2(N__32135),
            .in3(N__32120),
            .lcout(\ALU.mult_17_14 ),
            .ltout(),
            .carryin(\ALU.mult_17_c13 ),
            .carryout(\ALU.mult_17_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_424_c_RNIUVTAL4_LC_14_11_5 .C_ON=1'b0;
    defparam \ALU.mult_424_c_RNIUVTAL4_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_424_c_RNIUVTAL4_LC_14_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_424_c_RNIUVTAL4_LC_14_11_5  (
            .in0(N__32117),
            .in1(N__32108),
            .in2(N__33815),
            .in3(N__32102),
            .lcout(\ALU.mult_424_c_RNIUVTALZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHU6RL_1_LC_14_11_7 .C_ON=1'b0;
    defparam \ALU.d_RNIHU6RL_1_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHU6RL_1_LC_14_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIHU6RL_1_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__65521),
            .in2(_gnd_net_),
            .in3(N__68728),
            .lcout(\ALU.d_RNIHU6RLZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2E4JE1_4_LC_14_12_0 .C_ON=1'b0;
    defparam \ALU.d_RNI2E4JE1_4_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2E4JE1_4_LC_14_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI2E4JE1_4_LC_14_12_0  (
            .in0(N__65715),
            .in1(N__68660),
            .in2(N__59624),
            .in3(N__59903),
            .lcout(\ALU.d_RNI2E4JE1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISLOMK_0_1_LC_14_12_1 .C_ON=1'b0;
    defparam \ALU.d_RNISLOMK_0_1_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISLOMK_0_1_LC_14_12_1 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \ALU.d_RNISLOMK_0_1_LC_14_12_1  (
            .in0(N__34100),
            .in1(N__34685),
            .in2(N__53249),
            .in3(N__34067),
            .lcout(\ALU.addsub_axb_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFCCRV4_4_LC_14_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNIFCCRV4_4_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFCCRV4_4_LC_14_12_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNIFCCRV4_4_LC_14_12_4  (
            .in0(N__39229),
            .in1(N__68661),
            .in2(_gnd_net_),
            .in3(N__32078),
            .lcout(\ALU.N_920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_5_c_RNO_LC_14_12_5 .C_ON=1'b0;
    defparam \ALU.mult_5_c_RNO_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_5_c_RNO_LC_14_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_5_c_RNO_LC_14_12_5  (
            .in0(N__60539),
            .in1(N__65446),
            .in2(N__66755),
            .in3(N__65711),
            .lcout(\ALU.mult_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI290AE1_0_LC_14_12_6 .C_ON=1'b0;
    defparam \ALU.d_RNI290AE1_0_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI290AE1_0_LC_14_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI290AE1_0_LC_14_12_6  (
            .in0(N__65445),
            .in1(N__68659),
            .in2(N__65826),
            .in3(N__60540),
            .lcout(\ALU.d_RNI290AE1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5MTIO_1_LC_14_12_7 .C_ON=1'b0;
    defparam \ALU.d_RNI5MTIO_1_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5MTIO_1_LC_14_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI5MTIO_1_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__65444),
            .in2(_gnd_net_),
            .in3(N__65710),
            .lcout(\ALU.d_RNI5MTIOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNICT0U1_2_LC_14_13_0 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNICT0U1_2_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNICT0U1_2_LC_14_13_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \CONTROL.busState_1_RNICT0U1_2_LC_14_13_0  (
            .in0(N__49519),
            .in1(N__50337),
            .in2(N__32357),
            .in3(N__50197),
            .lcout(busState_1_RNICT0U1_2),
            .ltout(busState_1_RNICT0U1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8U1VH_2_LC_14_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNI8U1VH_2_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8U1VH_2_LC_14_13_1 .LUT_INIT=16'b1111011111000100;
    LogicCell40 \ALU.d_RNI8U1VH_2_LC_14_13_1  (
            .in0(N__32758),
            .in1(N__53204),
            .in2(N__32396),
            .in3(N__32937),
            .lcout(\ALU.status_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8U1VH_0_2_LC_14_13_3 .C_ON=1'b0;
    defparam \ALU.d_RNI8U1VH_0_2_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8U1VH_0_2_LC_14_13_3 .LUT_INIT=16'b1111011111000100;
    LogicCell40 \ALU.d_RNI8U1VH_0_2_LC_14_13_3  (
            .in0(N__32759),
            .in1(N__53205),
            .in2(N__32393),
            .in3(N__32938),
            .lcout(\ALU.lshift_15_0_sx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNILM6T5_2_LC_14_13_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNILM6T5_2_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNILM6T5_2_LC_14_13_4 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \CONTROL.busState_1_RNILM6T5_2_LC_14_13_4  (
            .in0(N__66228),
            .in1(N__32392),
            .in2(N__49582),
            .in3(N__50198),
            .lcout(N_227_0),
            .ltout(N_227_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_2_c_RNO_LC_14_13_5 .C_ON=1'b0;
    defparam \ALU.status_18_cry_2_c_RNO_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_2_c_RNO_LC_14_13_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \ALU.status_18_cry_2_c_RNO_LC_14_13_5  (
            .in0(N__53216),
            .in1(N__66229),
            .in2(N__32381),
            .in3(N__32939),
            .lcout(\ALU.status_18_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI8MJL_2_LC_14_13_6 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI8MJL_2_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI8MJL_2_LC_14_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI8MJL_2_LC_14_13_6  (
            .in0(N__32330),
            .in1(N__32347),
            .in2(_gnd_net_),
            .in3(N__32322),
            .lcout(DROM_ROMDATA_dintern_2ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_2_LC_14_13_7 .C_ON=1'b0;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_2_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \DROM.ROMDATA.dintern_0_0_OLD_ne_2_LC_14_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DROM.ROMDATA.dintern_0_0_OLD_ne_2_LC_14_13_7  (
            .in0(N__32348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DROM.ROMDATA.dintern_0_0_OLDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C_net ),
            .ce(N__32323),
            .sr(_gnd_net_));
    defparam \ALU.e_2_LC_14_14_0 .C_ON=1'b0;
    defparam \ALU.e_2_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.e_2_LC_14_14_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.e_2_LC_14_14_0  (
            .in0(N__39456),
            .in1(N__39604),
            .in2(_gnd_net_),
            .in3(N__39516),
            .lcout(\ALU.eZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73153),
            .ce(N__69244),
            .sr(_gnd_net_));
    defparam \ALU.e_4_LC_14_14_1 .C_ON=1'b0;
    defparam \ALU.e_4_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.e_4_LC_14_14_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.e_4_LC_14_14_1  (
            .in0(N__39391),
            .in1(N__57420),
            .in2(_gnd_net_),
            .in3(N__42551),
            .lcout(\ALU.eZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73153),
            .ce(N__69244),
            .sr(_gnd_net_));
    defparam \ALU.e_5_LC_14_14_2 .C_ON=1'b0;
    defparam \ALU.e_5_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.e_5_LC_14_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_5_LC_14_14_2  (
            .in0(N__57419),
            .in1(N__52627),
            .in2(_gnd_net_),
            .in3(N__39322),
            .lcout(\ALU.eZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73153),
            .ce(N__69244),
            .sr(_gnd_net_));
    defparam \ALU.e_6_LC_14_14_3 .C_ON=1'b0;
    defparam \ALU.e_6_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.e_6_LC_14_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_6_LC_14_14_3  (
            .in0(N__43067),
            .in1(N__43121),
            .in2(_gnd_net_),
            .in3(N__42991),
            .lcout(\ALU.eZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73153),
            .ce(N__69244),
            .sr(_gnd_net_));
    defparam \ALU.e_3_LC_14_14_4 .C_ON=1'b0;
    defparam \ALU.e_3_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.e_3_LC_14_14_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.e_3_LC_14_14_4  (
            .in0(N__58799),
            .in1(N__58757),
            .in2(_gnd_net_),
            .in3(N__58666),
            .lcout(\ALU.eZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73153),
            .ce(N__69244),
            .sr(_gnd_net_));
    defparam \ALU.e_10_LC_14_14_5 .C_ON=1'b0;
    defparam \ALU.e_10_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \ALU.e_10_LC_14_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_10_LC_14_14_5  (
            .in0(N__58510),
            .in1(N__58371),
            .in2(_gnd_net_),
            .in3(N__58300),
            .lcout(\ALU.eZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73153),
            .ce(N__69244),
            .sr(_gnd_net_));
    defparam \ALU.e_11_LC_14_14_6 .C_ON=1'b0;
    defparam \ALU.e_11_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \ALU.e_11_LC_14_14_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.e_11_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__58194),
            .in2(N__58126),
            .in3(N__58058),
            .lcout(\ALU.eZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73153),
            .ce(N__69244),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_14_14_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_14_14_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_14_14_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_14_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIAHH51_6_LC_14_15_0 .C_ON=1'b0;
    defparam \ALU.b_RNIAHH51_6_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIAHH51_6_LC_14_15_0 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \ALU.b_RNIAHH51_6_LC_14_15_0  (
            .in0(N__43912),
            .in1(N__70603),
            .in2(N__39895),
            .in3(N__34556),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMOPK1_6_LC_14_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIMOPK1_6_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMOPK1_6_LC_14_15_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIMOPK1_6_LC_14_15_1  (
            .in0(N__37434),
            .in1(N__36055),
            .in2(N__32735),
            .in3(N__47188),
            .lcout(\ALU.N_1139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI8BB31_6_LC_14_15_2 .C_ON=1'b0;
    defparam \ALU.e_RNI8BB31_6_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI8BB31_6_LC_14_15_2 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.e_RNI8BB31_6_LC_14_15_2  (
            .in0(N__43913),
            .in1(N__42941),
            .in2(N__32728),
            .in3(N__34557),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIICD02_6_LC_14_15_3 .C_ON=1'b0;
    defparam \ALU.c_RNIICD02_6_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIICD02_6_LC_14_15_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNIICD02_6_LC_14_15_3  (
            .in0(N__35764),
            .in1(N__35833),
            .in2(N__32708),
            .in3(N__47189),
            .lcout(),
            .ltout(\ALU.N_1091_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIB9LU3_6_LC_14_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNIB9LU3_6_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIB9LU3_6_LC_14_15_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIB9LU3_6_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__54110),
            .in2(N__32705),
            .in3(N__32702),
            .lcout(aluOut_6),
            .ltout(aluOut_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIR3N75_6_LC_14_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNIR3N75_6_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIR3N75_6_LC_14_15_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.d_RNIR3N75_6_LC_14_15_5  (
            .in0(N__53144),
            .in1(N__49563),
            .in2(N__32696),
            .in3(N__50143),
            .lcout(\ALU.d_RNIR3N75Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI3N941_1_LC_14_16_0 .C_ON=1'b0;
    defparam \ALU.b_RNI3N941_1_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI3N941_1_LC_14_16_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.b_RNI3N941_1_LC_14_16_0  (
            .in0(N__47144),
            .in1(N__49164),
            .in2(N__47271),
            .in3(N__48410),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5KHJ1_1_LC_14_16_1 .C_ON=1'b0;
    defparam \ALU.d_RNI5KHJ1_1_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5KHJ1_1_LC_14_16_1 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNI5KHJ1_1_LC_14_16_1  (
            .in0(N__37512),
            .in1(N__47145),
            .in2(N__32675),
            .in3(N__52165),
            .lcout(ALU_N_1134),
            .ltout(ALU_N_1134_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_RNIR8FK7_0_LC_14_16_2 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_RNIR8FK7_0_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_ne_RNIR8FK7_0_LC_14_16_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \CONTROL.operand1_ne_RNIR8FK7_0_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__32669),
            .in2(N__32672),
            .in3(N__34286),
            .lcout(operand1_ne_RNIR8FK7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_RNIBQE03_0_LC_14_16_3 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_RNIBQE03_0_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_ne_RNIBQE03_0_LC_14_16_3 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \CONTROL.operand1_ne_RNIBQE03_0_LC_14_16_3  (
            .in0(N__54113),
            .in1(N__50131),
            .in2(N__49579),
            .in3(N__34298),
            .lcout(\CONTROL.operand1_ne_RNIBQE03Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI9P5V3_2_LC_14_16_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI9P5V3_2_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI9P5V3_2_LC_14_16_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \CONTROL.busState_1_RNI9P5V3_2_LC_14_16_4  (
            .in0(N__50132),
            .in1(N__49512),
            .in2(_gnd_net_),
            .in3(N__66127),
            .lcout(busState_1_RNI9P5V3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI1H321_1_LC_14_16_5 .C_ON=1'b0;
    defparam \ALU.e_RNI1H321_1_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI1H321_1_LC_14_16_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.e_RNI1H321_1_LC_14_16_5  (
            .in0(N__37234),
            .in1(N__47142),
            .in2(N__46351),
            .in3(N__47246),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI185V1_1_LC_14_16_6 .C_ON=1'b0;
    defparam \ALU.c_RNI185V1_1_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI185V1_1_LC_14_16_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNI185V1_1_LC_14_16_6  (
            .in0(N__47143),
            .in1(N__48942),
            .in2(N__32747),
            .in3(N__46462),
            .lcout(ALU_N_1086),
            .ltout(ALU_N_1086_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI905S3_1_LC_14_16_7 .C_ON=1'b0;
    defparam \ALU.d_RNI905S3_1_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI905S3_1_LC_14_16_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNI905S3_1_LC_14_16_7  (
            .in0(N__54114),
            .in1(_gnd_net_),
            .in2(N__32744),
            .in3(N__32741),
            .lcout(aluOut_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_1_LC_14_17_0 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_1_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_ne_1_LC_14_17_0 .LUT_INIT=16'b0001111100001110;
    LogicCell40 \CONTROL.operand1_ne_1_LC_14_17_0  (
            .in0(N__79431),
            .in1(N__72722),
            .in2(N__34433),
            .in3(N__54362),
            .lcout(aluOperand1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_ne_1C_net ),
            .ce(N__36240),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_fast_ne_2_LC_14_17_1 .C_ON=1'b0;
    defparam \CONTROL.operand1_fast_ne_2_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_fast_ne_2_LC_14_17_1 .LUT_INIT=16'b0100111101001010;
    LogicCell40 \CONTROL.operand1_fast_ne_2_LC_14_17_1  (
            .in0(N__72721),
            .in1(N__50487),
            .in2(N__45059),
            .in3(N__41052),
            .lcout(aluOperand1_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_ne_1C_net ),
            .ce(N__36240),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_2_rep1_ne_LC_14_17_2 .C_ON=1'b0;
    defparam \CONTROL.operand1_2_rep1_ne_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_2_rep1_ne_LC_14_17_2 .LUT_INIT=16'b0101010111100100;
    LogicCell40 \CONTROL.operand1_2_rep1_ne_LC_14_17_2  (
            .in0(N__45050),
            .in1(N__41053),
            .in2(N__50494),
            .in3(N__72723),
            .lcout(aluOperand1_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_ne_1C_net ),
            .ce(N__36240),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_2_rep2_ne_LC_14_17_3 .C_ON=1'b0;
    defparam \CONTROL.operand1_2_rep2_ne_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_2_rep2_ne_LC_14_17_3 .LUT_INIT=16'b0100111101001010;
    LogicCell40 \CONTROL.operand1_2_rep2_ne_LC_14_17_3  (
            .in0(N__72720),
            .in1(N__50486),
            .in2(N__45058),
            .in3(N__41051),
            .lcout(aluOperand1_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_ne_1C_net ),
            .ce(N__36240),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_2_LC_14_17_4 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_2_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_ne_2_LC_14_17_4 .LUT_INIT=16'b0101010111100100;
    LogicCell40 \CONTROL.operand1_ne_2_LC_14_17_4  (
            .in0(N__45051),
            .in1(N__41054),
            .in2(N__50495),
            .in3(N__72724),
            .lcout(aluOperand1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_ne_1C_net ),
            .ce(N__36240),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPTT4O_0_8_LC_14_17_5 .C_ON=1'b0;
    defparam \ALU.d_RNIPTT4O_0_8_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPTT4O_0_8_LC_14_17_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNIPTT4O_0_8_LC_14_17_5  (
            .in0(N__61881),
            .in1(N__62191),
            .in2(_gnd_net_),
            .in3(N__66569),
            .lcout(\ALU.N_610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHD7AO_7_LC_14_17_7 .C_ON=1'b0;
    defparam \ALU.d_RNIHD7AO_7_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHD7AO_7_LC_14_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIHD7AO_7_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__62190),
            .in2(_gnd_net_),
            .in3(N__65931),
            .lcout(\ALU.d_RNIHD7AOZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNICDG51_0_LC_14_18_0 .C_ON=1'b0;
    defparam \ALU.b_RNICDG51_0_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNICDG51_0_LC_14_18_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.b_RNICDG51_0_LC_14_18_0  (
            .in0(N__48376),
            .in1(N__36315),
            .in2(N__49132),
            .in3(N__32809),
            .lcout(\ALU.dout_6_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_RNIHKCU2_0_LC_14_18_1 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_RNIHKCU2_0_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_ne_RNIHKCU2_0_LC_14_18_1 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \CONTROL.operand1_ne_RNIHKCU2_0_LC_14_18_1  (
            .in0(N__50103),
            .in1(N__54061),
            .in2(N__49528),
            .in3(N__32767),
            .lcout(),
            .ltout(\CONTROL.operand1_ne_RNIHKCU2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_RNIDN8E7_0_LC_14_18_2 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_RNIDN8E7_0_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_ne_RNIDN8E7_0_LC_14_18_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \CONTROL.operand1_ne_RNIDN8E7_0_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__32776),
            .in2(N__32849),
            .in3(N__32783),
            .lcout(operand1_ne_RNIDN8E7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBEFH1_0_LC_14_18_3 .C_ON=1'b0;
    defparam \ALU.d_RNIBEFH1_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBEFH1_0_LC_14_18_3 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \ALU.d_RNIBEFH1_0_LC_14_18_3  (
            .in0(N__51971),
            .in1(N__54236),
            .in2(N__37561),
            .in3(N__32831),
            .lcout(ALU_N_1133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIA7A31_0_LC_14_18_4 .C_ON=1'b0;
    defparam \ALU.e_RNIA7A31_0_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIA7A31_0_LC_14_18_4 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \ALU.e_RNIA7A31_0_LC_14_18_4  (
            .in0(N__46324),
            .in1(N__32810),
            .in2(N__37589),
            .in3(N__36316),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI723T1_0_LC_14_18_5 .C_ON=1'b0;
    defparam \ALU.c_RNI723T1_0_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI723T1_0_LC_14_18_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNI723T1_0_LC_14_18_5  (
            .in0(N__48900),
            .in1(N__46433),
            .in2(N__32789),
            .in3(N__54235),
            .lcout(ALU_N_1085),
            .ltout(ALU_N_1085_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_RNIHKCU2_0_0_LC_14_18_6 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_RNIHKCU2_0_0_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_ne_RNIHKCU2_0_0_LC_14_18_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \CONTROL.operand1_ne_RNIHKCU2_0_0_LC_14_18_6  (
            .in0(N__54060),
            .in1(N__49431),
            .in2(N__32786),
            .in3(N__50102),
            .lcout(\CONTROL.operand1_ne_RNIHKCU2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILK0O3_0_LC_14_18_7 .C_ON=1'b0;
    defparam \ALU.d_RNILK0O3_0_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILK0O3_0_LC_14_18_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNILK0O3_0_LC_14_18_7  (
            .in0(N__32777),
            .in1(N__54062),
            .in2(_gnd_net_),
            .in3(N__32768),
            .lcout(aluOut_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI1C5B1_2_LC_14_19_0 .C_ON=1'b0;
    defparam \ALU.b_RNI1C5B1_2_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI1C5B1_2_LC_14_19_0 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.b_RNI1C5B1_2_LC_14_19_0  (
            .in0(N__53584),
            .in1(N__35632),
            .in2(N__39422),
            .in3(N__53480),
            .lcout(\ALU.operand2_6_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIV5V81_2_LC_14_19_1 .C_ON=1'b0;
    defparam \ALU.e_RNIV5V81_2_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIV5V81_2_LC_14_19_1 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNIV5V81_2_LC_14_19_1  (
            .in0(N__34352),
            .in1(N__53583),
            .in2(N__34334),
            .in3(N__53479),
            .lcout(),
            .ltout(\ALU.operand2_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI0C2B2_2_LC_14_19_2 .C_ON=1'b0;
    defparam \ALU.c_RNI0C2B2_2_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI0C2B2_2_LC_14_19_2 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNI0C2B2_2_LC_14_19_2  (
            .in0(N__35566),
            .in1(N__35876),
            .in2(N__32960),
            .in3(N__53429),
            .lcout(\ALU.N_1199 ),
            .ltout(\ALU.N_1199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJ1JO4_2_LC_14_19_3 .C_ON=1'b0;
    defparam \ALU.c_RNIJ1JO4_2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJ1JO4_2_LC_14_19_3 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \ALU.c_RNIJ1JO4_2_LC_14_19_3  (
            .in0(N__43494),
            .in1(N__71320),
            .in2(N__32957),
            .in3(N__53941),
            .lcout(\ALU.c_RNIJ1JO4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJ1JO4_0_2_LC_14_19_4 .C_ON=1'b0;
    defparam \ALU.c_RNIJ1JO4_0_2_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJ1JO4_0_2_LC_14_19_4 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \ALU.c_RNIJ1JO4_0_2_LC_14_19_4  (
            .in0(N__53942),
            .in1(N__32954),
            .in2(N__71384),
            .in3(N__43495),
            .lcout(),
            .ltout(\ALU.c_RNIJ1JO4_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIARKGB_2_LC_14_19_5 .C_ON=1'b0;
    defparam \ALU.d_RNIARKGB_2_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIARKGB_2_LC_14_19_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIARKGB_2_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__32918),
            .in2(N__32948),
            .in3(N__32945),
            .lcout(\ALU.d_RNIARKGBZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4OEV1_2_LC_14_19_6 .C_ON=1'b0;
    defparam \ALU.d_RNI4OEV1_2_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4OEV1_2_LC_14_19_6 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \ALU.d_RNI4OEV1_2_LC_14_19_6  (
            .in0(N__36083),
            .in1(N__32924),
            .in2(N__34403),
            .in3(N__53430),
            .lcout(\ALU.N_1247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI48DU_13_LC_14_20_0 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI48DU_13_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI48DU_13_LC_14_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNI48DU_13_LC_14_20_0  (
            .in0(N__32912),
            .in1(N__43669),
            .in2(_gnd_net_),
            .in3(N__50009),
            .lcout(),
            .ltout(\CONTROL.N_174_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIEJJS1_2_LC_14_20_1 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIEJJS1_2_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIEJJS1_2_LC_14_20_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \CONTROL.busState_1_RNIEJJS1_2_LC_14_20_1  (
            .in0(N__50010),
            .in1(N__32891),
            .in2(N__32867),
            .in3(N__49341),
            .lcout(\CONTROL.N_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIAHKF1_2_LC_14_20_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIAHKF1_2_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIAHKF1_2_LC_14_20_2 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \CONTROL.busState_1_RNIAHKF1_2_LC_14_20_2  (
            .in0(N__49340),
            .in1(N__33200),
            .in2(N__33191),
            .in3(N__50008),
            .lcout(\CONTROL.N_185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_2_LC_14_20_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_2_LC_14_20_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.busState_1_2_LC_14_20_3 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \CONTROL.busState_1_2_LC_14_20_3  (
            .in0(N__41615),
            .in1(N__40625),
            .in2(N__49505),
            .in3(N__34697),
            .lcout(busState_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.busState_1_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIU83C1_0_2_LC_14_20_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIU83C1_0_2_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIU83C1_0_2_LC_14_20_4 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \CONTROL.busState_1_RNIU83C1_0_2_LC_14_20_4  (
            .in0(N__49342),
            .in1(N__37993),
            .in2(N__33139),
            .in3(N__50011),
            .lcout(\CONTROL.busState_1_RNIU83C1_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIOKAQ1_2_LC_14_20_6 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIOKAQ1_2_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIOKAQ1_2_LC_14_20_6 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \CONTROL.busState_1_RNIOKAQ1_2_LC_14_20_6  (
            .in0(N__49339),
            .in1(N__34829),
            .in2(N__33086),
            .in3(N__50007),
            .lcout(N_179),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIBKBS7_0_LC_14_20_7 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIBKBS7_0_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIBKBS7_0_LC_14_20_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \CONTROL.busState_1_RNIBKBS7_0_LC_14_20_7  (
            .in0(N__33065),
            .in1(N__33380),
            .in2(_gnd_net_),
            .in3(N__49802),
            .lcout(bus_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNILAEH1_2_LC_14_21_0 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNILAEH1_2_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNILAEH1_2_LC_14_21_0 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \CONTROL.busState_1_RNILAEH1_2_LC_14_21_0  (
            .in0(N__49946),
            .in1(N__49322),
            .in2(N__32993),
            .in3(N__32984),
            .lcout(\CONTROL.busState_1_RNILAEH1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNIUDOJ_1_LC_14_21_1 .C_ON=1'b0;
    defparam \CONTROL.dout_RNIUDOJ_1_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNIUDOJ_1_LC_14_21_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNIUDOJ_1_LC_14_21_1  (
            .in0(N__33017),
            .in1(N__50662),
            .in2(_gnd_net_),
            .in3(N__49942),
            .lcout(N_162),
            .ltout(N_162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.combOperand2_d_bm_1_LC_14_21_2 .C_ON=1'b0;
    defparam \ALU.combOperand2_d_bm_1_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \ALU.combOperand2_d_bm_1_LC_14_21_2 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \ALU.combOperand2_d_bm_1_LC_14_21_2  (
            .in0(N__49943),
            .in1(N__32983),
            .in2(N__32963),
            .in3(N__49320),
            .lcout(\ALU.combOperand2_d_bmZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_1_LC_14_21_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_1_LC_14_21_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.busState_1_1_LC_14_21_3 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \CONTROL.busState_1_1_LC_14_21_3  (
            .in0(N__34868),
            .in1(N__40637),
            .in2(N__50186),
            .in3(N__34712),
            .lcout(busState_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.busState_1_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_a7_3_LC_14_21_4 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_a7_3_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_a7_3_LC_14_21_4 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \CONTROL.g0_3_i_a7_3_LC_14_21_4  (
            .in0(N__39779),
            .in1(N__45410),
            .in2(N__45515),
            .in3(N__54660),
            .lcout(\CONTROL.g0_3_i_a7_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIRU6J1_2_LC_14_21_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIRU6J1_2_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIRU6J1_2_LC_14_21_5 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \CONTROL.busState_1_RNIRU6J1_2_LC_14_21_5  (
            .in0(N__49323),
            .in1(N__33344),
            .in2(N__33353),
            .in3(N__49947),
            .lcout(\CONTROL.N_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI2IOJ_3_LC_14_21_6 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI2IOJ_3_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI2IOJ_3_LC_14_21_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.dout_RNI2IOJ_3_LC_14_21_6  (
            .in0(N__49944),
            .in1(N__33374),
            .in2(_gnd_net_),
            .in3(N__45280),
            .lcout(N_164),
            .ltout(N_164_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.combOperand2_d_bm_3_LC_14_21_7 .C_ON=1'b0;
    defparam \ALU.combOperand2_d_bm_3_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \ALU.combOperand2_d_bm_3_LC_14_21_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \ALU.combOperand2_d_bm_3_LC_14_21_7  (
            .in0(N__49321),
            .in1(N__33343),
            .in2(N__33320),
            .in3(N__49945),
            .lcout(\ALU.combOperand2_d_bmZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_0_LC_14_22_0 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_0_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_0_LC_14_22_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \CONTROL.romAddReg_7_0_LC_14_22_0  (
            .in0(N__71828),
            .in1(N__33306),
            .in2(N__48914),
            .in3(N__72178),
            .lcout(CONTROL_romAddReg_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_17dflt_LC_14_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_17dflt_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_17dflt_LC_14_22_1 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_17dflt_LC_14_22_1  (
            .in0(N__72177),
            .in1(N__38869),
            .in2(N__63968),
            .in3(N__72681),
            .lcout(controlWord_17),
            .ltout(controlWord_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_1_LC_14_22_2 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_1_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_1_LC_14_22_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \CONTROL.romAddReg_7_1_LC_14_22_2  (
            .in0(N__71829),
            .in1(N__48950),
            .in2(N__33236),
            .in3(N__72179),
            .lcout(CONTROL_romAddReg_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m375_am_LC_14_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m375_am_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m375_am_LC_14_22_3 .LUT_INIT=16'b0000001110001011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m375_am_LC_14_22_3  (
            .in0(N__74480),
            .in1(N__76593),
            .in2(N__73394),
            .in3(N__75969),
            .lcout(\PROM.ROMDATA.m375_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_1_LC_14_22_6 .C_ON=1'b0;
    defparam \CONTROL.dout_1_LC_14_22_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_1_LC_14_22_6 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \CONTROL.dout_1_LC_14_22_6  (
            .in0(N__72682),
            .in1(N__63967),
            .in2(N__38873),
            .in3(N__72180),
            .lcout(\CONTROL.ctrlOut_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_1C_net ),
            .ce(N__44434),
            .sr(_gnd_net_));
    defparam \CONTROL.busState104_2_LC_14_22_7 .C_ON=1'b0;
    defparam \CONTROL.busState104_2_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState104_2_LC_14_22_7 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \CONTROL.busState104_2_LC_14_22_7  (
            .in0(N__72176),
            .in1(N__71827),
            .in2(_gnd_net_),
            .in3(N__44679),
            .lcout(\CONTROL.N_384_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_35_LC_14_23_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_35_LC_14_23_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_35_LC_14_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \CONTROL.programCounter_ret_35_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__50841),
            .in2(_gnd_net_),
            .in3(N__50906),
            .lcout(CONTROL_programCounter11_reto),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73232),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI7IMQ_15_LC_14_23_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI7IMQ_15_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI7IMQ_15_LC_14_23_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI7IMQ_15_LC_14_23_1  (
            .in0(N__33440),
            .in1(N__33422),
            .in2(_gnd_net_),
            .in3(N__42082),
            .lcout(\CONTROL.N_430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState98_1_1_0_0_LC_14_23_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState98_1_1_0_0_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState98_1_1_0_0_LC_14_23_2 .LUT_INIT=16'b1111111110111001;
    LogicCell40 \CONTROL.un1_busState98_1_1_0_0_LC_14_23_2  (
            .in0(N__44702),
            .in1(N__36680),
            .in2(N__41261),
            .in3(N__54655),
            .lcout(\CONTROL.un1_busState98_1_1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_15_LC_14_23_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_15_LC_14_23_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_15_LC_14_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_15_LC_14_23_3  (
            .in0(N__33461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73232),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_15_LC_14_23_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_15_LC_14_23_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_15_LC_14_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_15_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33434),
            .lcout(\CONTROL.dout_reto_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73232),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m465_am_LC_14_23_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m465_am_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m465_am_LC_14_23_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m465_am_LC_14_23_5  (
            .in0(N__74491),
            .in1(N__76633),
            .in2(_gnd_net_),
            .in3(N__75973),
            .lcout(\PROM.ROMDATA.m465_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m299_LC_14_23_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m299_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m299_LC_14_23_6 .LUT_INIT=16'b0000110000100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m299_LC_14_23_6  (
            .in0(N__78853),
            .in1(N__78060),
            .in2(N__76004),
            .in3(N__77308),
            .lcout(\PROM.ROMDATA.m299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_7_LC_14_23_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_7_LC_14_23_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_7_LC_14_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_7_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33401),
            .lcout(\CONTROL.dout_reto_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73232),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_0_LC_14_24_1 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_0_LC_14_24_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_0_LC_14_24_1 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \CONTROL.tempCounter_0_LC_14_24_1  (
            .in0(N__47408),
            .in1(N__73636),
            .in2(_gnd_net_),
            .in3(N__50969),
            .lcout(\CONTROL.tempCounterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_0C_net ),
            .ce(N__34954),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_5_LC_14_24_2 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_5_LC_14_24_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_5_LC_14_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_5_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41740),
            .lcout(\CONTROL.tempCounterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_0C_net ),
            .ce(N__34954),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_3_LC_14_24_3 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_3_LC_14_24_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_3_LC_14_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_3_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51148),
            .lcout(\CONTROL.tempCounterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_0C_net ),
            .ce(N__34954),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_8_LC_14_24_4 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_8_LC_14_24_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_8_LC_14_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_8_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33587),
            .lcout(\CONTROL.tempCounterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_0C_net ),
            .ce(N__34954),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_4_LC_14_25_0 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_4_LC_14_25_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_4_LC_14_25_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.tempCounter_4_LC_14_25_0  (
            .in0(N__45262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.tempCounterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_4C_net ),
            .ce(N__34965),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_1_LC_14_25_2 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_1_LC_14_25_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_1_LC_14_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_1_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45188),
            .lcout(\CONTROL.tempCounterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_4C_net ),
            .ce(N__34965),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_7_LC_14_25_3 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_7_LC_14_25_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_7_LC_14_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_7_LC_14_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73348),
            .lcout(\CONTROL.tempCounterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_4C_net ),
            .ce(N__34965),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_12_LC_14_25_6 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_12_LC_14_25_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_12_LC_14_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_12_LC_14_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36778),
            .lcout(\CONTROL.tempCounterZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_4C_net ),
            .ce(N__34965),
            .sr(_gnd_net_));
    defparam \CONTROL.tempCounter_2_LC_14_25_7 .C_ON=1'b0;
    defparam \CONTROL.tempCounter_2_LC_14_25_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.tempCounter_2_LC_14_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.tempCounter_2_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45316),
            .lcout(\CONTROL.tempCounterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.tempCounter_4C_net ),
            .ce(N__34965),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstack_addrstack_0_0_RNO_LC_15_8_0 .C_ON=1'b0;
    defparam \CONTROL.addrstack_addrstack_0_0_RNO_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstack_addrstack_0_0_RNO_LC_15_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \CONTROL.addrstack_addrstack_0_0_RNO_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57751),
            .lcout(\CONTROL.addrstack_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNII2KJ41_4_LC_15_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNII2KJ41_4_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNII2KJ41_4_LC_15_8_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNII2KJ41_4_LC_15_8_2  (
            .in0(N__56415),
            .in1(N__59618),
            .in2(N__59902),
            .in3(N__56266),
            .lcout(\ALU.d_RNII2KJ41Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIR6J013_2_LC_15_8_5 .C_ON=1'b0;
    defparam \ALU.d_RNIR6J013_2_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIR6J013_2_LC_15_8_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \ALU.d_RNIR6J013_2_LC_15_8_5  (
            .in0(N__33744),
            .in1(N__56473),
            .in2(N__68932),
            .in3(N__69977),
            .lcout(\ALU.d_RNIR6J013Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_173_c_RNO_LC_15_8_6 .C_ON=1'b0;
    defparam \ALU.mult_173_c_RNO_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_173_c_RNO_LC_15_8_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.mult_173_c_RNO_LC_15_8_6  (
            .in0(N__59884),
            .in1(N__59619),
            .in2(N__66029),
            .in3(N__66754),
            .lcout(\ALU.mult_173_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI68LSH_9_LC_15_8_7 .C_ON=1'b0;
    defparam \ALU.d_RNI68LSH_9_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI68LSH_9_LC_15_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI68LSH_9_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__62785),
            .in2(_gnd_net_),
            .in3(N__56414),
            .lcout(\ALU.d_RNI68LSHZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_173_c_RNIO8AO16_LC_15_9_0 .C_ON=1'b1;
    defparam \ALU.mult_173_c_RNIO8AO16_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_173_c_RNIO8AO16_LC_15_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ALU.mult_173_c_RNIO8AO16_LC_15_9_0  (
            .in0(N__35236),
            .in1(N__35330),
            .in2(N__33707),
            .in3(_gnd_net_),
            .lcout(\ALU.mult_173_c_RNIO8AOZ0Z16 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\ALU.mult_19_c6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_432_c_RNI5DJ6A3_LC_15_9_1 .C_ON=1'b1;
    defparam \ALU.mult_432_c_RNI5DJ6A3_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_432_c_RNI5DJ6A3_LC_15_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_432_c_RNI5DJ6A3_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__33698),
            .in2(N__33689),
            .in3(N__33680),
            .lcout(\ALU.mult_19_7 ),
            .ltout(),
            .carryin(\ALU.mult_19_c6 ),
            .carryout(\ALU.mult_19_c7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_435_c_RNIOA29R3_LC_15_9_2 .C_ON=1'b1;
    defparam \ALU.mult_435_c_RNIOA29R3_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_435_c_RNIOA29R3_LC_15_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_435_c_RNIOA29R3_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__33677),
            .in2(N__33665),
            .in3(N__33656),
            .lcout(\ALU.mult_19_8 ),
            .ltout(),
            .carryin(\ALU.mult_19_c7 ),
            .carryout(\ALU.mult_19_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_438_c_RNIG9IJJ3_LC_15_9_3 .C_ON=1'b1;
    defparam \ALU.mult_438_c_RNIG9IJJ3_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_438_c_RNIG9IJJ3_LC_15_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_438_c_RNIG9IJJ3_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__33653),
            .in2(N__33644),
            .in3(N__33935),
            .lcout(\ALU.mult_19_9 ),
            .ltout(),
            .carryin(\ALU.mult_19_c8 ),
            .carryout(\ALU.mult_19_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_441_c_RNIE942B3_LC_15_9_4 .C_ON=1'b1;
    defparam \ALU.mult_441_c_RNIE942B3_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_441_c_RNIE942B3_LC_15_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_441_c_RNIE942B3_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__33932),
            .in2(N__33923),
            .in3(N__33914),
            .lcout(\ALU.mult_19_10 ),
            .ltout(),
            .carryin(\ALU.mult_19_c9 ),
            .carryout(\ALU.mult_19_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_444_c_RNIOQ6GB3_LC_15_9_5 .C_ON=1'b1;
    defparam \ALU.mult_444_c_RNIOQ6GB3_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_444_c_RNIOQ6GB3_LC_15_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_444_c_RNIOQ6GB3_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__33911),
            .in2(N__33902),
            .in3(N__33890),
            .lcout(\ALU.mult_19_11 ),
            .ltout(),
            .carryin(\ALU.mult_19_c10 ),
            .carryout(\ALU.mult_19_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_447_c_RNIE3M1A3_LC_15_9_6 .C_ON=1'b1;
    defparam \ALU.mult_447_c_RNIE3M1A3_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_447_c_RNIE3M1A3_LC_15_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_447_c_RNIE3M1A3_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__33887),
            .in2(N__33881),
            .in3(N__33869),
            .lcout(\ALU.mult_19_12 ),
            .ltout(),
            .carryin(\ALU.mult_19_c11 ),
            .carryout(\ALU.mult_19_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_450_c_RNIB3GKA3_LC_15_9_7 .C_ON=1'b1;
    defparam \ALU.mult_450_c_RNIB3GKA3_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_450_c_RNIB3GKA3_LC_15_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_450_c_RNIB3GKA3_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__33866),
            .in2(N__33860),
            .in3(N__33845),
            .lcout(\ALU.mult_19_13 ),
            .ltout(),
            .carryin(\ALU.mult_19_c12 ),
            .carryout(\ALU.mult_19_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_453_c_RNI9IGIB3_LC_15_10_0 .C_ON=1'b1;
    defparam \ALU.mult_453_c_RNI9IGIB3_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_453_c_RNI9IGIB3_LC_15_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_453_c_RNI9IGIB3_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__33842),
            .in2(N__33836),
            .in3(N__33821),
            .lcout(\ALU.mult_19_14 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\ALU.mult_19_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_19_c14_THRU_LUT4_0_LC_15_10_1 .C_ON=1'b0;
    defparam \ALU.mult_19_c14_THRU_LUT4_0_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_19_c14_THRU_LUT4_0_LC_15_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.mult_19_c14_THRU_LUT4_0_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33818),
            .lcout(\ALU.mult_19_c14_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINP3HG_2_LC_15_10_2 .C_ON=1'b0;
    defparam \ALU.d_RNINP3HG_2_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINP3HG_2_LC_15_10_2 .LUT_INIT=16'b0010111000000000;
    LogicCell40 \ALU.d_RNINP3HG_2_LC_15_10_2  (
            .in0(N__39101),
            .in1(N__53290),
            .in2(N__39047),
            .in3(N__66176),
            .lcout(\ALU.mult_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIMNQ8E1_12_LC_15_10_4 .C_ON=1'b0;
    defparam \ALU.c_RNIMNQ8E1_12_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIMNQ8E1_12_LC_15_10_4 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.c_RNIMNQ8E1_12_LC_15_10_4  (
            .in0(N__65936),
            .in1(N__60953),
            .in2(N__61210),
            .in3(N__66753),
            .lcout(\ALU.mult_13_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_486_c_RNIPJD0I5_LC_15_10_6 .C_ON=1'b0;
    defparam \ALU.mult_486_c_RNIPJD0I5_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_486_c_RNIPJD0I5_LC_15_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.mult_486_c_RNIPJD0I5_LC_15_10_6  (
            .in0(N__58987),
            .in1(N__35252),
            .in2(_gnd_net_),
            .in3(N__51334),
            .lcout(),
            .ltout(\ALU.mult_486_c_RNIPJD0IZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_4_c_RNI2R6596_LC_15_10_7 .C_ON=1'b0;
    defparam \ALU.addsub_cry_4_c_RNI2R6596_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_4_c_RNI2R6596_LC_15_10_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.addsub_cry_4_c_RNI2R6596_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__67065),
            .in2(N__34019),
            .in3(N__59369),
            .lcout(\ALU.addsub_cry_4_c_RNI2RZ0Z6596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5S4HI_5_LC_15_11_0 .C_ON=1'b0;
    defparam \ALU.d_RNI5S4HI_5_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5S4HI_5_LC_15_11_0 .LUT_INIT=16'b1011100110010100;
    LogicCell40 \ALU.d_RNI5S4HI_5_LC_15_11_0  (
            .in0(N__34011),
            .in1(N__74882),
            .in2(N__63302),
            .in3(N__59602),
            .lcout(\ALU.log_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICGRJG_1_LC_15_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNICGRJG_1_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICGRJG_1_LC_15_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNICGRJG_1_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__65522),
            .in2(_gnd_net_),
            .in3(N__55953),
            .lcout(\ALU.d_RNICGRJGZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_4_c_RNI5L6IQA_LC_15_11_3 .C_ON=1'b0;
    defparam \ALU.addsub_cry_4_c_RNI5L6IQA_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_4_c_RNI5L6IQA_LC_15_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.addsub_cry_4_c_RNI5L6IQA_LC_15_11_3  (
            .in0(N__34177),
            .in1(N__35594),
            .in2(_gnd_net_),
            .in3(N__33965),
            .lcout(\ALU.addsub_cry_4_c_RNI5L6IQAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBVMTL_5_LC_15_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNIBVMTL_5_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBVMTL_5_LC_15_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIBVMTL_5_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__59601),
            .in2(_gnd_net_),
            .in3(N__68729),
            .lcout(\ALU.d_RNIBVMTLZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7ATTC1_8_LC_15_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNI7ATTC1_8_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7ATTC1_8_LC_15_11_5 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.d_RNI7ATTC1_8_LC_15_11_5  (
            .in0(N__65717),
            .in1(N__62820),
            .in2(N__62000),
            .in3(N__66629),
            .lcout(\ALU.mult_9_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVMDLO_5_LC_15_11_6 .C_ON=1'b0;
    defparam \ALU.d_RNIVMDLO_5_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVMDLO_5_LC_15_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIVMDLO_5_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__59600),
            .in2(_gnd_net_),
            .in3(N__65716),
            .lcout(\ALU.d_RNIVMDLOZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9QA4D1_1_0_LC_15_11_7 .C_ON=1'b0;
    defparam \ALU.d_RNI9QA4D1_1_0_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9QA4D1_1_0_LC_15_11_7 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \ALU.d_RNI9QA4D1_1_0_LC_15_11_7  (
            .in0(N__65718),
            .in1(N__60585),
            .in2(N__65564),
            .in3(N__66630),
            .lcout(\ALU.N_806_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNILV28R1_15_LC_15_12_0 .C_ON=1'b0;
    defparam \ALU.c_RNILV28R1_15_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNILV28R1_15_LC_15_12_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ALU.c_RNILV28R1_15_LC_15_12_0  (
            .in0(N__68727),
            .in1(N__65720),
            .in2(N__63670),
            .in3(N__66579),
            .lcout(\ALU.N_1030 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9QA4D1_0_0_LC_15_12_1 .C_ON=1'b0;
    defparam \ALU.d_RNI9QA4D1_0_0_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9QA4D1_0_0_LC_15_12_1 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.d_RNI9QA4D1_0_0_LC_15_12_1  (
            .in0(N__66580),
            .in1(N__60575),
            .in2(N__65827),
            .in3(N__65527),
            .lcout(\ALU.rshift_3_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIF6GEF1_12_LC_15_12_2 .C_ON=1'b0;
    defparam \ALU.c_RNIF6GEF1_12_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIF6GEF1_12_LC_15_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.c_RNIF6GEF1_12_LC_15_12_2  (
            .in0(N__60954),
            .in1(N__68721),
            .in2(N__65928),
            .in3(N__61170),
            .lcout(\ALU.c_RNIF6GEF1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN3QUB1_2_LC_15_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNIN3QUB1_2_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN3QUB1_2_LC_15_12_4 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.d_RNIN3QUB1_2_LC_15_12_4  (
            .in0(N__66175),
            .in1(N__65719),
            .in2(N__60205),
            .in3(N__66577),
            .lcout(\ALU.mult_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISLOMK_1_LC_15_12_5 .C_ON=1'b0;
    defparam \ALU.d_RNISLOMK_1_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISLOMK_1_LC_15_12_5 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \ALU.d_RNISLOMK_1_LC_15_12_5  (
            .in0(N__34095),
            .in1(N__34681),
            .in2(N__53301),
            .in3(N__34066),
            .lcout(\ALU.status_19_0 ),
            .ltout(\ALU.status_19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_95_c_RNO_LC_15_12_6 .C_ON=1'b0;
    defparam \ALU.mult_95_c_RNO_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_95_c_RNO_LC_15_12_6 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \ALU.mult_95_c_RNO_LC_15_12_6  (
            .in0(N__60133),
            .in1(N__66174),
            .in2(N__34049),
            .in3(N__66581),
            .lcout(\ALU.mult_95_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID4IDO_0_LC_15_12_7 .C_ON=1'b0;
    defparam \ALU.d_RNID4IDO_0_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID4IDO_0_LC_15_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNID4IDO_0_LC_15_12_7  (
            .in0(N__66578),
            .in1(N__60574),
            .in2(_gnd_net_),
            .in3(N__65526),
            .lcout(\ALU.N_765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_388_c_RNIBULDP3_LC_15_13_0 .C_ON=1'b0;
    defparam \ALU.mult_388_c_RNIBULDP3_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_388_c_RNIBULDP3_LC_15_13_0 .LUT_INIT=16'b1010001010101110;
    LogicCell40 \ALU.mult_388_c_RNIBULDP3_LC_15_13_0  (
            .in0(N__34034),
            .in1(N__70184),
            .in2(N__59050),
            .in3(N__47936),
            .lcout(\ALU.mult_388_c_RNIBULDPZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_2_c_RNIUFTGN3_LC_15_13_1 .C_ON=1'b0;
    defparam \ALU.addsub_cry_2_c_RNIUFTGN3_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_2_c_RNIUFTGN3_LC_15_13_1 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \ALU.addsub_cry_2_c_RNIUFTGN3_LC_15_13_1  (
            .in0(N__57231),
            .in1(N__59936),
            .in2(N__46508),
            .in3(N__67064),
            .lcout(),
            .ltout(\ALU.addsub_cry_2_c_RNIUFTGNZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_388_c_RNIEAAJH7_LC_15_13_2 .C_ON=1'b0;
    defparam \ALU.mult_388_c_RNIEAAJH7_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_388_c_RNIEAAJH7_LC_15_13_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.mult_388_c_RNIEAAJH7_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__34133),
            .in2(N__34022),
            .in3(N__34253),
            .lcout(\ALU.mult_388_c_RNIEAAJHZ0Z7 ),
            .ltout(\ALU.mult_388_c_RNIEAAJHZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_388_c_RNIPGN6Q7_0_LC_15_13_3 .C_ON=1'b0;
    defparam \ALU.mult_388_c_RNIPGN6Q7_0_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_388_c_RNIPGN6Q7_0_LC_15_13_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ALU.mult_388_c_RNIPGN6Q7_0_LC_15_13_3  (
            .in0(N__34241),
            .in1(N__57384),
            .in2(N__34247),
            .in3(N__69998),
            .lcout(\ALU.mult_388_c_RNIPGN6Q7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_388_c_RNIPGN6Q7_LC_15_13_4 .C_ON=1'b0;
    defparam \ALU.mult_388_c_RNIPGN6Q7_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_388_c_RNIPGN6Q7_LC_15_13_4 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \ALU.mult_388_c_RNIPGN6Q7_LC_15_13_4  (
            .in0(N__69999),
            .in1(N__34242),
            .in2(N__57405),
            .in3(N__34187),
            .lcout(\ALU.mult_388_c_RNIPGN6QZ0Z7 ),
            .ltout(\ALU.mult_388_c_RNIPGN6QZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_3_LC_15_13_5 .C_ON=1'b0;
    defparam \ALU.a_3_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.a_3_LC_15_13_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.a_3_LC_15_13_5  (
            .in0(N__58740),
            .in1(_gnd_net_),
            .in2(N__34181),
            .in3(N__58665),
            .lcout(\ALU.aZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73145),
            .ce(N__71189),
            .sr(_gnd_net_));
    defparam \ALU.a_15_d_s_5_LC_15_13_6 .C_ON=1'b0;
    defparam \ALU.a_15_d_s_5_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_d_s_5_LC_15_13_6 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \ALU.a_15_d_s_5_LC_15_13_6  (
            .in0(N__59009),
            .in1(_gnd_net_),
            .in2(N__67115),
            .in3(N__70186),
            .lcout(\ALU.a_15_d_sZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a32_LC_15_13_7 .C_ON=1'b0;
    defparam \ALU.a32_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.a32_LC_15_13_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ALU.a32_LC_15_13_7  (
            .in0(N__70185),
            .in1(N__67060),
            .in2(_gnd_net_),
            .in3(N__59005),
            .lcout(\ALU.aZ0Z32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_5_c_RNI6ET5D3_LC_15_14_0 .C_ON=1'b0;
    defparam \ALU.mult_5_c_RNI6ET5D3_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_5_c_RNI6ET5D3_LC_15_14_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \ALU.mult_5_c_RNI6ET5D3_LC_15_14_0  (
            .in0(N__70089),
            .in1(N__59001),
            .in2(N__34157),
            .in3(N__34142),
            .lcout(\ALU.mult_5_c_RNI6ET5DZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_d_s_3_LC_15_14_1 .C_ON=1'b0;
    defparam \ALU.a_15_d_s_3_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_d_s_3_LC_15_14_1 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \ALU.a_15_d_s_3_LC_15_14_1  (
            .in0(N__67052),
            .in1(_gnd_net_),
            .in2(N__59049),
            .in3(N__70090),
            .lcout(\ALU.a_15_d_sZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_1_c_RNI8FKPL3_LC_15_14_2 .C_ON=1'b0;
    defparam \ALU.addsub_cry_1_c_RNI8FKPL3_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_1_c_RNI8FKPL3_LC_15_14_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \ALU.addsub_cry_1_c_RNI8FKPL3_LC_15_14_2  (
            .in0(N__57227),
            .in1(N__60290),
            .in2(N__43164),
            .in3(N__67053),
            .lcout(),
            .ltout(\ALU.addsub_cry_1_c_RNI8FKPLZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_1_c_RNIJP8K37_LC_15_14_3 .C_ON=1'b0;
    defparam \ALU.addsub_cry_1_c_RNIJP8K37_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_1_c_RNIJP8K37_LC_15_14_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.addsub_cry_1_c_RNIJP8K37_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__34132),
            .in2(N__34121),
            .in3(N__34118),
            .lcout(\ALU.addsub_cry_1_c_RNIJP8KZ0Z37 ),
            .ltout(\ALU.addsub_cry_1_c_RNIJP8KZ0Z37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_1_c_RNIICPEC7_0_LC_15_14_4 .C_ON=1'b0;
    defparam \ALU.addsub_cry_1_c_RNIICPEC7_0_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_1_c_RNIICPEC7_0_LC_15_14_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ALU.addsub_cry_1_c_RNIICPEC7_0_LC_15_14_4  (
            .in0(N__57372),
            .in1(N__70000),
            .in2(N__34280),
            .in3(N__43574),
            .lcout(\ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_1_c_RNIICPEC7_LC_15_14_5 .C_ON=1'b0;
    defparam \ALU.addsub_cry_1_c_RNIICPEC7_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_1_c_RNIICPEC7_LC_15_14_5 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \ALU.addsub_cry_1_c_RNIICPEC7_LC_15_14_5  (
            .in0(N__43573),
            .in1(N__57371),
            .in2(N__70011),
            .in3(N__34277),
            .lcout(\ALU.addsub_cry_1_c_RNIICPECZ0Z7 ),
            .ltout(\ALU.addsub_cry_1_c_RNIICPECZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_2_LC_15_14_6 .C_ON=1'b0;
    defparam \ALU.a_2_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \ALU.a_2_LC_15_14_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.a_2_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__39603),
            .in2(N__34271),
            .in3(N__39514),
            .lcout(\ALU.aZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73150),
            .ce(N__71213),
            .sr(_gnd_net_));
    defparam \ALU.un1_operation_5_LC_15_14_7 .C_ON=1'b0;
    defparam \ALU.un1_operation_5_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_operation_5_LC_15_14_7 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \ALU.un1_operation_5_LC_15_14_7  (
            .in0(N__67051),
            .in1(_gnd_net_),
            .in2(N__59048),
            .in3(N__70088),
            .lcout(\ALU.un1_operation_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIG7RU_9_LC_15_15_0 .C_ON=1'b0;
    defparam \ALU.e_RNIG7RU_9_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIG7RU_9_LC_15_15_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNIG7RU_9_LC_15_15_0  (
            .in0(N__43553),
            .in1(N__47277),
            .in2(N__46211),
            .in3(N__54284),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI0FTR1_9_LC_15_15_1 .C_ON=1'b0;
    defparam \ALU.c_RNI0FTR1_9_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI0FTR1_9_LC_15_15_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNI0FTR1_9_LC_15_15_1  (
            .in0(N__72353),
            .in1(N__46667),
            .in2(N__34268),
            .in3(N__47194),
            .lcout(\ALU.N_1094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIID111_9_LC_15_15_2 .C_ON=1'b0;
    defparam \ALU.b_RNIID111_9_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIID111_9_LC_15_15_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNIID111_9_LC_15_15_2  (
            .in0(N__48833),
            .in1(N__47276),
            .in2(N__48991),
            .in3(N__54285),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4R9G1_9_LC_15_15_3 .C_ON=1'b0;
    defparam \ALU.d_RNI4R9G1_9_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4R9G1_9_LC_15_15_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNI4R9G1_9_LC_15_15_3  (
            .in0(N__37960),
            .in1(N__52745),
            .in2(N__34265),
            .in3(N__47195),
            .lcout(),
            .ltout(\ALU.N_1142_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7ELL3_9_LC_15_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNI7ELL3_9_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7ELL3_9_LC_15_15_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.d_RNI7ELL3_9_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__34262),
            .in2(N__34256),
            .in3(N__54134),
            .lcout(aluOut_9),
            .ltout(aluOut_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN8NU4_9_LC_15_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNIN8NU4_9_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN8NU4_9_LC_15_15_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.d_RNIN8NU4_9_LC_15_15_5  (
            .in0(N__53231),
            .in1(N__49577),
            .in2(N__34406),
            .in3(N__50153),
            .lcout(\ALU.d_RNIN8NU4Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIVLMT_2_LC_15_16_0 .C_ON=1'b0;
    defparam \ALU.b_RNIVLMT_2_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIVLMT_2_LC_15_16_0 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.b_RNIVLMT_2_LC_15_16_0  (
            .in0(N__36361),
            .in1(N__39415),
            .in2(N__35631),
            .in3(N__36317),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2RL91_2_LC_15_16_1 .C_ON=1'b0;
    defparam \ALU.d_RNI2RL91_2_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2RL91_2_LC_15_16_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNI2RL91_2_LC_15_16_1  (
            .in0(N__34392),
            .in1(N__36073),
            .in2(N__34355),
            .in3(N__54234),
            .lcout(\ALU.N_1135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNITFGR_2_LC_15_16_2 .C_ON=1'b0;
    defparam \ALU.e_RNITFGR_2_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNITFGR_2_LC_15_16_2 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.e_RNITFGR_2_LC_15_16_2  (
            .in0(N__36362),
            .in1(N__34348),
            .in2(N__34333),
            .in3(N__36318),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNITB6K1_2_LC_15_16_3 .C_ON=1'b0;
    defparam \ALU.c_RNITB6K1_2_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNITB6K1_2_LC_15_16_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNITB6K1_2_LC_15_16_3  (
            .in0(N__43896),
            .in1(N__35550),
            .in2(N__34310),
            .in3(N__35872),
            .lcout(),
            .ltout(\ALU.N_1087_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2BA73_2_LC_15_16_4 .C_ON=1'b0;
    defparam \ALU.d_RNI2BA73_2_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2BA73_2_LC_15_16_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNI2BA73_2_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__54112),
            .in2(N__34307),
            .in3(N__34304),
            .lcout(aluOut_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_RNIBQE03_0_0_LC_15_16_5 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_RNIBQE03_0_0_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_ne_RNIBQE03_0_0_LC_15_16_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \CONTROL.operand1_ne_RNIBQE03_0_0_LC_15_16_5  (
            .in0(N__54111),
            .in1(N__50152),
            .in2(N__49578),
            .in3(N__34297),
            .lcout(\CONTROL.operand1_ne_RNIBQE03_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m217_LC_15_17_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m217_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m217_LC_15_17_0 .LUT_INIT=16'b0010100000001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m217_LC_15_17_0  (
            .in0(N__77315),
            .in1(N__75879),
            .in2(N__78863),
            .in3(N__78063),
            .lcout(\PROM.ROMDATA.m217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m238_am_1_LC_15_17_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m238_am_1_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m238_am_1_LC_15_17_1 .LUT_INIT=16'b0000111010100011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m238_am_1_LC_15_17_1  (
            .in0(N__75880),
            .in1(N__78849),
            .in2(N__76634),
            .in3(N__77316),
            .lcout(),
            .ltout(\PROM.ROMDATA.m238_am_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m238_am_LC_15_17_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m238_am_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m238_am_LC_15_17_2 .LUT_INIT=16'b1001011000100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m238_am_LC_15_17_2  (
            .in0(N__78850),
            .in1(N__75881),
            .in2(N__34442),
            .in3(N__78064),
            .lcout(),
            .ltout(\PROM.ROMDATA.m238_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_1_LC_15_17_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_1_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_1_LC_15_17_3 .LUT_INIT=16'b1000110010011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m244_ns_1_LC_15_17_3  (
            .in0(N__72693),
            .in1(N__45092),
            .in2(N__34439),
            .in3(N__45539),
            .lcout(\PROM.ROMDATA.m244_ns_1 ),
            .ltout(\PROM.ROMDATA.m244_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_LC_15_17_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_LC_15_17_4 .LUT_INIT=16'b0001111100001110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m244_ns_LC_15_17_4  (
            .in0(N__72689),
            .in1(N__79420),
            .in2(N__34436),
            .in3(N__54355),
            .lcout(PROM_ROMDATA_dintern_8ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_fast_ne_1_LC_15_17_5 .C_ON=1'b0;
    defparam \CONTROL.operand1_fast_ne_1_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_fast_ne_1_LC_15_17_5 .LUT_INIT=16'b0011001100111010;
    LogicCell40 \CONTROL.operand1_fast_ne_1_LC_15_17_5  (
            .in0(N__54358),
            .in1(N__34428),
            .in2(N__79489),
            .in3(N__72692),
            .lcout(aluOperand1_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_fast_ne_1C_net ),
            .ce(N__36241),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_1_rep1_ne_LC_15_17_6 .C_ON=1'b0;
    defparam \CONTROL.operand1_1_rep1_ne_LC_15_17_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_1_rep1_ne_LC_15_17_6 .LUT_INIT=16'b0001111100001110;
    LogicCell40 \CONTROL.operand1_1_rep1_ne_LC_15_17_6  (
            .in0(N__72690),
            .in1(N__79421),
            .in2(N__34432),
            .in3(N__54356),
            .lcout(aluOperand1_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_fast_ne_1C_net ),
            .ce(N__36241),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_1_rep2_ne_LC_15_17_7 .C_ON=1'b0;
    defparam \CONTROL.operand1_1_rep2_ne_LC_15_17_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_1_rep2_ne_LC_15_17_7 .LUT_INIT=16'b0011001100111010;
    LogicCell40 \CONTROL.operand1_1_rep2_ne_LC_15_17_7  (
            .in0(N__54357),
            .in1(N__34427),
            .in2(N__79488),
            .in3(N__72691),
            .lcout(aluOperand1_1_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_fast_ne_1C_net ),
            .ce(N__36241),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI1OMT_3_LC_15_18_0 .C_ON=1'b0;
    defparam \ALU.b_RNI1OMT_3_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI1OMT_3_LC_15_18_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI1OMT_3_LC_15_18_0  (
            .in0(N__39866),
            .in1(N__36363),
            .in2(N__44242),
            .in3(N__36324),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6VL91_3_LC_15_18_1 .C_ON=1'b0;
    defparam \ALU.d_RNI6VL91_3_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6VL91_3_LC_15_18_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.d_RNI6VL91_3_LC_15_18_1  (
            .in0(N__37850),
            .in1(N__58606),
            .in2(N__34409),
            .in3(N__54249),
            .lcout(\ALU.N_1136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIVHGR_3_LC_15_18_2 .C_ON=1'b0;
    defparam \ALU.e_RNIVHGR_3_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIVHGR_3_LC_15_18_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNIVHGR_3_LC_15_18_2  (
            .in0(N__37822),
            .in1(N__36364),
            .in2(N__37801),
            .in3(N__36325),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI1G6K1_3_LC_15_18_3 .C_ON=1'b0;
    defparam \ALU.c_RNI1G6K1_3_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI1G6K1_3_LC_15_18_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.c_RNI1G6K1_3_LC_15_18_3  (
            .in0(N__37768),
            .in1(N__37741),
            .in2(N__34601),
            .in3(N__43897),
            .lcout(),
            .ltout(\ALU.N_1088_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAJA73_3_LC_15_18_4 .C_ON=1'b0;
    defparam \ALU.d_RNIAJA73_3_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAJA73_3_LC_15_18_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.d_RNIAJA73_3_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__34598),
            .in2(N__34592),
            .in3(N__54041),
            .lcout(aluOut_3),
            .ltout(aluOut_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIH16V3_2_LC_15_18_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIH16V3_2_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIH16V3_2_LC_15_18_5 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \CONTROL.busState_1_RNIH16V3_2_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__49501),
            .in2(N__34589),
            .in3(N__50157),
            .lcout(busState_1_RNIH16V3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI48EA1_13_LC_15_19_0 .C_ON=1'b0;
    defparam \ALU.a_RNI48EA1_13_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI48EA1_13_LC_15_19_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.a_RNI48EA1_13_LC_15_19_0  (
            .in0(N__57166),
            .in1(N__34559),
            .in2(N__52487),
            .in3(N__43919),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIAAVQ1_13_LC_15_19_1 .C_ON=1'b0;
    defparam \ALU.c_RNIAAVQ1_13_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIAAVQ1_13_LC_15_19_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNIAAVQ1_13_LC_15_19_1  (
            .in0(N__52358),
            .in1(N__67352),
            .in2(N__34571),
            .in3(N__47201),
            .lcout(\ALU.N_1098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI6GQI1_13_LC_15_19_2 .C_ON=1'b0;
    defparam \ALU.b_RNI6GQI1_13_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI6GQI1_13_LC_15_19_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI6GQI1_13_LC_15_19_2  (
            .in0(N__51548),
            .in1(N__34558),
            .in2(N__57638),
            .in3(N__43918),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEQNB2_13_LC_15_19_3 .C_ON=1'b0;
    defparam \ALU.d_RNIEQNB2_13_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEQNB2_13_LC_15_19_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIEQNB2_13_LC_15_19_3  (
            .in0(N__57892),
            .in1(N__65056),
            .in2(N__34511),
            .in3(N__47202),
            .lcout(),
            .ltout(\ALU.N_1146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIR85G4_13_LC_15_19_4 .C_ON=1'b0;
    defparam \ALU.c_RNIR85G4_13_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIR85G4_13_LC_15_19_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.c_RNIR85G4_13_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__34508),
            .in2(N__34502),
            .in3(N__54059),
            .lcout(aluOut_13),
            .ltout(aluOut_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIKLFS7_0_LC_15_19_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIKLFS7_0_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIKLFS7_0_LC_15_19_5 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \CONTROL.busState_1_RNIKLFS7_0_LC_15_19_5  (
            .in0(N__34499),
            .in1(N__34490),
            .in2(N__34460),
            .in3(N__49806),
            .lcout(\CONTROL.bus_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI4KP71_1_LC_15_20_0 .C_ON=1'b0;
    defparam \ALU.b_RNI4KP71_1_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI4KP71_1_LC_15_20_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI4KP71_1_LC_15_20_0  (
            .in0(N__48409),
            .in1(N__46925),
            .in2(N__49177),
            .in3(N__46812),
            .lcout(\ALU.operand2_6_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJMOB4_0_1_LC_15_20_1 .C_ON=1'b0;
    defparam \ALU.c_RNIJMOB4_0_1_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJMOB4_0_1_LC_15_20_1 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \ALU.c_RNIJMOB4_0_1_LC_15_20_1  (
            .in0(N__53964),
            .in1(N__34652),
            .in2(N__71435),
            .in3(N__34645),
            .lcout(),
            .ltout(\ALU.c_RNIJMOB4_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID42JA_1_LC_15_20_2 .C_ON=1'b0;
    defparam \ALU.d_RNID42JA_1_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID42JA_1_LC_15_20_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNID42JA_1_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__34661),
            .in2(N__34688),
            .in3(N__34634),
            .lcout(\ALU.d_RNID42JAZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7NGR1_1_LC_15_20_3 .C_ON=1'b0;
    defparam \ALU.d_RNI7NGR1_1_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7NGR1_1_LC_15_20_3 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \ALU.d_RNI7NGR1_1_LC_15_20_3  (
            .in0(N__46815),
            .in1(N__52166),
            .in2(N__37516),
            .in3(N__34667),
            .lcout(\ALU.N_1246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI2EJ51_1_LC_15_20_4 .C_ON=1'b0;
    defparam \ALU.e_RNI2EJ51_1_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI2EJ51_1_LC_15_20_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNI2EJ51_1_LC_15_20_4  (
            .in0(N__37238),
            .in1(N__46926),
            .in2(N__46358),
            .in3(N__46813),
            .lcout(),
            .ltout(\ALU.operand2_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3B472_1_LC_15_20_5 .C_ON=1'b0;
    defparam \ALU.c_RNI3B472_1_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3B472_1_LC_15_20_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNI3B472_1_LC_15_20_5  (
            .in0(N__46814),
            .in1(N__48943),
            .in2(N__34655),
            .in3(N__46463),
            .lcout(\ALU.N_1198 ),
            .ltout(\ALU.N_1198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJMOB4_1_LC_15_20_6 .C_ON=1'b0;
    defparam \ALU.c_RNIJMOB4_1_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJMOB4_1_LC_15_20_6 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \ALU.c_RNIJMOB4_1_LC_15_20_6  (
            .in0(N__34646),
            .in1(N__71380),
            .in2(N__34637),
            .in3(N__53963),
            .lcout(\ALU.c_RNIJMOB4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI7FBMHV_7_LC_15_21_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI7FBMHV_7_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI7FBMHV_7_LC_15_21_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI7FBMHV_7_LC_15_21_0  (
            .in0(N__34628),
            .in1(N__34856),
            .in2(N__36263),
            .in3(N__34823),
            .lcout(\CONTROL.N_5 ),
            .ltout(\CONTROL.N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNIPON8992_3_LC_15_21_1 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNIPON8992_3_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNIPON8992_3_LC_15_21_1 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \CONTROL.addrstackptr_RNIPON8992_3_LC_15_21_1  (
            .in0(N__34807),
            .in1(N__34739),
            .in2(N__34622),
            .in3(N__34816),
            .lcout(\CONTROL.addrstackptr_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI0GOJ_2_LC_15_21_2 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI0GOJ_2_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI0GOJ_2_LC_15_21_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNI0GOJ_2_LC_15_21_2  (
            .in0(N__34847),
            .in1(N__54814),
            .in2(_gnd_net_),
            .in3(N__49948),
            .lcout(\CONTROL.N_163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI060HM91_2_LC_15_21_3 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI060HM91_2_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI060HM91_2_LC_15_21_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI060HM91_2_LC_15_21_3  (
            .in0(N__38437),
            .in1(N__57792),
            .in2(N__60743),
            .in3(N__41923),
            .lcout(\CONTROL.un1_addrstackptr_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_2_7_LC_15_21_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_2_7_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_2_7_LC_15_21_4 .LUT_INIT=16'b1011101010111111;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIO2O5VB_2_7_LC_15_21_4  (
            .in0(N__41489),
            .in1(N__54661),
            .in2(N__71852),
            .in3(N__44712),
            .lcout(\CONTROL.g0_3_i_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_3_LC_15_21_6 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_3_LC_15_21_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_3_LC_15_21_6 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \CONTROL.addrstackptr_3_LC_15_21_6  (
            .in0(N__34817),
            .in1(N__34808),
            .in2(N__34753),
            .in3(N__34778),
            .lcout(\CONTROL.addrstackptrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.addrstackptr_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_ne_1_LC_15_22_0 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_ne_1_LC_15_22_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_ne_1_LC_15_22_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \CONTROL.aluOperation_ne_1_LC_15_22_0  (
            .in0(N__42196),
            .in1(N__71831),
            .in2(N__72305),
            .in3(N__54587),
            .lcout(aluOperation_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluOperation_ne_1C_net ),
            .ce(N__38125),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState101_3_0_a2_308_LC_15_22_1 .C_ON=1'b0;
    defparam \CONTROL.un1_busState101_3_0_a2_308_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState101_3_0_a2_308_LC_15_22_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \CONTROL.un1_busState101_3_0_a2_308_LC_15_22_1  (
            .in0(N__72297),
            .in1(N__71830),
            .in2(_gnd_net_),
            .in3(N__42195),
            .lcout(\CONTROL.N_83_0 ),
            .ltout(\CONTROL.N_83_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_4_LC_15_22_2 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_4_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_4_LC_15_22_2 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \CONTROL.busState_cnst_2_0__m28_0_120_i_i_4_LC_15_22_2  (
            .in0(N__41258),
            .in1(N__34883),
            .in2(N__34715),
            .in3(N__34706),
            .lcout(\CONTROL.m28_0_120_i_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_12_i_o2_6_LC_15_22_3 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_12_i_o2_6_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_12_i_o2_6_LC_15_22_3 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \CONTROL.aluOperation_12_i_o2_6_LC_15_22_3  (
            .in0(N__40958),
            .in1(N__41602),
            .in2(_gnd_net_),
            .in3(N__41257),
            .lcout(\CONTROL.N_75_0 ),
            .ltout(\CONTROL.N_75_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m38_i_2_LC_15_22_4 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m38_i_2_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m38_i_2_LC_15_22_4 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \CONTROL.busState_cnst_2_0__m38_i_2_LC_15_22_4  (
            .in0(N__41603),
            .in1(N__36797),
            .in2(N__34700),
            .in3(N__44749),
            .lcout(\CONTROL.m38_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_3_LC_15_22_5 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_3_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_3_LC_15_22_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_3_LC_15_22_5  (
            .in0(N__44748),
            .in1(N__44663),
            .in2(N__41696),
            .in3(N__44840),
            .lcout(\CONTROL.N_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState103_0_a2_2_LC_15_22_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState103_0_a2_2_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState103_0_a2_2_LC_15_22_6 .LUT_INIT=16'b0101010101011111;
    LogicCell40 \CONTROL.un1_busState103_0_a2_2_LC_15_22_6  (
            .in0(N__72264),
            .in1(_gnd_net_),
            .in2(N__42220),
            .in3(N__55444),
            .lcout(\CONTROL.N_219 ),
            .ltout(\CONTROL.N_219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_1_0_LC_15_22_7 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_1_0_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_1_0_LC_15_22_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \CONTROL.busState_cnst_2_0__m11_0_a2_1_0_LC_15_22_7  (
            .in0(N__54586),
            .in1(N__44662),
            .in2(N__34877),
            .in3(N__44839),
            .lcout(\CONTROL.N_350_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_1_LC_15_23_0 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_1_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_1_LC_15_23_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \CONTROL.busState_cnst_2_0__m38_i_a2_1_LC_15_23_0  (
            .in0(N__41650),
            .in1(N__38579),
            .in2(_gnd_net_),
            .in3(N__72293),
            .lcout(\CONTROL.N_246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_2_LC_15_23_1 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_2_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m11_0_a2_2_LC_15_23_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \CONTROL.busState_cnst_2_0__m11_0_a2_2_LC_15_23_1  (
            .in0(N__54656),
            .in1(N__44866),
            .in2(N__44759),
            .in3(N__44703),
            .lcout(\CONTROL.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_0_0_LC_15_23_2 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_0_0_LC_15_23_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_0_0_LC_15_23_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_0_0_LC_15_23_2  (
            .in0(N__41651),
            .in1(N__38580),
            .in2(_gnd_net_),
            .in3(N__55466),
            .lcout(),
            .ltout(\CONTROL.m28_0_120_i_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNO_1_1_LC_15_23_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNO_1_1_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNO_1_1_LC_15_23_3 .LUT_INIT=16'b0011001100000011;
    LogicCell40 \CONTROL.busState_1_RNO_1_1_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__38606),
            .in2(N__34874),
            .in3(N__54707),
            .lcout(),
            .ltout(\CONTROL.busState_1_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNO_0_1_LC_15_23_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNO_0_1_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNO_0_1_LC_15_23_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \CONTROL.busState_1_RNO_0_1_LC_15_23_4  (
            .in0(N__38624),
            .in1(_gnd_net_),
            .in2(N__34871),
            .in3(N__38633),
            .lcout(\CONTROL.busState_1_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_7_LC_15_23_5 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_7_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_7_LC_15_23_5 .LUT_INIT=16'b1101111101111111;
    LogicCell40 \CONTROL.g0_3_i_7_LC_15_23_5  (
            .in0(N__55465),
            .in1(N__42216),
            .in2(N__72317),
            .in3(N__54654),
            .lcout(\CONTROL.g0_3_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramWrite_5_m9_0_a2_LC_15_23_6 .C_ON=1'b0;
    defparam \CONTROL.ramWrite_5_m9_0_a2_LC_15_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.ramWrite_5_m9_0_a2_LC_15_23_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \CONTROL.ramWrite_5_m9_0_a2_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__38581),
            .in2(_gnd_net_),
            .in3(N__35182),
            .lcout(\CONTROL.N_345 ),
            .ltout(\CONTROL.N_345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramWrite_LC_15_23_7 .C_ON=1'b0;
    defparam \CONTROL.ramWrite_LC_15_23_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramWrite_LC_15_23_7 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \CONTROL.ramWrite_LC_15_23_7  (
            .in0(N__35156),
            .in1(N__35134),
            .in2(N__35120),
            .in3(N__36817),
            .lcout(ramWrite),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramWriteC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState114_1_0_LC_15_24_0 .C_ON=1'b0;
    defparam \CONTROL.un1_busState114_1_0_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState114_1_0_LC_15_24_0 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \CONTROL.un1_busState114_1_0_LC_15_24_0  (
            .in0(N__54653),
            .in1(N__47043),
            .in2(N__36833),
            .in3(N__47015),
            .lcout(\CONTROL.un1_busState114_1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_12_i_a2_6_LC_15_24_1 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_12_i_a2_6_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_12_i_a2_6_LC_15_24_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \CONTROL.aluOperation_12_i_a2_6_LC_15_24_1  (
            .in0(N__44882),
            .in1(N__54652),
            .in2(N__41433),
            .in3(N__44700),
            .lcout(\CONTROL.N_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_10_LC_15_24_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_10_LC_15_24_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_10_LC_15_24_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_19_10_LC_15_24_2  (
            .in0(N__34919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.dout_reto_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73233),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m1_LC_15_24_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m1_LC_15_24_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m1_LC_15_24_3 .LUT_INIT=16'b0000000000110101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m1_LC_15_24_3  (
            .in0(N__64747),
            .in1(N__64711),
            .in2(N__73661),
            .in3(N__77282),
            .lcout(\PROM.ROMDATA.m1 ),
            .ltout(\PROM.ROMDATA.m1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m312_am_LC_15_24_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m312_am_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m312_am_LC_15_24_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m312_am_LC_15_24_4  (
            .in0(N__78855),
            .in1(N__73857),
            .in2(N__34886),
            .in3(N__75906),
            .lcout(\PROM.ROMDATA.m312_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m298_am_LC_15_24_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m298_am_LC_15_24_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m298_am_LC_15_24_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m298_am_LC_15_24_5  (
            .in0(N__75905),
            .in1(N__64877),
            .in2(N__73873),
            .in3(N__78856),
            .lcout(\PROM.ROMDATA.m298_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m2_LC_15_24_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m2_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m2_LC_15_24_6 .LUT_INIT=16'b0000101000100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m2_LC_15_24_6  (
            .in0(N__77283),
            .in1(N__64748),
            .in2(N__64715),
            .in3(N__73627),
            .lcout(\PROM.ROMDATA.m2 ),
            .ltout(\PROM.ROMDATA.m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m451_am_LC_15_24_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m451_am_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m451_am_LC_15_24_7 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m451_am_LC_15_24_7  (
            .in0(N__75904),
            .in1(N__78996),
            .in2(N__35333),
            .in3(N__78854),
            .lcout(\PROM.ROMDATA.m451_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0OE8H_6_LC_16_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNI0OE8H_6_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0OE8H_6_LC_16_8_1 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \ALU.d_RNI0OE8H_6_LC_16_8_1  (
            .in0(N__39086),
            .in1(N__62571),
            .in2(N__39044),
            .in3(N__53302),
            .lcout(\ALU.mult_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIG7E8H_4_LC_16_8_3 .C_ON=1'b0;
    defparam \ALU.d_RNIG7E8H_4_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIG7E8H_4_LC_16_8_3 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \ALU.d_RNIG7E8H_4_LC_16_8_3  (
            .in0(N__39087),
            .in1(N__59898),
            .in2(N__39045),
            .in3(N__53303),
            .lcout(\ALU.mult_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_18_cry_0_c_RNO_LC_16_8_5 .C_ON=1'b0;
    defparam \ALU.status_18_cry_0_c_RNO_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_18_cry_0_c_RNO_LC_16_8_5 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \ALU.status_18_cry_0_c_RNO_LC_16_8_5  (
            .in0(N__39088),
            .in1(N__60624),
            .in2(N__39046),
            .in3(N__53304),
            .lcout(\ALU.status_18_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIDBF7E1_14_LC_16_8_6 .C_ON=1'b0;
    defparam \ALU.c_RNIDBF7E1_14_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIDBF7E1_14_LC_16_8_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.c_RNIDBF7E1_14_LC_16_8_6  (
            .in0(N__60994),
            .in1(N__65989),
            .in2(N__63854),
            .in3(N__66715),
            .lcout(\ALU.lshift_3_ns_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_391_c_RNIEC73T4_LC_16_9_0 .C_ON=1'b1;
    defparam \ALU.mult_391_c_RNIEC73T4_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_391_c_RNIEC73T4_LC_16_9_0 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \ALU.mult_391_c_RNIEC73T4_LC_16_9_0  (
            .in0(N__59124),
            .in1(N__35306),
            .in2(N__35297),
            .in3(N__51491),
            .lcout(\ALU.mult_391_c_RNIEC73TZ0Z4 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\ALU.mult_25_c4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_486_c_RNINTF5V4_LC_16_9_1 .C_ON=1'b1;
    defparam \ALU.mult_486_c_RNINTF5V4_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_486_c_RNINTF5V4_LC_16_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_486_c_RNINTF5V4_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__36986),
            .in2(N__35267),
            .in3(N__35246),
            .lcout(\ALU.mult_5 ),
            .ltout(),
            .carryin(\ALU.mult_25_c4 ),
            .carryout(\ALU.mult_25_c5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_489_c_RNIPFFTA9_LC_16_9_2 .C_ON=1'b1;
    defparam \ALU.mult_489_c_RNIPFFTA9_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_489_c_RNIPFFTA9_LC_16_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_489_c_RNIPFFTA9_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__35243),
            .in2(N__35237),
            .in3(N__35216),
            .lcout(\ALU.mult_6 ),
            .ltout(),
            .carryin(\ALU.mult_25_c5 ),
            .carryout(\ALU.mult_25_c6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_492_c_RNION7CK6_LC_16_9_3 .C_ON=1'b1;
    defparam \ALU.mult_492_c_RNION7CK6_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_492_c_RNION7CK6_LC_16_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_492_c_RNION7CK6_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__35213),
            .in2(N__35207),
            .in3(N__35192),
            .lcout(\ALU.mult_7 ),
            .ltout(),
            .carryin(\ALU.mult_25_c6 ),
            .carryout(\ALU.mult_25_c7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_495_c_RNI449047_LC_16_9_4 .C_ON=1'b1;
    defparam \ALU.mult_495_c_RNI449047_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_495_c_RNI449047_LC_16_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_495_c_RNI449047_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__35516),
            .in2(N__35504),
            .in3(N__35495),
            .lcout(\ALU.mult_25_8 ),
            .ltout(),
            .carryin(\ALU.mult_25_c7 ),
            .carryout(\ALU.mult_25_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_498_c_RNI5QTSS6_LC_16_9_5 .C_ON=1'b1;
    defparam \ALU.mult_498_c_RNI5QTSS6_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_498_c_RNI5QTSS6_LC_16_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_498_c_RNI5QTSS6_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__35492),
            .in2(N__35480),
            .in3(N__35471),
            .lcout(\ALU.mult_25_9 ),
            .ltout(),
            .carryin(\ALU.mult_25_c8 ),
            .carryout(\ALU.mult_25_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_501_c_RNII3J3L6_LC_16_9_6 .C_ON=1'b1;
    defparam \ALU.mult_501_c_RNII3J3L6_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_501_c_RNII3J3L6_LC_16_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_501_c_RNII3J3L6_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__35468),
            .in2(N__35462),
            .in3(N__35447),
            .lcout(\ALU.mult_25_10 ),
            .ltout(),
            .carryin(\ALU.mult_25_c9 ),
            .carryout(\ALU.mult_25_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_504_c_RNIA6C9P6_LC_16_9_7 .C_ON=1'b1;
    defparam \ALU.mult_504_c_RNIA6C9P6_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_504_c_RNIA6C9P6_LC_16_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_504_c_RNIA6C9P6_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__35444),
            .in2(N__35432),
            .in3(N__35423),
            .lcout(\ALU.mult_25_11 ),
            .ltout(),
            .carryin(\ALU.mult_25_c10 ),
            .carryout(\ALU.mult_25_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_507_c_RNIBABOO6_LC_16_10_0 .C_ON=1'b1;
    defparam \ALU.mult_507_c_RNIBABOO6_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_507_c_RNIBABOO6_LC_16_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_507_c_RNIBABOO6_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__35420),
            .in2(N__35408),
            .in3(N__35399),
            .lcout(\ALU.mult_25_12 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\ALU.mult_25_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_510_c_RNIHTE1V6_LC_16_10_1 .C_ON=1'b1;
    defparam \ALU.mult_510_c_RNIHTE1V6_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_510_c_RNIHTE1V6_LC_16_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_510_c_RNIHTE1V6_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__35396),
            .in2(N__35384),
            .in3(N__35375),
            .lcout(\ALU.mult_25_13 ),
            .ltout(),
            .carryin(\ALU.mult_25_c12 ),
            .carryout(\ALU.mult_25_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_513_c_RNIGEHOR6_LC_16_10_2 .C_ON=1'b1;
    defparam \ALU.mult_513_c_RNIGEHOR6_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_513_c_RNIGEHOR6_LC_16_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_513_c_RNIGEHOR6_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__35372),
            .in2(N__35360),
            .in3(N__35351),
            .lcout(\ALU.mult_25_14 ),
            .ltout(),
            .carryin(\ALU.mult_25_c13 ),
            .carryout(\ALU.mult_25_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_516_c_RNI98SKDC_LC_16_10_3 .C_ON=1'b0;
    defparam \ALU.mult_516_c_RNI98SKDC_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_516_c_RNI98SKDC_LC_16_10_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_516_c_RNI98SKDC_LC_16_10_3  (
            .in0(N__42347),
            .in1(N__35348),
            .in2(N__38894),
            .in3(N__35336),
            .lcout(\ALU.mult_516_c_RNI98SKDCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDR5C61_8_LC_16_10_5 .C_ON=1'b0;
    defparam \ALU.d_RNIDR5C61_8_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDR5C61_8_LC_16_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIDR5C61_8_LC_16_10_5  (
            .in0(N__62859),
            .in1(N__68315),
            .in2(N__68908),
            .in3(N__61983),
            .lcout(\ALU.d_RNIDR5C61Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIUT8OG4_0_LC_16_11_0 .C_ON=1'b0;
    defparam \ALU.d_RNIUT8OG4_0_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIUT8OG4_0_LC_16_11_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.d_RNIUT8OG4_0_LC_16_11_0  (
            .in0(N__68845),
            .in1(N__48082),
            .in2(N__68460),
            .in3(N__48023),
            .lcout(\ALU.d_RNIUT8OG4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI8FSDB2_12_LC_16_11_1 .C_ON=1'b0;
    defparam \ALU.c_RNI8FSDB2_12_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI8FSDB2_12_LC_16_11_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.c_RNI8FSDB2_12_LC_16_11_1  (
            .in0(N__65755),
            .in1(N__61157),
            .in2(N__35588),
            .in3(N__61425),
            .lcout(),
            .ltout(\ALU.N_646_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIMNASS6_12_LC_16_11_2 .C_ON=1'b0;
    defparam \ALU.c_RNIMNASS6_12_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIMNASS6_12_LC_16_11_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.c_RNIMNASS6_12_LC_16_11_2  (
            .in0(N__68846),
            .in1(N__68468),
            .in2(N__35576),
            .in3(N__39175),
            .lcout(),
            .ltout(\ALU.lshift_15_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNICF0UCB_12_LC_16_11_3 .C_ON=1'b0;
    defparam \ALU.c_RNICF0UCB_12_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNICF0UCB_12_LC_16_11_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.c_RNICF0UCB_12_LC_16_11_3  (
            .in0(N__43166),
            .in1(N__43603),
            .in2(N__35573),
            .in3(N__68378),
            .lcout(\ALU.lshift_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINUT6P_13_LC_16_11_4 .C_ON=1'b0;
    defparam \ALU.c_RNINUT6P_13_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINUT6P_13_LC_16_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.c_RNINUT6P_13_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__60938),
            .in2(_gnd_net_),
            .in3(N__65754),
            .lcout(\ALU.c_RNINUT6PZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_365_c_RNO_LC_16_11_6 .C_ON=1'b0;
    defparam \ALU.mult_365_c_RNO_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_365_c_RNO_LC_16_11_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_365_c_RNO_LC_16_11_6  (
            .in0(N__61156),
            .in1(N__65753),
            .in2(N__66717),
            .in3(N__60940),
            .lcout(\ALU.mult_365_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIS83N71_12_LC_16_11_7 .C_ON=1'b0;
    defparam \ALU.c_RNIS83N71_12_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIS83N71_12_LC_16_11_7 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.c_RNIS83N71_12_LC_16_11_7  (
            .in0(N__60939),
            .in1(N__68374),
            .in2(N__61194),
            .in3(N__68844),
            .lcout(\ALU.c_RNIS83N71Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_2_LC_16_12_0 .C_ON=1'b0;
    defparam \ALU.g_2_LC_16_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.g_2_LC_16_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.g_2_LC_16_12_0  (
            .in0(N__39605),
            .in1(N__39531),
            .in2(_gnd_net_),
            .in3(N__39475),
            .lcout(g_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73140),
            .ce(N__70994),
            .sr(_gnd_net_));
    defparam \ALU.g_4_LC_16_12_1 .C_ON=1'b0;
    defparam \ALU.g_4_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.g_4_LC_16_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_4_LC_16_12_1  (
            .in0(N__57382),
            .in1(N__42536),
            .in2(_gnd_net_),
            .in3(N__39394),
            .lcout(g_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73140),
            .ce(N__70994),
            .sr(_gnd_net_));
    defparam \ALU.g_5_LC_16_12_2 .C_ON=1'b0;
    defparam \ALU.g_5_LC_16_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.g_5_LC_16_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_5_LC_16_12_2  (
            .in0(N__57378),
            .in1(N__52628),
            .in2(_gnd_net_),
            .in3(N__39301),
            .lcout(g_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73140),
            .ce(N__70994),
            .sr(_gnd_net_));
    defparam \ALU.g_6_LC_16_12_3 .C_ON=1'b0;
    defparam \ALU.g_6_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.g_6_LC_16_12_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_6_LC_16_12_3  (
            .in0(N__43066),
            .in1(N__43120),
            .in2(_gnd_net_),
            .in3(N__42992),
            .lcout(g_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73140),
            .ce(N__70994),
            .sr(_gnd_net_));
    defparam \ALU.g_3_LC_16_12_4 .C_ON=1'b0;
    defparam \ALU.g_3_LC_16_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.g_3_LC_16_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.g_3_LC_16_12_4  (
            .in0(N__58679),
            .in1(N__58717),
            .in2(_gnd_net_),
            .in3(N__58816),
            .lcout(g_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73140),
            .ce(N__70994),
            .sr(_gnd_net_));
    defparam \ALU.g_10_LC_16_12_5 .C_ON=1'b0;
    defparam \ALU.g_10_LC_16_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.g_10_LC_16_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_10_LC_16_12_5  (
            .in0(N__58526),
            .in1(N__58370),
            .in2(_gnd_net_),
            .in3(N__58284),
            .lcout(g_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73140),
            .ce(N__70994),
            .sr(_gnd_net_));
    defparam \ALU.g_11_LC_16_12_6 .C_ON=1'b0;
    defparam \ALU.g_11_LC_16_12_6 .SEQ_MODE=4'b1000;
    defparam \ALU.g_11_LC_16_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.g_11_LC_16_12_6  (
            .in0(N__58196),
            .in1(N__58110),
            .in2(_gnd_net_),
            .in3(N__58052),
            .lcout(g_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73140),
            .ce(N__70994),
            .sr(_gnd_net_));
    defparam \ALU.f_2_LC_16_13_0 .C_ON=1'b0;
    defparam \ALU.f_2_LC_16_13_0 .SEQ_MODE=4'b1000;
    defparam \ALU.f_2_LC_16_13_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.f_2_LC_16_13_0  (
            .in0(N__39530),
            .in1(N__39607),
            .in2(_gnd_net_),
            .in3(N__39458),
            .lcout(f_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73142),
            .ce(N__67871),
            .sr(_gnd_net_));
    defparam \ALU.f_4_LC_16_13_1 .C_ON=1'b0;
    defparam \ALU.f_4_LC_16_13_1 .SEQ_MODE=4'b1000;
    defparam \ALU.f_4_LC_16_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_4_LC_16_13_1  (
            .in0(N__57389),
            .in1(N__42547),
            .in2(_gnd_net_),
            .in3(N__39387),
            .lcout(f_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73142),
            .ce(N__67871),
            .sr(_gnd_net_));
    defparam \ALU.f_5_LC_16_13_2 .C_ON=1'b0;
    defparam \ALU.f_5_LC_16_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.f_5_LC_16_13_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.f_5_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__57388),
            .in2(N__52636),
            .in3(N__39315),
            .lcout(f_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73142),
            .ce(N__67871),
            .sr(_gnd_net_));
    defparam \ALU.f_6_LC_16_13_3 .C_ON=1'b0;
    defparam \ALU.f_6_LC_16_13_3 .SEQ_MODE=4'b1000;
    defparam \ALU.f_6_LC_16_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_6_LC_16_13_3  (
            .in0(N__43051),
            .in1(N__43119),
            .in2(_gnd_net_),
            .in3(N__42983),
            .lcout(f_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73142),
            .ce(N__67871),
            .sr(_gnd_net_));
    defparam \ALU.f_3_LC_16_13_4 .C_ON=1'b0;
    defparam \ALU.f_3_LC_16_13_4 .SEQ_MODE=4'b1000;
    defparam \ALU.f_3_LC_16_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.f_3_LC_16_13_4  (
            .in0(N__58739),
            .in1(N__58663),
            .in2(_gnd_net_),
            .in3(N__58800),
            .lcout(f_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73142),
            .ce(N__67871),
            .sr(_gnd_net_));
    defparam \ALU.f_10_LC_16_13_5 .C_ON=1'b0;
    defparam \ALU.f_10_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.f_10_LC_16_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_10_LC_16_13_5  (
            .in0(N__58494),
            .in1(N__58366),
            .in2(_gnd_net_),
            .in3(N__58294),
            .lcout(f_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73142),
            .ce(N__67871),
            .sr(_gnd_net_));
    defparam \ALU.f_11_LC_16_13_6 .C_ON=1'b0;
    defparam \ALU.f_11_LC_16_13_6 .SEQ_MODE=4'b1000;
    defparam \ALU.f_11_LC_16_13_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.f_11_LC_16_13_6  (
            .in0(N__58118),
            .in1(N__58188),
            .in2(_gnd_net_),
            .in3(N__58049),
            .lcout(f_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73142),
            .ce(N__67871),
            .sr(_gnd_net_));
    defparam CONSTANT_ZERO_LUT4_LC_16_13_7.C_ON=1'b0;
    defparam CONSTANT_ZERO_LUT4_LC_16_13_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ZERO_LUT4_LC_16_13_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 CONSTANT_ZERO_LUT4_LC_16_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ZERO_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_2_LC_16_14_0 .C_ON=1'b0;
    defparam \ALU.c_2_LC_16_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.c_2_LC_16_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.c_2_LC_16_14_0  (
            .in0(N__39515),
            .in1(N__39599),
            .in2(_gnd_net_),
            .in3(N__39455),
            .lcout(\ALU.cZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73144),
            .ce(N__71554),
            .sr(_gnd_net_));
    defparam \ALU.c_4_LC_16_14_1 .C_ON=1'b0;
    defparam \ALU.c_4_LC_16_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.c_4_LC_16_14_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ALU.c_4_LC_16_14_1  (
            .in0(N__42546),
            .in1(_gnd_net_),
            .in2(N__57383),
            .in3(N__39392),
            .lcout(\ALU.cZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73144),
            .ce(N__71554),
            .sr(_gnd_net_));
    defparam \ALU.c_5_LC_16_14_2 .C_ON=1'b0;
    defparam \ALU.c_5_LC_16_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.c_5_LC_16_14_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_5_LC_16_14_2  (
            .in0(N__52612),
            .in1(N__39314),
            .in2(_gnd_net_),
            .in3(N__57351),
            .lcout(\ALU.cZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73144),
            .ce(N__71554),
            .sr(_gnd_net_));
    defparam \ALU.c_6_LC_16_14_3 .C_ON=1'b0;
    defparam \ALU.c_6_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.c_6_LC_16_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_6_LC_16_14_3  (
            .in0(N__43041),
            .in1(N__43105),
            .in2(_gnd_net_),
            .in3(N__42978),
            .lcout(\ALU.cZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73144),
            .ce(N__71554),
            .sr(_gnd_net_));
    defparam \ALU.c_3_LC_16_14_4 .C_ON=1'b0;
    defparam \ALU.c_3_LC_16_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.c_3_LC_16_14_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_3_LC_16_14_4  (
            .in0(N__58741),
            .in1(N__58664),
            .in2(_gnd_net_),
            .in3(N__58801),
            .lcout(\ALU.cZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73144),
            .ce(N__71554),
            .sr(_gnd_net_));
    defparam \ALU.c_10_LC_16_14_5 .C_ON=1'b0;
    defparam \ALU.c_10_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \ALU.c_10_LC_16_14_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_10_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__58495),
            .in2(N__58373),
            .in3(N__58295),
            .lcout(\ALU.cZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73144),
            .ce(N__71554),
            .sr(_gnd_net_));
    defparam \ALU.c_11_LC_16_14_6 .C_ON=1'b0;
    defparam \ALU.c_11_LC_16_14_6 .SEQ_MODE=4'b1000;
    defparam \ALU.c_11_LC_16_14_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.c_11_LC_16_14_6  (
            .in0(N__58109),
            .in1(N__58189),
            .in2(_gnd_net_),
            .in3(N__58051),
            .lcout(\ALU.cZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73144),
            .ce(N__71554),
            .sr(_gnd_net_));
    defparam \ALU.d_2_LC_16_15_0 .C_ON=1'b0;
    defparam \ALU.d_2_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \ALU.d_2_LC_16_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_2_LC_16_15_0  (
            .in0(N__39598),
            .in1(N__39517),
            .in2(_gnd_net_),
            .in3(N__39457),
            .lcout(\ALU.dZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73147),
            .ce(N__70249),
            .sr(_gnd_net_));
    defparam \ALU.d_4_LC_16_15_1 .C_ON=1'b0;
    defparam \ALU.d_4_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \ALU.d_4_LC_16_15_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_4_LC_16_15_1  (
            .in0(N__42548),
            .in1(N__57396),
            .in2(_gnd_net_),
            .in3(N__39393),
            .lcout(\ALU.dZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73147),
            .ce(N__70249),
            .sr(_gnd_net_));
    defparam \ALU.d_5_LC_16_15_2 .C_ON=1'b0;
    defparam \ALU.d_5_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \ALU.d_5_LC_16_15_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ALU.d_5_LC_16_15_2  (
            .in0(N__52623),
            .in1(_gnd_net_),
            .in2(N__57412),
            .in3(N__39321),
            .lcout(\ALU.dZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73147),
            .ce(N__70249),
            .sr(_gnd_net_));
    defparam \ALU.d_6_LC_16_15_3 .C_ON=1'b0;
    defparam \ALU.d_6_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \ALU.d_6_LC_16_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_6_LC_16_15_3  (
            .in0(N__43065),
            .in1(N__43118),
            .in2(_gnd_net_),
            .in3(N__42982),
            .lcout(\ALU.dZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73147),
            .ce(N__70249),
            .sr(_gnd_net_));
    defparam \ALU.d_3_LC_16_15_4 .C_ON=1'b0;
    defparam \ALU.d_3_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \ALU.d_3_LC_16_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_3_LC_16_15_4  (
            .in0(N__58752),
            .in1(N__58808),
            .in2(_gnd_net_),
            .in3(N__58676),
            .lcout(\ALU.dZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73147),
            .ce(N__70249),
            .sr(_gnd_net_));
    defparam \ALU.d_10_LC_16_15_5 .C_ON=1'b0;
    defparam \ALU.d_10_LC_16_15_5 .SEQ_MODE=4'b1000;
    defparam \ALU.d_10_LC_16_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_10_LC_16_15_5  (
            .in0(N__58525),
            .in1(N__58365),
            .in2(_gnd_net_),
            .in3(N__58299),
            .lcout(\ALU.dZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73147),
            .ce(N__70249),
            .sr(_gnd_net_));
    defparam \ALU.d_11_LC_16_15_6 .C_ON=1'b0;
    defparam \ALU.d_11_LC_16_15_6 .SEQ_MODE=4'b1000;
    defparam \ALU.d_11_LC_16_15_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.d_11_LC_16_15_6  (
            .in0(N__58119),
            .in1(N__58190),
            .in2(_gnd_net_),
            .in3(N__58057),
            .lcout(\ALU.dZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73147),
            .ce(N__70249),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_fast_ne_2_LC_16_16_0 .C_ON=1'b0;
    defparam \CONTROL.operand2_fast_ne_2_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_fast_ne_2_LC_16_16_0 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \CONTROL.operand2_fast_ne_2_LC_16_16_0  (
            .in0(N__44497),
            .in1(N__40297),
            .in2(N__40925),
            .in3(N__79507),
            .lcout(aluOperand2_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_fast_ne_2C_net ),
            .ce(N__40647),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_ne_2_LC_16_16_1 .C_ON=1'b0;
    defparam \CONTROL.operand2_ne_2_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_ne_2_LC_16_16_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \CONTROL.operand2_ne_2_LC_16_16_1  (
            .in0(N__40296),
            .in1(N__40920),
            .in2(N__79527),
            .in3(N__44498),
            .lcout(aluOperand2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_fast_ne_2C_net ),
            .ce(N__40647),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6DCT_11_LC_16_16_2 .C_ON=1'b0;
    defparam \ALU.d_RNI6DCT_11_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6DCT_11_LC_16_16_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNI6DCT_11_LC_16_16_2  (
            .in0(N__57997),
            .in1(N__36184),
            .in2(_gnd_net_),
            .in3(N__43237),
            .lcout(\ALU.d_RNI6DCTZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICJCT_14_LC_16_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNICJCT_14_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICJCT_14_LC_16_16_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNICJCT_14_LC_16_16_3  (
            .in0(N__43238),
            .in1(N__57852),
            .in2(_gnd_net_),
            .in3(N__67783),
            .lcout(\ALU.d_RNICJCTZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_ne_0_LC_16_16_4 .C_ON=1'b0;
    defparam \CONTROL.operand2_ne_0_LC_16_16_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_ne_0_LC_16_16_4 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \CONTROL.operand2_ne_0_LC_16_16_4  (
            .in0(N__72694),
            .in1(N__44927),
            .in2(N__41072),
            .in3(N__50720),
            .lcout(aluOperand2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_fast_ne_2C_net ),
            .ce(N__40647),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI02EVNB_4_LC_16_16_6 .C_ON=1'b0;
    defparam \ALU.d_RNI02EVNB_4_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI02EVNB_4_LC_16_16_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNI02EVNB_4_LC_16_16_6  (
            .in0(N__36158),
            .in1(N__39251),
            .in2(_gnd_net_),
            .in3(N__68516),
            .lcout(\ALU.d_RNI02EVNBZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIG2L52_15_LC_16_17_0 .C_ON=1'b0;
    defparam \ALU.c_RNIG2L52_15_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIG2L52_15_LC_16_17_0 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \ALU.c_RNIG2L52_15_LC_16_17_0  (
            .in0(N__46684),
            .in1(N__36146),
            .in2(N__50404),
            .in3(N__53425),
            .lcout(\ALU.N_1212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI7F2G1_15_LC_16_17_1 .C_ON=1'b0;
    defparam \ALU.a_RNI7F2G1_15_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI7F2G1_15_LC_16_17_1 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.a_RNI7F2G1_15_LC_16_17_1  (
            .in0(N__46549),
            .in1(N__53574),
            .in2(N__46237),
            .in3(N__53477),
            .lcout(\ALU.operand2_3_ns_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI5PJ21_15_LC_16_17_2 .C_ON=1'b0;
    defparam \ALU.a_RNI5PJ21_15_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI5PJ21_15_LC_16_17_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.a_RNI5PJ21_15_LC_16_17_2  (
            .in0(N__46550),
            .in1(N__36371),
            .in2(N__46238),
            .in3(N__36326),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNID2PE1_15_LC_16_17_3 .C_ON=1'b0;
    defparam \ALU.c_RNID2PE1_15_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNID2PE1_15_LC_16_17_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNID2PE1_15_LC_16_17_3  (
            .in0(N__43903),
            .in1(N__50400),
            .in2(N__36140),
            .in3(N__46685),
            .lcout(\ALU.N_1100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI710B1_15_LC_16_17_4 .C_ON=1'b0;
    defparam \ALU.b_RNI710B1_15_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI710B1_15_LC_16_17_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI710B1_15_LC_16_17_4  (
            .in0(N__53612),
            .in1(N__36370),
            .in2(N__53530),
            .in3(N__36327),
            .lcout(\ALU.dout_6_ns_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIE4B6N4_15_LC_16_17_5 .C_ON=1'b0;
    defparam \ALU.c_RNIE4B6N4_15_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIE4B6N4_15_LC_16_17_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ALU.c_RNIE4B6N4_15_LC_16_17_5  (
            .in0(N__37637),
            .in1(N__63615),
            .in2(N__69168),
            .in3(N__50351),
            .lcout(\ALU.c_RNIE4B6N4Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_16_LC_16_18_0 .C_ON=1'b0;
    defparam \CONTROL.g0_16_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_16_LC_16_18_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \CONTROL.g0_16_LC_16_18_0  (
            .in0(N__38248),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63463),
            .lcout(\CONTROL.increment28lto5_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_11_LC_16_18_1 .C_ON=1'b0;
    defparam \CONTROL.g0_11_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_11_LC_16_18_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \CONTROL.g0_11_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__63462),
            .in2(_gnd_net_),
            .in3(N__38249),
            .lcout(),
            .ltout(\CONTROL.increment28lto5_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_a7_4_LC_16_18_2 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_a7_4_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_a7_4_LC_16_18_2 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \CONTROL.g0_3_i_a7_4_LC_16_18_2  (
            .in0(N__48468),
            .in1(N__40826),
            .in2(N__36266),
            .in3(N__38209),
            .lcout(\CONTROL.g0_3_i_a7Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m221cf1_LC_16_18_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf1_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf1_LC_16_18_3 .LUT_INIT=16'b1000100000001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m221cf1_LC_16_18_3  (
            .in0(N__36206),
            .in1(N__74038),
            .in2(N__73412),
            .in3(N__72688),
            .lcout(\PROM.ROMDATA.m221cf1 ),
            .ltout(\PROM.ROMDATA.m221cf1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m221_LC_16_18_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m221_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m221_LC_16_18_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m221_LC_16_18_4  (
            .in0(N__45238),
            .in1(_gnd_net_),
            .in2(N__36251),
            .in3(N__36196),
            .lcout(PROM_ROMDATA_dintern_7ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_ne_0_LC_16_18_5 .C_ON=1'b0;
    defparam \CONTROL.operand1_ne_0_LC_16_18_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_ne_0_LC_16_18_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.operand1_ne_0_LC_16_18_5  (
            .in0(N__36197),
            .in1(N__36248),
            .in2(_gnd_net_),
            .in3(N__45239),
            .lcout(aluOperand1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand1_ne_0C_net ),
            .ce(N__36242),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m221cf0_LC_16_18_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf0_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf0_LC_16_18_6 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m221cf0_LC_16_18_6  (
            .in0(N__74037),
            .in1(N__36205),
            .in2(N__72742),
            .in3(N__73433),
            .lcout(\PROM.ROMDATA.m221cf0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_7_LC_16_18_7 .C_ON=1'b0;
    defparam \CONTROL.g0_7_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_7_LC_16_18_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \CONTROL.g0_7_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__63461),
            .in2(_gnd_net_),
            .in3(N__38247),
            .lcout(\CONTROL.increment28lto5_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState103_0_a2_1_LC_16_19_0 .C_ON=1'b0;
    defparam \CONTROL.un1_busState103_0_a2_1_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState103_0_a2_1_LC_16_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \CONTROL.un1_busState103_0_a2_1_LC_16_19_0  (
            .in0(N__54584),
            .in1(N__36878),
            .in2(N__36397),
            .in3(N__41210),
            .lcout(),
            .ltout(\CONTROL.N_320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState103_0_LC_16_19_1 .C_ON=1'b0;
    defparam \CONTROL.un1_busState103_0_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState103_0_LC_16_19_1 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \CONTROL.un1_busState103_0_LC_16_19_1  (
            .in0(N__36452),
            .in1(N__36377),
            .in2(N__36410),
            .in3(N__41201),
            .lcout(\CONTROL.un1_busState103_0_0 ),
            .ltout(\CONTROL.un1_busState103_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_1_0_LC_16_19_2 .C_ON=1'b0;
    defparam \CONTROL.aluParams_1_0_LC_16_19_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluParams_1_0_LC_16_19_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \CONTROL.aluParams_1_0_LC_16_19_2  (
            .in0(N__63030),
            .in1(N__36713),
            .in2(N__36407),
            .in3(N__41582),
            .lcout(aluParams_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluParams_1_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState103_0_o2_LC_16_19_3 .C_ON=1'b0;
    defparam \CONTROL.un1_busState103_0_o2_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState103_0_o2_LC_16_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \CONTROL.un1_busState103_0_o2_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__71820),
            .in2(_gnd_net_),
            .in3(N__44661),
            .lcout(\CONTROL.N_95_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState103_0_a2_LC_16_19_4 .C_ON=1'b0;
    defparam \CONTROL.un1_busState103_0_a2_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState103_0_a2_LC_16_19_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \CONTROL.un1_busState103_0_a2_LC_16_19_4  (
            .in0(N__54583),
            .in1(N__41396),
            .in2(N__41235),
            .in3(N__44871),
            .lcout(\CONTROL.N_318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNITJ3GK_12_LC_16_19_6 .C_ON=1'b0;
    defparam \ALU.c_RNITJ3GK_12_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNITJ3GK_12_LC_16_19_6 .LUT_INIT=16'b0111011001101000;
    LogicCell40 \ALU.c_RNITJ3GK_12_LC_16_19_6  (
            .in0(N__56910),
            .in1(N__74682),
            .in2(N__63076),
            .in3(N__61151),
            .lcout(\ALU.N_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNITVOEK_12_LC_16_19_7 .C_ON=1'b0;
    defparam \ALU.c_RNITVOEK_12_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNITVOEK_12_LC_16_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.c_RNITVOEK_12_LC_16_19_7  (
            .in0(N__61152),
            .in1(N__63026),
            .in2(_gnd_net_),
            .in3(N__56909),
            .lcout(\ALU.c_RNITVOEKZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA7CLH_8_LC_16_20_0 .C_ON=1'b0;
    defparam \ALU.d_RNIA7CLH_8_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA7CLH_8_LC_16_20_0 .LUT_INIT=16'b0111011001101000;
    LogicCell40 \ALU.d_RNIA7CLH_8_LC_16_20_0  (
            .in0(N__55812),
            .in1(N__74681),
            .in2(N__63075),
            .in3(N__61930),
            .lcout(\ALU.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_1_ne_RNO_0_1_LC_16_20_1 .C_ON=1'b0;
    defparam \CONTROL.aluParams_1_ne_RNO_0_1_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluParams_1_ne_RNO_0_1_LC_16_20_1 .LUT_INIT=16'b0010001100010011;
    LogicCell40 \CONTROL.aluParams_1_ne_RNO_0_1_LC_16_20_1  (
            .in0(N__44656),
            .in1(N__74815),
            .in2(N__41357),
            .in3(N__44869),
            .lcout(),
            .ltout(\CONTROL.N_340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_1_ne_1_LC_16_20_2 .C_ON=1'b0;
    defparam \CONTROL.aluParams_1_ne_1_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluParams_1_ne_1_LC_16_20_2 .LUT_INIT=16'b0000110000001011;
    LogicCell40 \CONTROL.aluParams_1_ne_1_LC_16_20_2  (
            .in0(N__44870),
            .in1(N__54585),
            .in2(N__36533),
            .in3(N__44657),
            .lcout(aluParams_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluParams_1_ne_1C_net ),
            .ce(N__36530),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAJ1KH_8_LC_16_20_3 .C_ON=1'b0;
    defparam \ALU.d_RNIAJ1KH_8_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAJ1KH_8_LC_16_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.d_RNIAJ1KH_8_LC_16_20_3  (
            .in0(N__61931),
            .in1(N__63022),
            .in2(_gnd_net_),
            .in3(N__55811),
            .lcout(\ALU.d_RNIAJ1KHZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState114_2_0_0_x1_LC_16_20_4 .C_ON=1'b0;
    defparam \CONTROL.un1_busState114_2_0_0_x1_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState114_2_0_0_x1_LC_16_20_4 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \CONTROL.un1_busState114_2_0_0_x1_LC_16_20_4  (
            .in0(N__44867),
            .in1(N__41305),
            .in2(N__54651),
            .in3(N__44654),
            .lcout(\CONTROL.un1_busState114_2_0_0_xZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState114_2_0_0_x0_LC_16_20_5 .C_ON=1'b0;
    defparam \CONTROL.un1_busState114_2_0_0_x0_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState114_2_0_0_x0_LC_16_20_5 .LUT_INIT=16'b1110010011111010;
    LogicCell40 \CONTROL.un1_busState114_2_0_0_x0_LC_16_20_5  (
            .in0(N__44655),
            .in1(N__54579),
            .in2(N__41356),
            .in3(N__44868),
            .lcout(),
            .ltout(\CONTROL.un1_busState114_2_0_0_xZ0Z0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState114_2_0_0_ns_LC_16_20_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState114_2_0_0_ns_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState114_2_0_0_ns_LC_16_20_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \CONTROL.un1_busState114_2_0_0_ns_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__71745),
            .in2(N__36518),
            .in3(N__36515),
            .lcout(\CONTROL.un1_busState114_2_0_0_0 ),
            .ltout(\CONTROL.un1_busState114_2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState114_2_0_LC_16_20_7 .C_ON=1'b0;
    defparam \CONTROL.un1_busState114_2_0_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState114_2_0_LC_16_20_7 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \CONTROL.un1_busState114_2_0_LC_16_20_7  (
            .in0(N__47033),
            .in1(N__46984),
            .in2(N__36509),
            .in3(N__54580),
            .lcout(\CONTROL.un1_busState114_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_4_LC_16_21_1 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_4_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_4_LC_16_21_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \CONTROL.aluOperation_4_LC_16_21_1  (
            .in0(N__38127),
            .in1(N__41203),
            .in2(N__69885),
            .in3(N__41394),
            .lcout(aluOperation_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluOperation_4C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_2_0_LC_16_21_2 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_2_0_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluReadBus_1_sqmuxa_0_a2_2_0_LC_16_21_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \CONTROL.aluReadBus_1_sqmuxa_0_a2_2_0_LC_16_21_2  (
            .in0(N__55451),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54539),
            .lcout(\CONTROL.aluReadBus_1_sqmuxa_0_a2_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState96_1_i_2_LC_16_21_3 .C_ON=1'b0;
    defparam \CONTROL.un1_busState96_1_i_2_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState96_1_i_2_LC_16_21_3 .LUT_INIT=16'b0000010001010001;
    LogicCell40 \CONTROL.un1_busState96_1_i_2_LC_16_21_3  (
            .in0(N__40963),
            .in1(N__41575),
            .in2(N__36487),
            .in3(N__41202),
            .lcout(\CONTROL.N_48_0 ),
            .ltout(\CONTROL.N_48_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_2_LC_16_21_4 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_2_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_2_LC_16_21_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \CONTROL.aluOperation_2_LC_16_21_4  (
            .in0(N__41576),
            .in1(N__70054),
            .in2(N__36635),
            .in3(N__36632),
            .lcout(aluOperation_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluOperation_4C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_RNO_0_2_LC_16_21_5 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_RNO_0_2_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_RNO_0_2_LC_16_21_5 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \CONTROL.aluOperation_RNO_0_2_LC_16_21_5  (
            .in0(N__54541),
            .in1(N__41393),
            .in2(N__71853),
            .in3(N__44650),
            .lcout(\CONTROL.un1_controlWord_14_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_RNO_1_LC_16_21_6 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_RNO_1_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluReadBus_RNO_1_LC_16_21_6 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \CONTROL.aluReadBus_RNO_1_LC_16_21_6  (
            .in0(N__41392),
            .in1(N__38699),
            .in2(N__36625),
            .in3(N__38623),
            .lcout(\CONTROL.un1_busState97_1_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment_5_0__m6_i_0_LC_16_21_7 .C_ON=1'b0;
    defparam \CONTROL.increment_5_0__m6_i_0_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment_5_0__m6_i_0_LC_16_21_7 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \CONTROL.increment_5_0__m6_i_0_LC_16_21_7  (
            .in0(N__54540),
            .in1(N__42221),
            .in2(N__72316),
            .in3(N__55452),
            .lcout(\CONTROL.un1_busState114_2_0_o2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNII6GE_7_LC_16_22_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNII6GE_7_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNII6GE_7_LC_16_22_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNII6GE_7_LC_16_22_0  (
            .in0(N__73319),
            .in1(N__36566),
            .in2(_gnd_net_),
            .in3(N__45145),
            .lcout(),
            .ltout(\CONTROL.N_422_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNII9UU_7_LC_16_22_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNII9UU_7_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNII9UU_7_LC_16_22_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNII9UU_7_LC_16_22_1  (
            .in0(N__36554),
            .in1(_gnd_net_),
            .in2(N__36539),
            .in3(N__73677),
            .lcout(progRomAddress_7),
            .ltout(progRomAddress_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_2_LC_16_22_2 .C_ON=1'b0;
    defparam \CONTROL.dout_2_LC_16_22_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_2_LC_16_22_2 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \CONTROL.dout_2_LC_16_22_2  (
            .in0(N__72263),
            .in1(N__41008),
            .in2(N__36536),
            .in3(N__45766),
            .lcout(\CONTROL.ctrlOut_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_2C_net ),
            .ce(N__44396),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m90_LC_16_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m90_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m90_LC_16_22_3 .LUT_INIT=16'b0110110110011100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m90_LC_16_22_3  (
            .in0(N__77862),
            .in1(N__78779),
            .in2(N__75984),
            .in3(N__77174),
            .lcout(\PROM.ROMDATA.m90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_3dflt_LC_16_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_3dflt_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_3dflt_LC_16_22_4 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \PROM.ROMDATA.dintern_3dflt_LC_16_22_4  (
            .in0(N__72262),
            .in1(N__41834),
            .in2(N__72606),
            .in3(N__64397),
            .lcout(controlWord_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIE2GE_5_LC_16_22_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIE2GE_5_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIE2GE_5_LC_16_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIE2GE_5_LC_16_22_5  (
            .in0(N__45146),
            .in1(N__45662),
            .in2(_gnd_net_),
            .in3(N__41723),
            .lcout(),
            .ltout(\CONTROL.N_420_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIC3UU_5_LC_16_22_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIC3UU_5_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIC3UU_5_LC_16_22_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIC3UU_5_LC_16_22_6  (
            .in0(N__73679),
            .in1(_gnd_net_),
            .in2(N__36746),
            .in3(N__41771),
            .lcout(\CONTROL.programCounter_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_1_cry_0_c_RNO_LC_16_22_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_1_cry_0_c_RNO_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_1_cry_0_c_RNO_LC_16_22_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \CONTROL.programCounter_1_cry_0_c_RNO_LC_16_22_7  (
            .in0(N__47407),
            .in1(N__73678),
            .in2(_gnd_net_),
            .in3(N__50962),
            .lcout(\CONTROL.programCounter_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_1_RNO_0_0_LC_16_23_0 .C_ON=1'b0;
    defparam \CONTROL.aluParams_1_RNO_0_0_LC_16_23_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluParams_1_RNO_0_0_LC_16_23_0 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \CONTROL.aluParams_1_RNO_0_0_LC_16_23_0  (
            .in0(N__41108),
            .in1(N__41424),
            .in2(N__72626),
            .in3(N__41810),
            .lcout(\CONTROL.N_105_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI1CMQ_12_LC_16_23_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI1CMQ_12_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI1CMQ_12_LC_16_23_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI1CMQ_12_LC_16_23_1  (
            .in0(N__42070),
            .in1(N__36755),
            .in2(_gnd_net_),
            .in3(N__38753),
            .lcout(\CONTROL.N_427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m177_LC_16_23_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m177_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m177_LC_16_23_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m177_LC_16_23_2  (
            .in0(N__47309),
            .in1(N__72503),
            .in2(_gnd_net_),
            .in3(N__64900),
            .lcout(PROM_ROMDATA_dintern_5ro),
            .ltout(PROM_ROMDATA_dintern_5ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState111_0_202_a2_0_o2_LC_16_23_3 .C_ON=1'b0;
    defparam \CONTROL.busState111_0_202_a2_0_o2_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState111_0_202_a2_0_o2_LC_16_23_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \CONTROL.busState111_0_202_a2_0_o2_LC_16_23_3  (
            .in0(N__71802),
            .in1(_gnd_net_),
            .in2(N__36692),
            .in3(N__72226),
            .lcout(\CONTROL.N_80_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_0_LC_16_23_4 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_0_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_0_LC_16_23_4 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_0_LC_16_23_4  (
            .in0(N__72227),
            .in1(N__42208),
            .in2(_gnd_net_),
            .in3(N__71803),
            .lcout(\CONTROL.N_98_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_1_i_3_1_LC_16_23_5 .C_ON=1'b0;
    defparam \CONTROL.g0_1_i_3_1_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_1_i_3_1_LC_16_23_5 .LUT_INIT=16'b0001110000001000;
    LogicCell40 \CONTROL.g0_1_i_3_1_LC_16_23_5  (
            .in0(N__71804),
            .in1(N__54573),
            .in2(N__42235),
            .in3(N__44639),
            .lcout(\CONTROL.g0_1_i_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState114_1_0_a2_LC_16_23_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState114_1_0_a2_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState114_1_0_a2_LC_16_23_6 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \CONTROL.un1_busState114_1_0_a2_LC_16_23_6  (
            .in0(N__44640),
            .in1(N__42212),
            .in2(_gnd_net_),
            .in3(N__71805),
            .lcout(),
            .ltout(\CONTROL.N_209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState114_1_0_0_LC_16_23_7 .C_ON=1'b0;
    defparam \CONTROL.un1_busState114_1_0_0_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState114_1_0_0_LC_16_23_7 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \CONTROL.un1_busState114_1_0_0_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(N__36879),
            .in2(N__36836),
            .in3(N__54574),
            .lcout(\CONTROL.un1_busState114_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_0_LC_16_24_0 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_0_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_0_LC_16_24_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \CONTROL.busState_cnst_2_0__m38_i_a2_0_LC_16_24_0  (
            .in0(N__41423),
            .in1(N__54632),
            .in2(N__38582),
            .in3(N__44884),
            .lcout(),
            .ltout(\CONTROL.N_349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m38_i_1_LC_16_24_1 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m38_i_1_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m38_i_1_LC_16_24_1 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \CONTROL.busState_cnst_2_0__m38_i_1_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(N__36788),
            .in2(N__36824),
            .in3(N__36813),
            .lcout(\CONTROL.m38_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_LC_16_24_2 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m38_i_a2_LC_16_24_2 .LUT_INIT=16'b0000000000110101;
    LogicCell40 \CONTROL.busState_cnst_2_0__m38_i_a2_LC_16_24_2  (
            .in0(N__51065),
            .in1(N__45343),
            .in2(N__72698),
            .in3(N__44883),
            .lcout(\CONTROL.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_12_LC_16_24_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_12_LC_16_24_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_12_LC_16_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_1_12_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36782),
            .lcout(\CONTROL.programCounter_1_reto_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73217),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_2_LC_16_24_4 .C_ON=1'b0;
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_2_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_2_LC_16_24_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \CONTROL.un1_busState_0_sqmuxa_i_a2_2_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(N__41655),
            .in2(_gnd_net_),
            .in3(N__38567),
            .lcout(\CONTROL.N_362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_1dflt_LC_16_24_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_1dflt_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_1dflt_LC_16_24_5 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \PROM.ROMDATA.dintern_1dflt_LC_16_24_5  (
            .in0(N__72608),
            .in1(N__51064),
            .in2(N__45344),
            .in3(N__72224),
            .lcout(controlWord_1),
            .ltout(controlWord_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState_1_sqmuxa_i_a2_1_LC_16_24_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_a2_1_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState_1_sqmuxa_i_a2_1_LC_16_24_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \CONTROL.un1_busState_1_sqmuxa_i_a2_1_LC_16_24_6  (
            .in0(N__72225),
            .in1(_gnd_net_),
            .in2(N__36749),
            .in3(N__38566),
            .lcout(\CONTROL.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState97_i_i_o2_0_LC_16_26_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState97_i_i_o2_0_LC_16_26_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState97_i_i_o2_0_LC_16_26_2 .LUT_INIT=16'b0000101100001001;
    LogicCell40 \CONTROL.un1_busState97_i_i_o2_0_LC_16_26_2  (
            .in0(N__41580),
            .in1(N__41256),
            .in2(N__40962),
            .in3(N__41434),
            .lcout(\CONTROL.N_136_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m506_LC_16_26_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m506_LC_16_26_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m506_LC_16_26_4 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m506_LC_16_26_4  (
            .in0(N__74487),
            .in1(N__76600),
            .in2(N__65029),
            .in3(N__75907),
            .lcout(),
            .ltout(\PROM.ROMDATA.m506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m508_LC_16_26_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m508_LC_16_26_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m508_LC_16_26_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m508_LC_16_26_5  (
            .in0(_gnd_net_),
            .in1(N__79503),
            .in2(N__36953),
            .in3(N__79897),
            .lcout(\PROM.ROMDATA.N_571_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI64MA6_0_LC_17_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNI64MA6_0_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI64MA6_0_LC_17_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNI64MA6_0_LC_17_8_1  (
            .in0(N__71471),
            .in1(N__36932),
            .in2(_gnd_net_),
            .in3(N__37874),
            .lcout(\ALU.d_RNI64MA6Z0Z_0 ),
            .ltout(\ALU.d_RNI64MA6Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_21_0_LC_17_8_2 .C_ON=1'b0;
    defparam \ALU.status_RNO_21_0_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_21_0_LC_17_8_2 .LUT_INIT=16'b0011001111110000;
    LogicCell40 \ALU.status_RNO_21_0_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__39040),
            .in2(N__36899),
            .in3(N__53298),
            .lcout(),
            .ltout(\ALU.log_1_3_ns_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_17_0_LC_17_8_3 .C_ON=1'b0;
    defparam \ALU.status_RNO_17_0_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_17_0_LC_17_8_3 .LUT_INIT=16'b1111110011000011;
    LogicCell40 \ALU.status_RNO_17_0_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__63254),
            .in2(N__36896),
            .in3(N__60616),
            .lcout(),
            .ltout(\ALU.log_1_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_11_0_LC_17_8_4 .C_ON=1'b0;
    defparam \ALU.status_RNO_11_0_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_11_0_LC_17_8_4 .LUT_INIT=16'b0011010010101100;
    LogicCell40 \ALU.status_RNO_11_0_LC_17_8_4  (
            .in0(N__63255),
            .in1(N__74895),
            .in2(N__36893),
            .in3(N__66716),
            .lcout(),
            .ltout(\ALU.log_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_5_0_LC_17_8_5 .C_ON=1'b0;
    defparam \ALU.status_RNO_5_0_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_5_0_LC_17_8_5 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \ALU.status_RNO_5_0_LC_17_8_5  (
            .in0(N__63256),
            .in1(N__37193),
            .in2(N__36890),
            .in3(N__37373),
            .lcout(),
            .ltout(\ALU.status_8_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_2_0_LC_17_8_6 .C_ON=1'b0;
    defparam \ALU.status_RNO_2_0_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_2_0_LC_17_8_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ALU.status_RNO_2_0_LC_17_8_6  (
            .in0(N__48176),
            .in1(N__51458),
            .in2(N__36887),
            .in3(N__51203),
            .lcout(\ALU.status_RNO_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_365_c_LC_17_9_0 .C_ON=1'b1;
    defparam \ALU.mult_365_c_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_365_c_LC_17_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_365_c_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__37052),
            .in2(N__37385),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\ALU.mult_13_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_365_c_RNINK1M82_LC_17_9_1 .C_ON=1'b1;
    defparam \ALU.mult_365_c_RNINK1M82_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_365_c_RNINK1M82_LC_17_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_365_c_RNINK1M82_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__37040),
            .in2(N__37028),
            .in3(N__37016),
            .lcout(\ALU.mult_13_14 ),
            .ltout(),
            .carryin(\ALU.mult_13_c13 ),
            .carryout(\ALU.mult_13_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_371_c_RNIAJLO71_LC_17_9_2 .C_ON=1'b0;
    defparam \ALU.mult_371_c_RNIAJLO71_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_371_c_RNIAJLO71_LC_17_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.mult_371_c_RNIAJLO71_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__37013),
            .in2(_gnd_net_),
            .in3(N__37004),
            .lcout(\ALU.mult_13_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_365_c_RNI8ALO96_LC_17_9_3 .C_ON=1'b0;
    defparam \ALU.mult_365_c_RNI8ALO96_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_365_c_RNI8ALO96_LC_17_9_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALU.mult_365_c_RNI8ALO96_LC_17_9_3  (
            .in0(N__63835),
            .in1(N__38821),
            .in2(N__42377),
            .in3(N__66714),
            .lcout(\ALU.mult_365_c_RNI8ALOZ0Z96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIL4PC21_6_LC_17_9_4 .C_ON=1'b0;
    defparam \ALU.d_RNIL4PC21_6_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIL4PC21_6_LC_17_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIL4PC21_6_LC_17_9_4  (
            .in0(N__62232),
            .in1(N__55958),
            .in2(N__56130),
            .in3(N__62558),
            .lcout(\ALU.d_RNIL4PC21Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9VEDD1_4_LC_17_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNI9VEDD1_4_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9VEDD1_4_LC_17_9_7 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.d_RNI9VEDD1_4_LC_17_9_7  (
            .in0(N__59620),
            .in1(N__65990),
            .in2(N__59912),
            .in3(N__66713),
            .lcout(\ALU.mult_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_546_c_LC_17_10_0 .C_ON=1'b1;
    defparam \ALU.mult_546_c_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_546_c_LC_17_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_546_c_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__48790),
            .in2(N__48772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\ALU.mult_29_c8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_546_c_RNIUNL1A8_LC_17_10_1 .C_ON=1'b1;
    defparam \ALU.mult_546_c_RNIUNL1A8_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_546_c_RNIUNL1A8_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_546_c_RNIUNL1A8_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__36980),
            .in2(N__36968),
            .in3(N__36959),
            .lcout(\ALU.mult_9 ),
            .ltout(),
            .carryin(\ALU.mult_29_c8 ),
            .carryout(\ALU.mult_29_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_549_c_RNIV9413G_LC_17_10_2 .C_ON=1'b1;
    defparam \ALU.mult_549_c_RNIV9413G_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_549_c_RNIV9413G_LC_17_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_549_c_RNIV9413G_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__42437),
            .in2(N__42463),
            .in3(N__36956),
            .lcout(\ALU.mult_10 ),
            .ltout(),
            .carryin(\ALU.mult_29_c9 ),
            .carryout(\ALU.mult_29_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_552_c_RNIK1H74A_LC_17_10_3 .C_ON=1'b1;
    defparam \ALU.mult_552_c_RNIK1H74A_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_552_c_RNIK1H74A_LC_17_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_552_c_RNIK1H74A_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__42416),
            .in2(N__37172),
            .in3(N__37163),
            .lcout(\ALU.mult_11 ),
            .ltout(),
            .carryin(\ALU.mult_29_c10 ),
            .carryout(\ALU.mult_29_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_555_c_RNI9QLKVH_LC_17_10_4 .C_ON=1'b1;
    defparam \ALU.mult_555_c_RNI9QLKVH_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_555_c_RNI9QLKVH_LC_17_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_555_c_RNI9QLKVH_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__38957),
            .in2(N__38977),
            .in3(N__37160),
            .lcout(\ALU.mult_12 ),
            .ltout(),
            .carryin(\ALU.mult_29_c11 ),
            .carryout(\ALU.mult_29_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_558_c_RNIN3VB2C_LC_17_10_5 .C_ON=1'b1;
    defparam \ALU.mult_558_c_RNIN3VB2C_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_558_c_RNIN3VB2C_LC_17_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_558_c_RNIN3VB2C_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__37157),
            .in2(N__38930),
            .in3(N__37151),
            .lcout(\ALU.mult_13 ),
            .ltout(),
            .carryin(\ALU.mult_29_c12 ),
            .carryout(\ALU.mult_29_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_561_c_RNIL4S0IG_LC_17_10_6 .C_ON=1'b1;
    defparam \ALU.mult_561_c_RNIL4S0IG_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_561_c_RNIL4S0IG_LC_17_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_561_c_RNIL4S0IG_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__37148),
            .in2(N__38909),
            .in3(N__37142),
            .lcout(\ALU.mult_14 ),
            .ltout(),
            .carryin(\ALU.mult_29_c13 ),
            .carryout(\ALU.mult_29_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_564_c_RNIRTQTDC_LC_17_10_7 .C_ON=1'b0;
    defparam \ALU.mult_564_c_RNIRTQTDC_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_564_c_RNIRTQTDC_LC_17_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.mult_564_c_RNIRTQTDC_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__37139),
            .in2(_gnd_net_),
            .in3(N__37133),
            .lcout(\ALU.mult_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_9_c_RNI0ALKH7_LC_17_11_0 .C_ON=1'b0;
    defparam \ALU.addsub_cry_9_c_RNI0ALKH7_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_9_c_RNI0ALKH7_LC_17_11_0 .LUT_INIT=16'b0000001110100011;
    LogicCell40 \ALU.addsub_cry_9_c_RNI0ALKH7_LC_17_11_0  (
            .in0(N__39244),
            .in1(N__61505),
            .in2(N__66902),
            .in3(N__68459),
            .lcout(\ALU.a_15_am_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_549_c_RNIB6TIDG_LC_17_11_1 .C_ON=1'b0;
    defparam \ALU.mult_549_c_RNIB6TIDG_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_549_c_RNIB6TIDG_LC_17_11_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \ALU.mult_549_c_RNIB6TIDG_LC_17_11_1  (
            .in0(N__59044),
            .in1(N__37130),
            .in2(_gnd_net_),
            .in3(N__37094),
            .lcout(),
            .ltout(\ALU.mult_549_c_RNIB6TIDGZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_549_c_RNIE7260O_LC_17_11_2 .C_ON=1'b0;
    defparam \ALU.mult_549_c_RNIE7260O_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_549_c_RNIE7260O_LC_17_11_2 .LUT_INIT=16'b1011101001010100;
    LogicCell40 \ALU.mult_549_c_RNIE7260O_LC_17_11_2  (
            .in0(N__66901),
            .in1(N__67047),
            .in2(N__37088),
            .in3(N__37085),
            .lcout(\ALU.mult_549_c_RNIE7260OZ0 ),
            .ltout(\ALU.mult_549_c_RNIE7260OZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_10_LC_17_11_3 .C_ON=1'b0;
    defparam \ALU.a_10_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \ALU.a_10_LC_17_11_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.a_10_LC_17_11_3  (
            .in0(N__58455),
            .in1(_gnd_net_),
            .in2(N__37079),
            .in3(N__58343),
            .lcout(\ALU.aZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73141),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m3_s_13_LC_17_11_4 .C_ON=1'b0;
    defparam \ALU.a_15_m3_s_13_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m3_s_13_LC_17_11_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ALU.a_15_m3_s_13_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__59043),
            .in2(_gnd_net_),
            .in3(N__59295),
            .lcout(\ALU.a_15_m3_sZ0Z_13 ),
            .ltout(\ALU.a_15_m3_sZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_s_13_LC_17_11_5 .C_ON=1'b0;
    defparam \ALU.a_15_s_13_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_s_13_LC_17_11_5 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ALU.a_15_s_13_LC_17_11_5  (
            .in0(N__67046),
            .in1(_gnd_net_),
            .in2(N__37244),
            .in3(_gnd_net_),
            .lcout(\ALU.a_15_sZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a32_0_LC_17_11_6 .C_ON=1'b0;
    defparam \ALU.a32_0_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a32_0_LC_17_11_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ALU.a32_0_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__59042),
            .in2(_gnd_net_),
            .in3(N__67045),
            .lcout(\ALU.a32Z0Z_0 ),
            .ltout(\ALU.a32Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_1_LC_17_11_7 .C_ON=1'b0;
    defparam \ALU.a_1_LC_17_11_7 .SEQ_MODE=4'b1000;
    defparam \ALU.a_1_LC_17_11_7 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.a_1_LC_17_11_7  (
            .in0(N__59296),
            .in1(N__52205),
            .in2(N__37241),
            .in3(N__69014),
            .lcout(\ALU.aZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73141),
            .ce(N__71211),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICUA7B5_0_LC_17_12_0 .C_ON=1'b0;
    defparam \ALU.d_RNICUA7B5_0_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICUA7B5_0_LC_17_12_0 .LUT_INIT=16'b0000100011111101;
    LogicCell40 \ALU.d_RNICUA7B5_0_LC_17_12_0  (
            .in0(N__70168),
            .in1(N__37178),
            .in2(N__59139),
            .in3(N__40175),
            .lcout(),
            .ltout(\ALU.d_RNICUA7B5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_0_c_RNI43EE86_LC_17_12_1 .C_ON=1'b0;
    defparam \ALU.addsub_cry_0_c_RNI43EE86_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_0_c_RNI43EE86_LC_17_12_1 .LUT_INIT=16'b0000001111001111;
    LogicCell40 \ALU.addsub_cry_0_c_RNI43EE86_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__67044),
            .in2(N__37208),
            .in3(N__60326),
            .lcout(\ALU.a_15_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIL3JT71_0_LC_17_12_2 .C_ON=1'b0;
    defparam \ALU.d_RNIL3JT71_0_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIL3JT71_0_LC_17_12_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNIL3JT71_0_LC_17_12_2  (
            .in0(N__56929),
            .in1(N__65556),
            .in2(N__56804),
            .in3(N__60602),
            .lcout(\ALU.d_RNIL3JT71Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5A8KO_1_LC_17_12_3 .C_ON=1'b0;
    defparam \ALU.d_RNI5A8KO_1_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5A8KO_1_LC_17_12_3 .LUT_INIT=16'b0110011010001000;
    LogicCell40 \ALU.d_RNI5A8KO_1_LC_17_12_3  (
            .in0(N__74853),
            .in1(N__65551),
            .in2(_gnd_net_),
            .in3(N__65926),
            .lcout(\ALU.N_556 ),
            .ltout(\ALU.N_556_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3MGBH1_1_LC_17_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNI3MGBH1_1_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3MGBH1_1_LC_17_12_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \ALU.d_RNI3MGBH1_1_LC_17_12_4  (
            .in0(N__70167),
            .in1(N__63291),
            .in2(N__37181),
            .in3(N__37369),
            .lcout(\ALU.d_RNI3MGBH1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_39_c_RNO_LC_17_12_5 .C_ON=1'b0;
    defparam \ALU.status_17_I_39_c_RNO_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_39_c_RNO_LC_17_12_5 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \ALU.status_17_I_39_c_RNO_LC_17_12_5  (
            .in0(N__60965),
            .in1(N__56787),
            .in2(N__61216),
            .in3(N__56928),
            .lcout(\ALU.status_17_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_365_c_RNO_0_LC_17_12_6 .C_ON=1'b0;
    defparam \ALU.mult_365_c_RNO_0_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_365_c_RNO_0_LC_17_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_365_c_RNO_0_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__60964),
            .in2(_gnd_net_),
            .in3(N__66582),
            .lcout(\ALU.mult_365_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5A8KO_0_1_LC_17_12_7 .C_ON=1'b0;
    defparam \ALU.d_RNI5A8KO_0_1_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5A8KO_0_1_LC_17_12_7 .LUT_INIT=16'b0101010111101110;
    LogicCell40 \ALU.d_RNI5A8KO_0_1_LC_17_12_7  (
            .in0(N__74854),
            .in1(N__65552),
            .in2(_gnd_net_),
            .in3(N__65927),
            .lcout(\ALU.N_572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_10_c_RNISV0175_LC_17_13_0 .C_ON=1'b0;
    defparam \ALU.addsub_cry_10_c_RNISV0175_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_10_c_RNISV0175_LC_17_13_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.addsub_cry_10_c_RNISV0175_LC_17_13_0  (
            .in0(N__69944),
            .in1(N__61276),
            .in2(N__69679),
            .in3(N__37292),
            .lcout(\ALU.a_15_am_rn_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_552_c_RNI70R9DA_LC_17_13_1 .C_ON=1'b0;
    defparam \ALU.mult_552_c_RNI70R9DA_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_552_c_RNI70R9DA_LC_17_13_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.mult_552_c_RNI70R9DA_LC_17_13_1  (
            .in0(N__37341),
            .in1(N__69645),
            .in2(_gnd_net_),
            .in3(N__37304),
            .lcout(\ALU.mult_552_c_RNI70R9DAZ0 ),
            .ltout(\ALU.mult_552_c_RNI70R9DAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_552_c_RNIOT7VLF_0_LC_17_13_2 .C_ON=1'b0;
    defparam \ALU.mult_552_c_RNIOT7VLF_0_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_552_c_RNIOT7VLF_0_LC_17_13_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ALU.mult_552_c_RNIOT7VLF_0_LC_17_13_2  (
            .in0(N__37285),
            .in1(N__43037),
            .in2(N__37295),
            .in3(N__37532),
            .lcout(\ALU.mult_552_c_RNIOT7VLFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIP0VNF4_15_LC_17_13_3 .C_ON=1'b0;
    defparam \ALU.c_RNIP0VNF4_15_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIP0VNF4_15_LC_17_13_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ALU.c_RNIP0VNF4_15_LC_17_13_3  (
            .in0(N__43184),
            .in1(N__68464),
            .in2(N__42872),
            .in3(N__68809),
            .lcout(\ALU.rshift_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_552_c_RNIOT7VLF_LC_17_13_4 .C_ON=1'b0;
    defparam \ALU.mult_552_c_RNIOT7VLF_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_552_c_RNIOT7VLF_LC_17_13_4 .LUT_INIT=16'b1111111011011100;
    LogicCell40 \ALU.mult_552_c_RNIOT7VLF_LC_17_13_4  (
            .in0(N__37531),
            .in1(N__43038),
            .in2(N__37286),
            .in3(N__37274),
            .lcout(\ALU.mult_552_c_RNIOT7VLFZ0 ),
            .ltout(\ALU.mult_552_c_RNIOT7VLFZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_11_LC_17_13_5 .C_ON=1'b0;
    defparam \ALU.a_11_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.a_11_LC_17_13_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.a_11_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__58165),
            .in2(N__37268),
            .in3(N__58111),
            .lcout(\ALU.aZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73146),
            .ce(N__71216),
            .sr(_gnd_net_));
    defparam \ALU.a_15_am_sn_11_LC_17_13_6 .C_ON=1'b0;
    defparam \ALU.a_15_am_sn_11_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_am_sn_11_LC_17_13_6 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \ALU.a_15_am_sn_11_LC_17_13_6  (
            .in0(N__69641),
            .in1(N__67043),
            .in2(_gnd_net_),
            .in3(N__69943),
            .lcout(\ALU.a_15_am_snZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_1_LC_17_14_0 .C_ON=1'b0;
    defparam \ALU.h_1_LC_17_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_1_LC_17_14_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.h_1_LC_17_14_0  (
            .in0(N__59298),
            .in1(N__52223),
            .in2(N__69666),
            .in3(N__69013),
            .lcout(h_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73151),
            .ce(N__69453),
            .sr(_gnd_net_));
    defparam \ALU.a_15_s_11_LC_17_14_1 .C_ON=1'b0;
    defparam \ALU.a_15_s_11_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_s_11_LC_17_14_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.a_15_s_11_LC_17_14_1  (
            .in0(N__69646),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59297),
            .lcout(\ALU.a_15_sZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_489_c_RNIGEUL1A_LC_17_14_2 .C_ON=1'b0;
    defparam \ALU.mult_489_c_RNIGEUL1A_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_489_c_RNIGEUL1A_LC_17_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.mult_489_c_RNIGEUL1A_LC_17_14_2  (
            .in0(N__67042),
            .in1(N__62345),
            .in2(_gnd_net_),
            .in3(N__37478),
            .lcout(\ALU.mult_489_c_RNIGEUL1AZ0 ),
            .ltout(\ALU.mult_489_c_RNIGEUL1AZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_489_c_RNIPGBQMC_LC_17_14_3 .C_ON=1'b0;
    defparam \ALU.mult_489_c_RNIPGBQMC_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_489_c_RNIPGBQMC_LC_17_14_3 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \ALU.mult_489_c_RNIPGBQMC_LC_17_14_3  (
            .in0(N__69647),
            .in1(N__52678),
            .in2(N__37466),
            .in3(N__63319),
            .lcout(\ALU.mult_489_c_RNIPGBQMCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_489_c_RNIPGBQMC_0_LC_17_14_5 .C_ON=1'b0;
    defparam \ALU.mult_489_c_RNIPGBQMC_0_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_489_c_RNIPGBQMC_0_LC_17_14_5 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ALU.mult_489_c_RNIPGBQMC_0_LC_17_14_5  (
            .in0(N__52679),
            .in1(N__63320),
            .in2(N__69680),
            .in3(N__37463),
            .lcout(),
            .ltout(\ALU.mult_489_c_RNIPGBQMCZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_489_c_RNI1J3GCU_LC_17_14_6 .C_ON=1'b0;
    defparam \ALU.mult_489_c_RNI1J3GCU_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_489_c_RNI1J3GCU_LC_17_14_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.mult_489_c_RNI1J3GCU_LC_17_14_6  (
            .in0(N__39209),
            .in1(_gnd_net_),
            .in2(N__37457),
            .in3(N__37454),
            .lcout(\ALU.mult_489_c_RNI1J3GCUZ0 ),
            .ltout(\ALU.mult_489_c_RNI1J3GCUZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_6_LC_17_14_7 .C_ON=1'b0;
    defparam \ALU.h_6_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \ALU.h_6_LC_17_14_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.h_6_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(N__43039),
            .in2(N__37448),
            .in3(N__43104),
            .lcout(h_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73151),
            .ce(N__69453),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4HL061_0_LC_17_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNI4HL061_0_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4HL061_0_LC_17_15_0 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \ALU.d_RNI4HL061_0_LC_17_15_0  (
            .in0(N__66685),
            .in1(N__60365),
            .in2(N__67204),
            .in3(N__60566),
            .lcout(\ALU.d_RNI4HL061Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA4TMK_0_LC_17_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIA4TMK_0_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA4TMK_0_LC_17_15_1 .LUT_INIT=16'b0010110111010100;
    LogicCell40 \ALU.d_RNIA4TMK_0_LC_17_15_1  (
            .in0(N__50541),
            .in1(N__60572),
            .in2(N__74832),
            .in3(N__66686),
            .lcout(),
            .ltout(\ALU.a_15_m2_d_d_ns_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4D6E01_0_LC_17_15_2 .C_ON=1'b0;
    defparam \ALU.d_RNI4D6E01_0_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4D6E01_0_LC_17_15_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \ALU.d_RNI4D6E01_0_LC_17_15_2  (
            .in0(N__59282),
            .in1(N__50542),
            .in2(N__37691),
            .in3(N__37659),
            .lcout(),
            .ltout(\ALU.d_RNI4D6E01Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQQ9O83_0_LC_17_15_3 .C_ON=1'b0;
    defparam \ALU.d_RNIQQ9O83_0_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQQ9O83_0_LC_17_15_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ALU.d_RNIQQ9O83_0_LC_17_15_3  (
            .in0(N__59328),
            .in1(N__37636),
            .in2(N__37604),
            .in3(N__60573),
            .lcout(),
            .ltout(\ALU.d_RNIQQ9O83Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINUGCF4_0_LC_17_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNINUGCF4_0_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINUGCF4_0_LC_17_15_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNINUGCF4_0_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__69651),
            .in2(N__37601),
            .in3(N__37598),
            .lcout(\ALU.d_RNINUGCF4Z0Z_0 ),
            .ltout(\ALU.d_RNINUGCF4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_0_LC_17_15_5 .C_ON=1'b0;
    defparam \ALU.a_0_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \ALU.a_0_LC_17_15_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ALU.a_0_LC_17_15_5  (
            .in0(N__69160),
            .in1(N__69627),
            .in2(N__37592),
            .in3(N__52055),
            .lcout(\ALU.aZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73154),
            .ce(N__71193),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_s_15_LC_17_15_6 .C_ON=1'b0;
    defparam \ALU.a_15_m2_s_15_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_s_15_LC_17_15_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ALU.a_15_m2_s_15_LC_17_15_6  (
            .in0(N__59281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__70139),
            .lcout(\ALU.a_15_m2_sZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI933S_0_LC_17_15_7 .C_ON=1'b0;
    defparam \ALU.e_RNI933S_0_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI933S_0_LC_17_15_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.e_RNI933S_0_LC_17_15_7  (
            .in0(N__46325),
            .in1(N__37579),
            .in2(_gnd_net_),
            .in3(N__53572),
            .lcout(\ALU.e_RNI933SZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_0_LC_17_16_0 .C_ON=1'b0;
    defparam \ALU.h_0_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_0_LC_17_16_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \ALU.h_0_LC_17_16_0  (
            .in0(N__52080),
            .in1(N__69161),
            .in2(N__69689),
            .in3(N__52054),
            .lcout(h_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73160),
            .ce(N__69450),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0G5D_0_LC_17_16_1 .C_ON=1'b0;
    defparam \ALU.d_RNI0G5D_0_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0G5D_0_LC_17_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNI0G5D_0_LC_17_16_1  (
            .in0(N__43983),
            .in1(N__37548),
            .in2(_gnd_net_),
            .in3(N__51967),
            .lcout(\ALU.d_RNI0G5DZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIDFF01_0_LC_17_16_2 .C_ON=1'b0;
    defparam \ALU.c_RNIDFF01_0_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIDFF01_0_LC_17_16_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIDFF01_0_LC_17_16_2  (
            .in0(N__48901),
            .in1(N__46429),
            .in2(_gnd_net_),
            .in3(N__53573),
            .lcout(),
            .ltout(\ALU.c_RNIDFF01Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNITEVO2_0_LC_17_16_3 .C_ON=1'b0;
    defparam \ALU.e_RNITEVO2_0_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNITEVO2_0_LC_17_16_3 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.e_RNITEVO2_0_LC_17_16_3  (
            .in0(N__53859),
            .in1(N__37898),
            .in2(N__37892),
            .in3(N__53410),
            .lcout(\ALU.operand2_7_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIS3PO_0_LC_17_16_4 .C_ON=1'b0;
    defparam \ALU.b_RNIS3PO_0_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIS3PO_0_LC_17_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.b_RNIS3PO_0_LC_17_16_4  (
            .in0(N__49131),
            .in1(N__48380),
            .in2(_gnd_net_),
            .in3(N__43982),
            .lcout(),
            .ltout(\ALU.b_RNIS3POZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITCRC4_0_LC_17_16_5 .C_ON=1'b0;
    defparam \ALU.d_RNITCRC4_0_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITCRC4_0_LC_17_16_5 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \ALU.d_RNITCRC4_0_LC_17_16_5  (
            .in0(N__53860),
            .in1(N__37889),
            .in2(N__37883),
            .in3(N__37880),
            .lcout(\ALU.operand2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNICGJM_9_LC_17_16_6 .C_ON=1'b0;
    defparam \ALU.e_RNICGJM_9_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNICGJM_9_LC_17_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.e_RNICGJM_9_LC_17_16_6  (
            .in0(N__46207),
            .in1(N__43552),
            .in2(_gnd_net_),
            .in3(N__43981),
            .lcout(\ALU.e_RNICGJMZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI3E5B1_3_LC_17_17_0 .C_ON=1'b0;
    defparam \ALU.b_RNI3E5B1_3_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI3E5B1_3_LC_17_17_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI3E5B1_3_LC_17_17_0  (
            .in0(N__39862),
            .in1(N__53570),
            .in2(N__44235),
            .in3(N__53466),
            .lcout(),
            .ltout(\ALU.operand2_6_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8SEV1_3_LC_17_17_1 .C_ON=1'b0;
    defparam \ALU.d_RNI8SEV1_3_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8SEV1_3_LC_17_17_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.d_RNI8SEV1_3_LC_17_17_1  (
            .in0(N__37843),
            .in1(N__58602),
            .in2(N__37829),
            .in3(N__53405),
            .lcout(\ALU.N_1248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI18V81_3_LC_17_17_2 .C_ON=1'b0;
    defparam \ALU.e_RNI18V81_3_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI18V81_3_LC_17_17_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNI18V81_3_LC_17_17_2  (
            .in0(N__37826),
            .in1(N__53571),
            .in2(N__37802),
            .in3(N__53467),
            .lcout(),
            .ltout(\ALU.operand2_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI4G2B2_3_LC_17_17_3 .C_ON=1'b0;
    defparam \ALU.c_RNI4G2B2_3_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI4G2B2_3_LC_17_17_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.c_RNI4G2B2_3_LC_17_17_3  (
            .in0(N__37769),
            .in1(N__37737),
            .in2(N__37694),
            .in3(N__53406),
            .lcout(),
            .ltout(\ALU.N_1200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGMEO4_3_LC_17_17_4 .C_ON=1'b0;
    defparam \ALU.d_RNIGMEO4_3_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGMEO4_3_LC_17_17_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIGMEO4_3_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__53861),
            .in2(N__38093),
            .in3(N__38090),
            .lcout(),
            .ltout(\ALU.d_RNIGMEO4Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2CUG6_3_LC_17_17_5 .C_ON=1'b0;
    defparam \ALU.d_RNI2CUG6_3_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2CUG6_3_LC_17_17_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNI2CUG6_3_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__71400),
            .in2(N__38084),
            .in3(N__38081),
            .lcout(\ALU.d_RNI2CUG6Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNI4KOJ_4_LC_17_17_6 .C_ON=1'b0;
    defparam \CONTROL.dout_RNI4KOJ_4_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNI4KOJ_4_LC_17_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNI4KOJ_4_LC_17_17_6  (
            .in0(N__38027),
            .in1(N__55334),
            .in2(_gnd_net_),
            .in3(N__50168),
            .lcout(\CONTROL.N_165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_9_LC_17_18_0 .C_ON=1'b0;
    defparam \ALU.h_9_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_9_LC_17_18_0 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \ALU.h_9_LC_17_18_0  (
            .in0(N__66845),
            .in1(N__58498),
            .in2(N__52889),
            .in3(N__52808),
            .lcout(h_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73181),
            .ce(N__69454),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKKNJ_9_LC_17_18_1 .C_ON=1'b0;
    defparam \ALU.d_RNIKKNJ_9_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKKNJ_9_LC_17_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIKKNJ_9_LC_17_18_1  (
            .in0(N__43242),
            .in1(N__37941),
            .in2(_gnd_net_),
            .in3(N__52744),
            .lcout(\ALU.d_RNIKKNJZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIG8BV_9_LC_17_18_2 .C_ON=1'b0;
    defparam \ALU.b_RNIG8BV_9_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIG8BV_9_LC_17_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.b_RNIG8BV_9_LC_17_18_2  (
            .in0(N__48832),
            .in1(N__48981),
            .in2(_gnd_net_),
            .in3(N__43243),
            .lcout(\ALU.b_RNIG8BVZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI65HE2_9_LC_17_18_3 .C_ON=1'b0;
    defparam \ALU.e_RNI65HE2_9_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI65HE2_9_LC_17_18_3 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \ALU.e_RNI65HE2_9_LC_17_18_3  (
            .in0(N__37925),
            .in1(N__43415),
            .in2(N__53940),
            .in3(N__46782),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIECHF4_9_LC_17_18_4 .C_ON=1'b0;
    defparam \ALU.d_RNIECHF4_9_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIECHF4_9_LC_17_18_4 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNIECHF4_9_LC_17_18_4  (
            .in0(N__37916),
            .in1(N__53898),
            .in2(N__37910),
            .in3(N__37907),
            .lcout(),
            .ltout(\ALU.operand2_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4K8P6_9_LC_17_18_5 .C_ON=1'b0;
    defparam \ALU.d_RNI4K8P6_9_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4K8P6_9_LC_17_18_5 .LUT_INIT=16'b1010111100100111;
    LogicCell40 \ALU.d_RNI4K8P6_9_LC_17_18_5  (
            .in0(N__71401),
            .in1(N__40400),
            .in2(N__37901),
            .in3(N__49825),
            .lcout(\ALU.combOperand2_0_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_0_LC_17_19_0 .C_ON=1'b0;
    defparam \ALU.status_0_LC_17_19_0 .SEQ_MODE=4'b1000;
    defparam \ALU.status_0_LC_17_19_0 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.status_0_LC_17_19_0  (
            .in0(N__56573),
            .in1(N__38303),
            .in2(N__38285),
            .in3(N__48425),
            .lcout(aluStatus_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73190),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_0_0_LC_17_19_1 .C_ON=1'b0;
    defparam \ALU.status_RNO_0_0_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_0_0_LC_17_19_1 .LUT_INIT=16'b0011010100110011;
    LogicCell40 \ALU.status_RNO_0_0_LC_17_19_1  (
            .in0(N__56532),
            .in1(N__48463),
            .in2(N__71504),
            .in3(N__69318),
            .lcout(\ALU.status_e_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_LC_17_19_2 .C_ON=1'b0;
    defparam \ALU.un1_a41_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_LC_17_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ALU.un1_a41_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__69317),
            .in2(_gnd_net_),
            .in3(N__71500),
            .lcout(\ALU.un1_a41_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment28lto5_1_1_LC_17_19_3 .C_ON=1'b0;
    defparam \CONTROL.increment28lto5_1_1_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment28lto5_1_1_LC_17_19_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \CONTROL.increment28lto5_1_1_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__63459),
            .in2(_gnd_net_),
            .in3(N__38264),
            .lcout(),
            .ltout(\CONTROL.increment28lto5_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment28lto5_LC_17_19_4 .C_ON=1'b0;
    defparam \CONTROL.increment28lto5_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment28lto5_LC_17_19_4 .LUT_INIT=16'b1000000001010101;
    LogicCell40 \CONTROL.increment28lto5_LC_17_19_4  (
            .in0(N__72252),
            .in1(N__41018),
            .in2(N__38276),
            .in3(N__38160),
            .lcout(\CONTROL.N_361_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_14_LC_17_19_5 .C_ON=1'b0;
    defparam \CONTROL.g0_14_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_14_LC_17_19_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \CONTROL.g0_14_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__63460),
            .in2(_gnd_net_),
            .in3(N__38265),
            .lcout(),
            .ltout(\CONTROL.increment28lto5_1_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_2_i_a7_3_LC_17_19_6 .C_ON=1'b0;
    defparam \CONTROL.g0_2_i_a7_3_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_2_i_a7_3_LC_17_19_6 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \CONTROL.g0_2_i_a7_3_LC_17_19_6  (
            .in0(N__38205),
            .in1(N__40819),
            .in2(N__38219),
            .in3(N__48453),
            .lcout(\CONTROL.g0_2_i_a7Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment28lto5_1_2_LC_17_19_7 .C_ON=1'b0;
    defparam \CONTROL.increment28lto5_1_2_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment28lto5_1_2_LC_17_19_7 .LUT_INIT=16'b0001100110011001;
    LogicCell40 \CONTROL.increment28lto5_1_2_LC_17_19_7  (
            .in0(N__72251),
            .in1(N__40818),
            .in2(N__48464),
            .in3(N__38204),
            .lcout(\CONTROL.increment28lto5_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_ne_5_LC_17_20_0 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_ne_5_LC_17_20_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_ne_5_LC_17_20_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \CONTROL.aluOperation_ne_5_LC_17_20_0  (
            .in0(N__44660),
            .in1(N__54582),
            .in2(N__41397),
            .in3(N__44901),
            .lcout(aluOperation_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluOperation_ne_5C_net ),
            .ce(N__38126),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState96_1_i_i_a2_0_1_LC_17_20_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState96_1_i_i_a2_0_1_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState96_1_i_i_a2_0_1_LC_17_20_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \CONTROL.un1_busState96_1_i_i_a2_0_1_LC_17_20_2  (
            .in0(N__41689),
            .in1(N__38584),
            .in2(_gnd_net_),
            .in3(N__55456),
            .lcout(\CONTROL.un1_busState96_1_i_i_a2_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState96_1_i_i_o2_0_LC_17_20_3 .C_ON=1'b0;
    defparam \CONTROL.un1_busState96_1_i_i_o2_0_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState96_1_i_i_o2_0_LC_17_20_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \CONTROL.un1_busState96_1_i_i_o2_0_LC_17_20_3  (
            .in0(N__55455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44658),
            .lcout(\CONTROL.N_140_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_6dflt_LC_17_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_6dflt_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_6dflt_LC_17_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PROM.ROMDATA.dintern_6dflt_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__72273),
            .in2(_gnd_net_),
            .in3(N__55454),
            .lcout(controlWord_6),
            .ltout(controlWord_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState96_1_i_i_a2_1_1_LC_17_20_5 .C_ON=1'b0;
    defparam \CONTROL.un1_busState96_1_i_i_a2_1_1_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState96_1_i_i_a2_1_1_LC_17_20_5 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \CONTROL.un1_busState96_1_i_i_a2_1_1_LC_17_20_5  (
            .in0(N__38583),
            .in1(N__41688),
            .in2(N__38354),
            .in3(N__44659),
            .lcout(),
            .ltout(\CONTROL.un1_busState96_1_i_i_a2_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState96_1_i_i_0_LC_17_20_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState96_1_i_i_0_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState96_1_i_i_0_LC_17_20_6 .LUT_INIT=16'b0011101100111111;
    LogicCell40 \CONTROL.un1_busState96_1_i_i_0_LC_17_20_6  (
            .in0(N__38351),
            .in1(N__54719),
            .in2(N__38345),
            .in3(N__54581),
            .lcout(),
            .ltout(\CONTROL.un1_busState96_1_i_iZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI41SBR02_7_LC_17_20_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI41SBR02_7_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI41SBR02_7_LC_17_20_7 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI41SBR02_7_LC_17_20_7  (
            .in0(N__38330),
            .in1(N__38342),
            .in2(N__38336),
            .in3(N__41117),
            .lcout(\CONTROL.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_5dflt_LC_17_21_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_5dflt_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_5dflt_LC_17_21_0 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \PROM.ROMDATA.dintern_5dflt_LC_17_21_0  (
            .in0(N__47305),
            .in1(N__72272),
            .in2(N__72607),
            .in3(N__64904),
            .lcout(controlWord_5),
            .ltout(controlWord_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState96_1_i_i_o2_LC_17_21_1 .C_ON=1'b0;
    defparam \CONTROL.un1_busState96_1_i_i_o2_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState96_1_i_i_o2_LC_17_21_1 .LUT_INIT=16'b0001001100100011;
    LogicCell40 \CONTROL.un1_busState96_1_i_i_o2_LC_17_21_1  (
            .in0(N__44635),
            .in1(N__54571),
            .in2(N__38333),
            .in3(N__44862),
            .lcout(\CONTROL.N_134_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_LC_17_21_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_LC_17_21_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \CONTROL.un1_busState_0_sqmuxa_i_a2_LC_17_21_2  (
            .in0(N__44769),
            .in1(N__44863),
            .in2(N__38528),
            .in3(N__44636),
            .lcout(\CONTROL.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_2_i_a7_2_LC_17_21_3 .C_ON=1'b0;
    defparam \CONTROL.g0_2_i_a7_2_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_2_i_a7_2_LC_17_21_3 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \CONTROL.g0_2_i_a7_2_LC_17_21_3  (
            .in0(N__53627),
            .in1(N__45401),
            .in2(N__45479),
            .in3(N__54572),
            .lcout(\CONTROL.g0_2_i_a7Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_22_LC_17_21_4 .C_ON=1'b0;
    defparam \CONTROL.g0_22_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_22_LC_17_21_4 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \CONTROL.g0_22_LC_17_21_4  (
            .in0(N__54569),
            .in1(N__71758),
            .in2(_gnd_net_),
            .in3(N__44634),
            .lcout(\CONTROL.N_133_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m126_LC_17_21_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m126_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m126_LC_17_21_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m126_LC_17_21_5  (
            .in0(N__72504),
            .in1(N__64396),
            .in2(_gnd_net_),
            .in3(N__41833),
            .lcout(PROM_ROMDATA_dintern_3ro),
            .ltout(PROM_ROMDATA_dintern_3ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_6_LC_17_21_6 .C_ON=1'b0;
    defparam \CONTROL.g0_6_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_6_LC_17_21_6 .LUT_INIT=16'b0011000000111111;
    LogicCell40 \CONTROL.g0_6_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(N__54568),
            .in2(N__38504),
            .in3(N__44632),
            .lcout(\CONTROL.N_133_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_1_7_LC_17_21_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_1_7_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_1_7_LC_17_21_7 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIO2O5VB_1_7_LC_17_21_7  (
            .in0(N__44633),
            .in1(N__41464),
            .in2(N__71819),
            .in3(N__54570),
            .lcout(\CONTROL.g0_3_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_7_LC_17_22_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_7_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIO2O5VB_7_LC_17_22_0 .LUT_INIT=16'b1011101010111111;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIO2O5VB_7_LC_17_22_0  (
            .in0(N__41463),
            .in1(N__54575),
            .in2(N__71821),
            .in3(N__44649),
            .lcout(),
            .ltout(\CONTROL.g0_2_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI7FBMHV_0_7_LC_17_22_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI7FBMHV_0_7_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI7FBMHV_0_7_LC_17_22_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI7FBMHV_0_7_LC_17_22_1  (
            .in0(N__38486),
            .in1(N__38477),
            .in2(N__38471),
            .in3(N__42149),
            .lcout(\CONTROL.N_5_0 ),
            .ltout(\CONTROL.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNIJQC4JV_1_LC_17_22_2 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNIJQC4JV_1_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNIJQC4JV_1_LC_17_22_2 .LUT_INIT=16'b0011010111110101;
    LogicCell40 \CONTROL.addrstackptr_RNIJQC4JV_1_LC_17_22_2  (
            .in0(N__38468),
            .in1(N__38444),
            .in2(N__38375),
            .in3(N__57820),
            .lcout(\CONTROL.g0_12_1 ),
            .ltout(\CONTROL.g0_12_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNITKBIQ83_2_LC_17_22_3 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNITKBIQ83_2_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNITKBIQ83_2_LC_17_22_3 .LUT_INIT=16'b1000011110001011;
    LogicCell40 \CONTROL.addrstackptr_RNITKBIQ83_2_LC_17_22_3  (
            .in0(N__60682),
            .in1(N__38734),
            .in2(N__38372),
            .in3(N__41958),
            .lcout(\CONTROL.addrstackptr_8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_2dflt_LC_17_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_2dflt_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_2dflt_LC_17_22_4 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \PROM.ROMDATA.dintern_2dflt_LC_17_22_4  (
            .in0(N__41100),
            .in1(N__72261),
            .in2(N__72672),
            .in3(N__41805),
            .lcout(controlWord_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_4dflt_LC_17_22_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_4dflt_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_4dflt_LC_17_22_5 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \PROM.ROMDATA.dintern_4dflt_LC_17_22_5  (
            .in0(N__72260),
            .in1(N__72563),
            .in2(N__54389),
            .in3(N__74138),
            .lcout(controlWord_4),
            .ltout(controlWord_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIQ59BL4_7_LC_17_22_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIQ59BL4_7_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIQ59BL4_7_LC_17_22_6 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIQ59BL4_7_LC_17_22_6  (
            .in0(N__41101),
            .in1(N__72618),
            .in2(N__38738),
            .in3(N__41806),
            .lcout(\CONTROL.N_249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_2_LC_17_22_7 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_2_LC_17_22_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_2_LC_17_22_7 .LUT_INIT=16'b1001001110110001;
    LogicCell40 \CONTROL.addrstackptr_2_LC_17_22_7  (
            .in0(N__38735),
            .in1(N__38723),
            .in2(N__60701),
            .in3(N__41959),
            .lcout(\CONTROL.addrstackptrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.addrstackptr_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_0_LC_17_23_0 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_0_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_0_LC_17_23_0 .LUT_INIT=16'b0111000001110111;
    LogicCell40 \CONTROL.busState_cnst_2_0__m28_0_120_i_i_0_LC_17_23_0  (
            .in0(N__41233),
            .in1(N__38678),
            .in2(N__38810),
            .in3(N__38644),
            .lcout(\CONTROL.m28_0_120_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState97_1_0_a2_LC_17_23_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState97_1_0_a2_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState97_1_0_a2_LC_17_23_2 .LUT_INIT=16'b0000000010001100;
    LogicCell40 \CONTROL.un1_busState97_1_0_a2_LC_17_23_2  (
            .in0(N__44865),
            .in1(N__41581),
            .in2(N__41415),
            .in3(N__41234),
            .lcout(\CONTROL.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_2_LC_17_23_3 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_2_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_2_LC_17_23_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_2_LC_17_23_3  (
            .in0(N__54543),
            .in1(N__41372),
            .in2(N__41670),
            .in3(N__44864),
            .lcout(\CONTROL.N_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment_5_0__m6_i_x2_0_LC_17_23_4 .C_ON=1'b0;
    defparam \CONTROL.increment_5_0__m6_i_x2_0_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment_5_0__m6_i_x2_0_LC_17_23_4 .LUT_INIT=16'b1111000001011010;
    LogicCell40 \CONTROL.increment_5_0__m6_i_x2_0_LC_17_23_4  (
            .in0(N__44638),
            .in1(_gnd_net_),
            .in2(N__41416),
            .in3(N__71806),
            .lcout(\CONTROL.N_114_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m42_LC_17_23_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m42_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m42_LC_17_23_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m42_LC_17_23_5  (
            .in0(N__72511),
            .in1(N__74011),
            .in2(N__45554),
            .in3(N__47702),
            .lcout(PROM_ROMDATA_dintern_0ro),
            .ltout(PROM_ROMDATA_dintern_0ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_0_0_LC_17_23_6 .C_ON=1'b0;
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_0_0_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState_0_sqmuxa_i_a2_0_0_LC_17_23_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \CONTROL.un1_busState_0_sqmuxa_i_a2_0_0_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38531),
            .in3(N__54542),
            .lcout(\CONTROL.un1_busState_0_sqmuxa_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_1_LC_17_23_7 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_1_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_1_LC_17_23_7 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_1_LC_17_23_7  (
            .in0(N__55453),
            .in1(N__41371),
            .in2(N__72320),
            .in3(N__44637),
            .lcout(\CONTROL.N_304_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m433_ns_LC_17_24_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m433_ns_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m433_ns_LC_17_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m433_ns_LC_17_24_0  (
            .in0(N__38744),
            .in1(N__47798),
            .in2(_gnd_net_),
            .in3(N__79845),
            .lcout(\PROM.ROMDATA.m433_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m294_bm_LC_17_24_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m294_bm_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m294_bm_LC_17_24_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m294_bm_LC_17_24_1  (
            .in0(N__78838),
            .in1(N__74129),
            .in2(N__75967),
            .in3(N__78059),
            .lcout(),
            .ltout(\PROM.ROMDATA.m294_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m294_ns_LC_17_24_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m294_ns_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m294_ns_LC_17_24_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m294_ns_LC_17_24_2  (
            .in0(N__41081),
            .in1(_gnd_net_),
            .in2(N__38780),
            .in3(N__76592),
            .lcout(\PROM.ROMDATA.m294_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m31_LC_17_24_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m31_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m31_LC_17_24_3 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m31_LC_17_24_3  (
            .in0(N__78836),
            .in1(N__78055),
            .in2(_gnd_net_),
            .in3(N__77280),
            .lcout(\PROM.ROMDATA.m31 ),
            .ltout(\PROM.ROMDATA.m31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m353_bm_LC_17_24_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m353_bm_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m353_bm_LC_17_24_4 .LUT_INIT=16'b0011001111110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m353_bm_LC_17_24_4  (
            .in0(_gnd_net_),
            .in1(N__41819),
            .in2(N__38777),
            .in3(N__75846),
            .lcout(\PROM.ROMDATA.m353_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_12_LC_17_24_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_12_LC_17_24_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_12_LC_17_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_12_LC_17_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38774),
            .lcout(\CONTROL.dout_reto_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73234),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m391_LC_17_24_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m391_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m391_LC_17_24_6 .LUT_INIT=16'b0000001001000001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m391_LC_17_24_6  (
            .in0(N__77281),
            .in1(N__75847),
            .in2(N__78071),
            .in3(N__78837),
            .lcout(),
            .ltout(\PROM.ROMDATA.m391_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m433_bm_LC_17_24_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m433_bm_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m433_bm_LC_17_24_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m433_bm_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(N__76591),
            .in2(N__38747),
            .in3(N__74246),
            .lcout(\PROM.ROMDATA.m433_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m382_ns_LC_17_25_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m382_ns_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m382_ns_LC_17_25_2 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m382_ns_LC_17_25_2  (
            .in0(N__79342),
            .in1(N__42137),
            .in2(N__47363),
            .in3(N__42119),
            .lcout(\PROM.ROMDATA.m382_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI27KBD_0_LC_18_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNI27KBD_0_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI27KBD_0_LC_18_8_1 .LUT_INIT=16'b1010010100111100;
    LogicCell40 \ALU.d_RNI27KBD_0_LC_18_8_1  (
            .in0(N__39024),
            .in1(N__39089),
            .in2(N__63275),
            .in3(N__53292),
            .lcout(\ALU.d_RNI27KBDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA3Q1H_0_LC_18_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNIA3Q1H_0_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA3Q1H_0_LC_18_8_2 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \ALU.d_RNIA3Q1H_0_LC_18_8_2  (
            .in0(N__53294),
            .in1(N__39100),
            .in2(N__60627),
            .in3(N__39025),
            .lcout(\ALU.N_794_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI6USD6_2_LC_18_8_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI6USD6_2_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI6USD6_2_LC_18_8_4 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \CONTROL.busState_1_RNI6USD6_2_LC_18_8_4  (
            .in0(N__49604),
            .in1(N__50218),
            .in2(N__60626),
            .in3(N__38855),
            .lcout(N_225_0),
            .ltout(N_225_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNISBUGH_14_LC_18_8_5 .C_ON=1'b0;
    defparam \ALU.c_RNISBUGH_14_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNISBUGH_14_LC_18_8_5 .LUT_INIT=16'b0000101010001000;
    LogicCell40 \ALU.c_RNISBUGH_14_LC_18_8_5  (
            .in0(N__63843),
            .in1(N__39091),
            .in2(N__38834),
            .in3(N__53295),
            .lcout(),
            .ltout(\ALU.mult_15_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_371_c_RNIHIRFF5_LC_18_8_6 .C_ON=1'b0;
    defparam \ALU.mult_371_c_RNIHIRFF5_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_371_c_RNIHIRFF5_LC_18_8_6 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \ALU.mult_371_c_RNIHIRFF5_LC_18_8_6  (
            .in0(N__39200),
            .in1(N__38831),
            .in2(N__38825),
            .in3(N__38822),
            .lcout(\ALU.mult_23_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIIRAJH_10_LC_18_8_7 .C_ON=1'b0;
    defparam \ALU.c_RNIIRAJH_10_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIIRAJH_10_LC_18_8_7 .LUT_INIT=16'b0101000011000000;
    LogicCell40 \ALU.c_RNIIRAJH_10_LC_18_8_7  (
            .in0(N__39023),
            .in1(N__39090),
            .in2(N__61715),
            .in3(N__53293),
            .lcout(\ALU.mult_11_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA5S1H_8_LC_18_9_0 .C_ON=1'b0;
    defparam \ALU.d_RNIA5S1H_8_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA5S1H_8_LC_18_9_0 .LUT_INIT=16'b0011000010100000;
    LogicCell40 \ALU.d_RNIA5S1H_8_LC_18_9_0  (
            .in0(N__39095),
            .in1(N__39027),
            .in2(N__62022),
            .in3(N__53296),
            .lcout(\ALU.mult_9_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIRFM5I_11_LC_18_9_2 .C_ON=1'b0;
    defparam \ALU.c_RNIRFM5I_11_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIRFM5I_11_LC_18_9_2 .LUT_INIT=16'b0001111011101000;
    LogicCell40 \ALU.c_RNIRFM5I_11_LC_18_9_2  (
            .in0(N__63112),
            .in1(N__61466),
            .in2(N__74894),
            .in3(N__57046),
            .lcout(\ALU.log_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIKU5GD1_0_14_LC_18_9_4 .C_ON=1'b0;
    defparam \ALU.c_RNIKU5GD1_0_14_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIKU5GD1_0_14_LC_18_9_4 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.c_RNIKU5GD1_0_14_LC_18_9_4  (
            .in0(N__66027),
            .in1(N__63669),
            .in2(N__63853),
            .in3(N__66764),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIR6KVA2_12_LC_18_9_5 .C_ON=1'b0;
    defparam \ALU.c_RNIR6KVA2_12_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIR6KVA2_12_LC_18_9_5 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.c_RNIR6KVA2_12_LC_18_9_5  (
            .in0(N__61012),
            .in1(N__61203),
            .in2(N__39104),
            .in3(N__66028),
            .lcout(\ALU.N_647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI5O9IH_12_LC_18_9_6 .C_ON=1'b0;
    defparam \ALU.c_RNI5O9IH_12_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI5O9IH_12_LC_18_9_6 .LUT_INIT=16'b0011000010100000;
    LogicCell40 \ALU.c_RNI5O9IH_12_LC_18_9_6  (
            .in0(N__39096),
            .in1(N__39026),
            .in2(N__61217),
            .in3(N__53297),
            .lcout(\ALU.mult_13_12 ),
            .ltout(\ALU.mult_13_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_467_c_RNICRDK6B_LC_18_9_7 .C_ON=1'b0;
    defparam \ALU.mult_467_c_RNICRDK6B_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_467_c_RNICRDK6B_LC_18_9_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_467_c_RNICRDK6B_LC_18_9_7  (
            .in0(N__38981),
            .in1(_gnd_net_),
            .in2(N__38960),
            .in3(N__42400),
            .lcout(\ALU.mult_467_c_RNICRDK6BZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_526_c_LC_18_10_0 .C_ON=1'b1;
    defparam \ALU.mult_526_c_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_526_c_LC_18_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_526_c_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__42401),
            .in2(N__38951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\ALU.mult_27_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_526_c_RNIHBG235_LC_18_10_1 .C_ON=1'b1;
    defparam \ALU.mult_526_c_RNIHBG235_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_526_c_RNIHBG235_LC_18_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_526_c_RNIHBG235_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__42386),
            .in2(N__38942),
            .in3(N__38921),
            .lcout(\ALU.mult_27_13 ),
            .ltout(),
            .carryin(\ALU.mult_27_c12 ),
            .carryout(\ALU.mult_27_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_529_c_RNIM6FVL9_LC_18_10_2 .C_ON=1'b1;
    defparam \ALU.mult_529_c_RNIM6FVL9_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_529_c_RNIM6FVL9_LC_18_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_529_c_RNIM6FVL9_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(N__42370),
            .in2(N__38918),
            .in3(N__38900),
            .lcout(\ALU.mult_27_14 ),
            .ltout(),
            .carryin(\ALU.mult_27_c13 ),
            .carryout(\ALU.mult_27_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_27_c14_THRU_LUT4_0_LC_18_10_3 .C_ON=1'b0;
    defparam \ALU.mult_27_c14_THRU_LUT4_0_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_27_c14_THRU_LUT4_0_LC_18_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.mult_27_c14_THRU_LUT4_0_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38897),
            .lcout(\ALU.mult_27_c14_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_546_c_RNIG1E6I8_LC_18_10_4 .C_ON=1'b0;
    defparam \ALU.mult_546_c_RNIG1E6I8_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_546_c_RNIG1E6I8_LC_18_10_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.mult_546_c_RNIG1E6I8_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(N__59144),
            .in2(N__38882),
            .in3(N__40353),
            .lcout(\ALU.mult_546_c_RNIG1E6IZ0Z8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINMQ0E1_10_LC_18_10_5 .C_ON=1'b0;
    defparam \ALU.c_RNINMQ0E1_10_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINMQ0E1_10_LC_18_10_5 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.c_RNINMQ0E1_10_LC_18_10_5  (
            .in0(N__61465),
            .in1(N__65935),
            .in2(N__61716),
            .in3(N__66697),
            .lcout(\ALU.mult_11_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_558_c_RNIB3E8DC_LC_18_10_7 .C_ON=1'b0;
    defparam \ALU.mult_558_c_RNIB3E8DC_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_558_c_RNIB3E8DC_LC_18_10_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \ALU.mult_558_c_RNIB3E8DC_LC_18_10_7  (
            .in0(N__59145),
            .in1(N__39656),
            .in2(_gnd_net_),
            .in3(N__39182),
            .lcout(\ALU.mult_558_c_RNIB3E8DCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFCNKL_9_LC_18_11_1 .C_ON=1'b0;
    defparam \ALU.d_RNIFCNKL_9_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFCNKL_9_LC_18_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIFCNKL_9_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__62818),
            .in2(_gnd_net_),
            .in3(N__68841),
            .lcout(\ALU.d_RNIFCNKLZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIG61LG_9_LC_18_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNIG61LG_9_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIG61LG_9_LC_18_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIG61LG_9_LC_18_11_2  (
            .in0(N__62819),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68439),
            .lcout(\ALU.d_RNIG61LGZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIULN025_0_2_LC_18_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIULN025_0_2_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIULN025_0_2_LC_18_11_3 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \ALU.d_RNIULN025_0_2_LC_18_11_3  (
            .in0(N__68440),
            .in1(N__43599),
            .in2(N__43165),
            .in3(N__68842),
            .lcout(\ALU.d_RNIULN025_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIULN025_2_LC_18_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNIULN025_2_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIULN025_2_LC_18_11_4 .LUT_INIT=16'b0100010011110101;
    LogicCell40 \ALU.d_RNIULN025_2_LC_18_11_4  (
            .in0(N__68843),
            .in1(N__43160),
            .in2(N__43604),
            .in3(N__68441),
            .lcout(),
            .ltout(\ALU.d_RNIULN025Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPTFHMD_2_LC_18_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNIPTFHMD_2_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPTFHMD_2_LC_18_11_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIPTFHMD_2_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__39176),
            .in2(N__39152),
            .in3(N__39149),
            .lcout(),
            .ltout(\ALU.lshift_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIO0KOKE_10_LC_18_11_6 .C_ON=1'b0;
    defparam \ALU.c_RNIO0KOKE_10_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIO0KOKE_10_LC_18_11_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.c_RNIO0KOKE_10_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__70191),
            .in2(N__39143),
            .in3(N__51296),
            .lcout(\ALU.c_RNIO0KOKEZ0Z_10 ),
            .ltout(\ALU.c_RNIO0KOKEZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_10_LC_18_11_7 .C_ON=1'b0;
    defparam \ALU.b_10_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \ALU.b_10_LC_18_11_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.b_10_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__58456),
            .in2(N__39140),
            .in3(N__58283),
            .lcout(\ALU.bZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73143),
            .ce(N__67938),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI8TL4B6_12_LC_18_12_0 .C_ON=1'b0;
    defparam \ALU.c_RNI8TL4B6_12_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI8TL4B6_12_LC_18_12_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNI8TL4B6_12_LC_18_12_0  (
            .in0(N__42787),
            .in1(N__42794),
            .in2(_gnd_net_),
            .in3(N__39188),
            .lcout(\ALU.N_1025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIHOSI72_12_LC_18_12_1 .C_ON=1'b0;
    defparam \ALU.c_RNIHOSI72_12_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIHOSI72_12_LC_18_12_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNIHOSI72_12_LC_18_12_1  (
            .in0(N__65903),
            .in1(N__42811),
            .in2(_gnd_net_),
            .in3(N__42788),
            .lcout(),
            .ltout(\ALU.N_965_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFHCRU4_2_LC_18_12_2 .C_ON=1'b0;
    defparam \ALU.d_RNIFHCRU4_2_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFHCRU4_2_LC_18_12_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.d_RNIFHCRU4_2_LC_18_12_2  (
            .in0(N__39233),
            .in1(_gnd_net_),
            .in2(N__39212),
            .in3(N__68920),
            .lcout(\ALU.d_RNIFHCRU4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBN2FN8_11_LC_18_12_4 .C_ON=1'b0;
    defparam \ALU.c_RNIBN2FN8_11_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBN2FN8_11_LC_18_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIBN2FN8_11_LC_18_12_4  (
            .in0(N__70187),
            .in1(N__51322),
            .in2(_gnd_net_),
            .in3(N__42821),
            .lcout(\ALU.c_RNIBN2FN8Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINMQ0E1_0_10_LC_18_12_5 .C_ON=1'b0;
    defparam \ALU.c_RNINMQ0E1_0_10_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINMQ0E1_0_10_LC_18_12_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.c_RNINMQ0E1_0_10_LC_18_12_5  (
            .in0(N__61439),
            .in1(N__65904),
            .in2(N__61717),
            .in3(N__66699),
            .lcout(\ALU.lshift_3_ns_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIKU5GD1_14_LC_18_12_6 .C_ON=1'b0;
    defparam \ALU.c_RNIKU5GD1_14_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIKU5GD1_14_LC_18_12_6 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.c_RNIKU5GD1_14_LC_18_12_6  (
            .in0(N__66698),
            .in1(N__63644),
            .in2(N__63842),
            .in3(N__65902),
            .lcout(\ALU.mult_15_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINT9PO2_10_LC_18_12_7 .C_ON=1'b0;
    defparam \ALU.c_RNINT9PO2_10_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINT9PO2_10_LC_18_12_7 .LUT_INIT=16'b0101010111100100;
    LogicCell40 \ALU.c_RNINT9PO2_10_LC_18_12_7  (
            .in0(N__68919),
            .in1(N__42810),
            .in2(N__62656),
            .in3(N__65905),
            .lcout(\ALU.c_RNINT9PO2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI61KC1_13_LC_18_13_0 .C_ON=1'b0;
    defparam \ALU.b_RNI61KC1_13_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI61KC1_13_LC_18_13_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.b_RNI61KC1_13_LC_18_13_0  (
            .in0(N__51541),
            .in1(N__57631),
            .in2(_gnd_net_),
            .in3(N__43295),
            .lcout(\ALU.b_RNI61KC1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAHCT_13_LC_18_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIAHCT_13_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAHCT_13_LC_18_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIAHCT_13_LC_18_13_1  (
            .in0(N__43294),
            .in1(N__57891),
            .in2(_gnd_net_),
            .in3(N__65060),
            .lcout(\ALU.d_RNIAHCTZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI890L_13_LC_18_13_2 .C_ON=1'b0;
    defparam \ALU.c_RNI890L_13_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI890L_13_LC_18_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNI890L_13_LC_18_13_2  (
            .in0(N__52350),
            .in1(N__67348),
            .in2(_gnd_net_),
            .in3(N__43293),
            .lcout(\ALU.c_RNI890LZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI4P741_13_LC_18_13_3 .C_ON=1'b0;
    defparam \ALU.a_RNI4P741_13_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI4P741_13_LC_18_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_RNI4P741_13_LC_18_13_3  (
            .in0(N__43296),
            .in1(N__52477),
            .in2(_gnd_net_),
            .in3(N__57170),
            .lcout(),
            .ltout(\ALU.a_RNI4P741Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNILN2L2_13_LC_18_13_4 .C_ON=1'b0;
    defparam \ALU.c_RNILN2L2_13_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNILN2L2_13_LC_18_13_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.c_RNILN2L2_13_LC_18_13_4  (
            .in0(N__39698),
            .in1(N__53951),
            .in2(N__39692),
            .in3(N__46811),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9K0D5_13_LC_18_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNI9K0D5_13_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9K0D5_13_LC_18_13_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI9K0D5_13_LC_18_13_5  (
            .in0(N__53952),
            .in1(N__39689),
            .in2(N__39683),
            .in3(N__39680),
            .lcout(\ALU.operand2_13 ),
            .ltout(\ALU.operand2_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINGV4G_13_LC_18_13_6 .C_ON=1'b0;
    defparam \ALU.d_RNINGV4G_13_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINGV4G_13_LC_18_13_6 .LUT_INIT=16'b0011001111110000;
    LogicCell40 \ALU.d_RNINGV4G_13_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__39652),
            .in2(N__39614),
            .in3(N__71467),
            .lcout(\ALU.N_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJAJOO_10_LC_18_13_7 .C_ON=1'b0;
    defparam \ALU.c_RNIJAJOO_10_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJAJOO_10_LC_18_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIJAJOO_10_LC_18_13_7  (
            .in0(N__61697),
            .in1(N__62811),
            .in2(_gnd_net_),
            .in3(N__66721),
            .lcout(\ALU.N_837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_2_LC_18_14_0 .C_ON=1'b0;
    defparam \ALU.b_2_LC_18_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.b_2_LC_18_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.b_2_LC_18_14_0  (
            .in0(N__39606),
            .in1(N__39535),
            .in2(_gnd_net_),
            .in3(N__39468),
            .lcout(\ALU.bZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73155),
            .ce(N__67943),
            .sr(_gnd_net_));
    defparam \ALU.b_4_LC_18_14_1 .C_ON=1'b0;
    defparam \ALU.b_4_LC_18_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.b_4_LC_18_14_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.b_4_LC_18_14_1  (
            .in0(N__42529),
            .in1(N__57350),
            .in2(_gnd_net_),
            .in3(N__39395),
            .lcout(\ALU.bZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73155),
            .ce(N__67943),
            .sr(_gnd_net_));
    defparam \ALU.b_5_LC_18_14_2 .C_ON=1'b0;
    defparam \ALU.b_5_LC_18_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.b_5_LC_18_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_5_LC_18_14_2  (
            .in0(N__57349),
            .in1(N__52619),
            .in2(_gnd_net_),
            .in3(N__39320),
            .lcout(\ALU.bZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73155),
            .ce(N__67943),
            .sr(_gnd_net_));
    defparam \ALU.b_6_LC_18_14_3 .C_ON=1'b0;
    defparam \ALU.b_6_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.b_6_LC_18_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_6_LC_18_14_3  (
            .in0(N__43040),
            .in1(N__43086),
            .in2(_gnd_net_),
            .in3(N__42977),
            .lcout(\ALU.bZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73155),
            .ce(N__67943),
            .sr(_gnd_net_));
    defparam \ALU.b_3_LC_18_14_4 .C_ON=1'b0;
    defparam \ALU.b_3_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.b_3_LC_18_14_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.b_3_LC_18_14_4  (
            .in0(N__58812),
            .in1(N__58745),
            .in2(_gnd_net_),
            .in3(N__58678),
            .lcout(\ALU.bZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73155),
            .ce(N__67943),
            .sr(_gnd_net_));
    defparam \ALU.b_11_LC_18_14_5 .C_ON=1'b0;
    defparam \ALU.b_11_LC_18_14_5 .SEQ_MODE=4'b1000;
    defparam \ALU.b_11_LC_18_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.b_11_LC_18_14_5  (
            .in0(N__58184),
            .in1(N__58108),
            .in2(_gnd_net_),
            .in3(N__58050),
            .lcout(\ALU.bZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73155),
            .ce(N__67943),
            .sr(_gnd_net_));
    defparam \ALU.b_12_LC_18_14_6 .C_ON=1'b0;
    defparam \ALU.b_12_LC_18_14_6 .SEQ_MODE=4'b1000;
    defparam \ALU.b_12_LC_18_14_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \ALU.b_12_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__67757),
            .in2(N__67622),
            .in3(N__67691),
            .lcout(\ALU.bZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73155),
            .ce(N__67943),
            .sr(_gnd_net_));
    defparam \CONTROL.g3_LC_18_14_7 .C_ON=1'b0;
    defparam \CONTROL.g3_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g3_LC_18_14_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \CONTROL.g3_LC_18_14_7  (
            .in0(N__53720),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53668),
            .lcout(\CONTROL.gZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDC6LJ1_2_LC_18_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNIDC6LJ1_2_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDC6LJ1_2_LC_18_15_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ALU.d_RNIDC6LJ1_2_LC_18_15_0  (
            .in0(N__65957),
            .in1(N__39764),
            .in2(_gnd_net_),
            .in3(N__68515),
            .lcout(\ALU.lshift_15_0_1 ),
            .ltout(\ALU.lshift_15_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNITNPJL2_14_LC_18_15_1 .C_ON=1'b0;
    defparam \ALU.c_RNITNPJL2_14_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNITNPJL2_14_LC_18_15_1 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \ALU.c_RNITNPJL2_14_LC_18_15_1  (
            .in0(N__39732),
            .in1(N__69928),
            .in2(N__39707),
            .in3(N__39704),
            .lcout(\ALU.a_15_m0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI6KIQO_14_LC_18_15_2 .C_ON=1'b0;
    defparam \ALU.c_RNI6KIQO_14_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI6KIQO_14_LC_18_15_2 .LUT_INIT=16'b0011000001010000;
    LogicCell40 \ALU.c_RNI6KIQO_14_LC_18_15_2  (
            .in0(N__63802),
            .in1(N__63668),
            .in2(N__69965),
            .in3(N__66682),
            .lcout(\ALU.a_15_m0_sx_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI34ECO_9_LC_18_15_3 .C_ON=1'b0;
    defparam \ALU.d_RNI34ECO_9_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI34ECO_9_LC_18_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI34ECO_9_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__62764),
            .in2(_gnd_net_),
            .in3(N__65955),
            .lcout(\ALU.d_RNI34ECOZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9QA4D1_0_LC_18_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNI9QA4D1_0_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9QA4D1_0_LC_18_15_4 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.d_RNI9QA4D1_0_LC_18_15_4  (
            .in0(N__65958),
            .in1(N__60568),
            .in2(N__65575),
            .in3(N__66683),
            .lcout(),
            .ltout(\ALU.mult_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI05SGP3_0_LC_18_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNI05SGP3_0_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI05SGP3_0_LC_18_15_5 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.d_RNI05SGP3_0_LC_18_15_5  (
            .in0(N__59066),
            .in1(N__40184),
            .in2(N__40178),
            .in3(N__47986),
            .lcout(\ALU.a_15_m3_d_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJOQE21_0_LC_18_15_6 .C_ON=1'b0;
    defparam \ALU.d_RNIJOQE21_0_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJOQE21_0_LC_18_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIJOQE21_0_LC_18_15_6  (
            .in0(N__65569),
            .in1(N__60567),
            .in2(N__56141),
            .in3(N__55875),
            .lcout(\ALU.d_RNIJOQE21Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_293_c_RNO_LC_18_15_7 .C_ON=1'b0;
    defparam \ALU.mult_293_c_RNO_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_293_c_RNO_LC_18_15_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_293_c_RNO_LC_18_15_7  (
            .in0(N__66684),
            .in1(N__62765),
            .in2(N__61982),
            .in3(N__65956),
            .lcout(\ALU.mult_293_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI8KVQ_5_LC_18_16_0 .C_ON=1'b0;
    defparam \ALU.c_RNI8KVQ_5_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI8KVQ_5_LC_18_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNI8KVQ_5_LC_18_16_0  (
            .in0(N__40134),
            .in1(N__40090),
            .in2(_gnd_net_),
            .in3(N__43974),
            .lcout(\ALU.c_RNI8KVQZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI48JM_5_LC_18_16_1 .C_ON=1'b0;
    defparam \ALU.e_RNI48JM_5_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI48JM_5_LC_18_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_RNI48JM_5_LC_18_16_1  (
            .in0(N__43975),
            .in1(N__40069),
            .in2(_gnd_net_),
            .in3(N__40043),
            .lcout(),
            .ltout(\ALU.e_RNI48JMZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNILHDD2_5_LC_18_16_2 .C_ON=1'b0;
    defparam \ALU.e_RNILHDD2_5_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNILHDD2_5_LC_18_16_2 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \ALU.e_RNILHDD2_5_LC_18_16_2  (
            .in0(N__53887),
            .in1(N__40013),
            .in2(N__40007),
            .in3(N__46779),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBAG34_5_LC_18_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNIBAG34_5_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBAG34_5_LC_18_16_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIBAG34_5_LC_18_16_3  (
            .in0(N__40196),
            .in1(N__39905),
            .in2(N__40004),
            .in3(N__53888),
            .lcout(\ALU.operand2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI7HSP_5_LC_18_16_4 .C_ON=1'b0;
    defparam \ALU.b_RNI7HSP_5_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI7HSP_5_LC_18_16_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ALU.b_RNI7HSP_5_LC_18_16_4  (
            .in0(N__39973),
            .in1(_gnd_net_),
            .in2(N__46922),
            .in3(N__39922),
            .lcout(\ALU.b_RNI7HSPZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBT8E_5_LC_18_16_5 .C_ON=1'b0;
    defparam \ALU.d_RNIBT8E_5_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBT8E_5_LC_18_16_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIBT8E_5_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__46892),
            .in2(N__40267),
            .in3(N__40219),
            .lcout(\ALU.d_RNIBT8EZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_2_rep1_ne_LC_18_16_6 .C_ON=1'b0;
    defparam \CONTROL.operand2_2_rep1_ne_LC_18_16_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_2_rep1_ne_LC_18_16_6 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \CONTROL.operand2_2_rep1_ne_LC_18_16_6  (
            .in0(N__79411),
            .in1(N__40916),
            .in2(N__40298),
            .in3(N__44495),
            .lcout(aluOperand2_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_2_rep1_neC_net ),
            .ce(N__40657),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_2_rep2_ne_LC_18_16_7 .C_ON=1'b0;
    defparam \CONTROL.operand2_2_rep2_ne_LC_18_16_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_2_rep2_ne_LC_18_16_7 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \CONTROL.operand2_2_rep2_ne_LC_18_16_7  (
            .in0(N__44496),
            .in1(N__40292),
            .in2(N__40924),
            .in3(N__79412),
            .lcout(aluOperand2_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_2_rep1_neC_net ),
            .ce(N__40657),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m407_LC_18_17_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m407_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m407_LC_18_17_0 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m407_LC_18_17_0  (
            .in0(N__74492),
            .in1(N__76583),
            .in2(N__45805),
            .in3(N__75815),
            .lcout(),
            .ltout(\PROM.ROMDATA.m407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m418_ns_1_LC_18_17_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m418_ns_1_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m418_ns_1_LC_18_17_1 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m418_ns_1_LC_18_17_1  (
            .in0(N__79879),
            .in1(N__40796),
            .in2(N__40190),
            .in3(N__72727),
            .lcout(\PROM.ROMDATA.m418_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m134_LC_18_17_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m134_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m134_LC_18_17_2 .LUT_INIT=16'b0101010110011001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m134_LC_18_17_2  (
            .in0(N__78851),
            .in1(N__78050),
            .in2(_gnd_net_),
            .in3(N__77312),
            .lcout(\PROM.ROMDATA.m134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_fast_ne_1_LC_18_17_3 .C_ON=1'b0;
    defparam \CONTROL.operand2_fast_ne_1_LC_18_17_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_fast_ne_1_LC_18_17_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \CONTROL.operand2_fast_ne_1_LC_18_17_3  (
            .in0(N__79880),
            .in1(N__40800),
            .in2(N__79495),
            .in3(N__72729),
            .lcout(aluOperand2_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_fast_ne_1C_net ),
            .ce(N__40658),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_1_rep1_ne_LC_18_17_4 .C_ON=1'b0;
    defparam \CONTROL.operand2_1_rep1_ne_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_1_rep1_ne_LC_18_17_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \CONTROL.operand2_1_rep1_ne_LC_18_17_4  (
            .in0(N__72728),
            .in1(N__79433),
            .in2(N__40802),
            .in3(N__79882),
            .lcout(aluOperand2_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_fast_ne_1C_net ),
            .ce(N__40658),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m488_ns_LC_18_17_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m488_ns_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m488_ns_LC_18_17_5 .LUT_INIT=16'b0100000100011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m488_ns_LC_18_17_5  (
            .in0(N__77313),
            .in1(N__74087),
            .in2(N__78070),
            .in3(N__78852),
            .lcout(),
            .ltout(\PROM.ROMDATA.m488_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m500_ns_1_LC_18_17_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m500_ns_1_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m500_ns_1_LC_18_17_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m500_ns_1_LC_18_17_6  (
            .in0(N__64298),
            .in1(N__79432),
            .in2(N__40187),
            .in3(N__79878),
            .lcout(\PROM.ROMDATA.m500_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_ne_1_LC_18_17_7 .C_ON=1'b0;
    defparam \CONTROL.operand2_ne_1_LC_18_17_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_ne_1_LC_18_17_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \CONTROL.operand2_ne_1_LC_18_17_7  (
            .in0(N__79881),
            .in1(N__40801),
            .in2(N__79496),
            .in3(N__72730),
            .lcout(aluOperand2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.operand2_fast_ne_1C_net ),
            .ce(N__40658),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJP1AE_0_9_LC_18_18_1 .C_ON=1'b0;
    defparam \ALU.d_RNIJP1AE_0_9_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJP1AE_0_9_LC_18_18_1 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \ALU.d_RNIJP1AE_0_9_LC_18_18_1  (
            .in0(N__40601),
            .in1(N__40541),
            .in2(N__40499),
            .in3(N__40513),
            .lcout(\ALU.combOperand2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI27JA5_1_LC_18_18_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI27JA5_1_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI27JA5_1_LC_18_18_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \CONTROL.busState_1_RNI27JA5_1_LC_18_18_3  (
            .in0(N__50156),
            .in1(N__40498),
            .in2(N__62886),
            .in3(N__50342),
            .lcout(\CONTROL.N_202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_RNIEUOJ_9_LC_18_18_4 .C_ON=1'b0;
    defparam \CONTROL.dout_RNIEUOJ_9_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.dout_RNIEUOJ_9_LC_18_18_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.dout_RNIEUOJ_9_LC_18_18_4  (
            .in0(N__40463),
            .in1(N__40309),
            .in2(_gnd_net_),
            .in3(N__50154),
            .lcout(),
            .ltout(\CONTROL.N_170_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIDRGO1_2_LC_18_18_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIDRGO1_2_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIDRGO1_2_LC_18_18_5 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \CONTROL.busState_1_RNIDRGO1_2_LC_18_18_5  (
            .in0(N__50155),
            .in1(N__40433),
            .in2(N__40403),
            .in3(N__49575),
            .lcout(N_186),
            .ltout(N_186_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNILFVQ7_0_LC_18_18_6 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNILFVQ7_0_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNILFVQ7_0_LC_18_18_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \CONTROL.busState_1_RNILFVQ7_0_LC_18_18_6  (
            .in0(N__49576),
            .in1(N__40394),
            .in2(N__40388),
            .in3(N__49818),
            .lcout(bus_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_9_LC_18_18_7 .C_ON=1'b0;
    defparam \CONTROL.dout_9_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_9_LC_18_18_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \CONTROL.dout_9_LC_18_18_7  (
            .in0(N__72300),
            .in1(N__72380),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.ctrlOut_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_9C_net ),
            .ce(N__44398),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m284_LC_18_19_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m284_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m284_LC_18_19_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m284_LC_18_19_0  (
            .in0(N__50759),
            .in1(N__43714),
            .in2(N__79861),
            .in3(N__78956),
            .lcout(\PROM.ROMDATA.m284 ),
            .ltout(\PROM.ROMDATA.m284_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_12dflt_LC_18_19_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_12dflt_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_12dflt_LC_18_19_1 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \PROM.ROMDATA.dintern_12dflt_LC_18_19_1  (
            .in0(N__79298),
            .in1(N__40913),
            .in2(N__40832),
            .in3(N__44478),
            .lcout(controlWord_12),
            .ltout(controlWord_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment28lto5_0_ns_LC_18_19_2 .C_ON=1'b0;
    defparam \CONTROL.increment28lto5_0_ns_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment28lto5_0_ns_LC_18_19_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \CONTROL.increment28lto5_0_ns_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__40775),
            .in2(N__40829),
            .in3(N__40769),
            .lcout(\CONTROL.increment28lto5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m273_LC_18_19_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m273_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m273_LC_18_19_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m273_LC_18_19_3  (
            .in0(N__78955),
            .in1(N__75619),
            .in2(N__76619),
            .in3(N__78753),
            .lcout(\PROM.ROMDATA.m273 ),
            .ltout(\PROM.ROMDATA.m273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m276_LC_18_19_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m276_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m276_LC_18_19_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m276_LC_18_19_4  (
            .in0(N__72683),
            .in1(N__79297),
            .in2(N__40781),
            .in3(N__79783),
            .lcout(PROM_ROMDATA_dintern_11ro),
            .ltout(PROM_ROMDATA_dintern_11ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment28lto5_0_x1_LC_18_19_5 .C_ON=1'b0;
    defparam \CONTROL.increment28lto5_0_x1_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment28lto5_0_x1_LC_18_19_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \CONTROL.increment28lto5_0_x1_LC_18_19_5  (
            .in0(N__72249),
            .in1(N__40750),
            .in2(N__40778),
            .in3(N__56656),
            .lcout(\CONTROL.increment28lto5_0_xZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment28lto5_0_x0_LC_18_19_6 .C_ON=1'b0;
    defparam \CONTROL.increment28lto5_0_x0_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment28lto5_0_x0_LC_18_19_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \CONTROL.increment28lto5_0_x0_LC_18_19_6  (
            .in0(N__40749),
            .in1(N__72250),
            .in2(_gnd_net_),
            .in3(N__40762),
            .lcout(\CONTROL.increment28lto5_0_xZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_1_i_a6_0_LC_18_19_7 .C_ON=1'b0;
    defparam \CONTROL.g0_1_i_a6_0_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_1_i_a6_0_LC_18_19_7 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \CONTROL.g0_1_i_a6_0_LC_18_19_7  (
            .in0(N__40763),
            .in1(N__56657),
            .in2(N__40754),
            .in3(N__40715),
            .lcout(\CONTROL.g0_1_i_a6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_1_i_a6_1_LC_18_20_0 .C_ON=1'b0;
    defparam \CONTROL.g0_1_i_a6_1_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_1_i_a6_1_LC_18_20_0 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \CONTROL.g0_1_i_a6_1_LC_18_20_0  (
            .in0(N__53662),
            .in1(N__45509),
            .in2(N__53717),
            .in3(N__45392),
            .lcout(\CONTROL.g0_1_i_a6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_a7_0_LC_18_20_1 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_a7_0_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_a7_0_LC_18_20_1 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \CONTROL.g0_3_i_a7_0_LC_18_20_1  (
            .in0(N__45391),
            .in1(N__53705),
            .in2(N__45516),
            .in3(N__53661),
            .lcout(\CONTROL.g0_3_i_a7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m271_1_LC_18_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m271_1_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m271_1_LC_18_20_2 .LUT_INIT=16'b0011010111110101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m271_1_LC_18_20_2  (
            .in0(N__79210),
            .in1(N__47524),
            .in2(N__72726),
            .in3(N__47537),
            .lcout(\PROM.ROMDATA.m271_1 ),
            .ltout(\PROM.ROMDATA.m271_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m271_LC_18_20_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m271_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m271_LC_18_20_3 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m271_LC_18_20_3  (
            .in0(N__72655),
            .in1(N__44920),
            .in2(N__41057),
            .in3(N__50713),
            .lcout(PROM_ROMDATA_dintern_10ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m258_ns_LC_18_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m258_ns_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m258_ns_LC_18_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m258_ns_LC_18_20_4  (
            .in0(N__79818),
            .in1(N__45194),
            .in2(_gnd_net_),
            .in3(N__45356),
            .lcout(\PROM.ROMDATA.m258_ns ),
            .ltout(\PROM.ROMDATA.m258_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m260_LC_18_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m260_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m260_LC_18_20_5 .LUT_INIT=16'b0111011000110010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m260_LC_18_20_5  (
            .in0(N__72656),
            .in1(N__45031),
            .in2(N__41024),
            .in3(N__50470),
            .lcout(PROM_ROMDATA_dintern_9ro),
            .ltout(PROM_ROMDATA_dintern_9ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment28lto5_1_0_LC_18_20_6 .C_ON=1'b0;
    defparam \CONTROL.increment28lto5_1_0_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.increment28lto5_1_0_LC_18_20_6 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \CONTROL.increment28lto5_1_0_LC_18_20_6  (
            .in0(N__53704),
            .in1(N__45505),
            .in2(N__41021),
            .in3(N__45390),
            .lcout(\CONTROL.increment28lto5_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m404_LC_18_20_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m404_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m404_LC_18_20_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m404_LC_18_20_7  (
            .in0(N__79299),
            .in1(N__64246),
            .in2(N__47528),
            .in3(N__75708),
            .lcout(\PROM.ROMDATA.N_566_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m470_bm_LC_18_21_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m470_bm_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m470_bm_LC_18_21_0 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m470_bm_LC_18_21_0  (
            .in0(N__64245),
            .in1(N__76470),
            .in2(N__69359),
            .in3(N__75598),
            .lcout(\PROM.ROMDATA.m470_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_RNO_0_6_LC_18_21_1 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_RNO_0_6_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_RNO_0_6_LC_18_21_1 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \CONTROL.aluOperation_RNO_0_6_LC_18_21_1  (
            .in0(N__41194),
            .in1(N__54766),
            .in2(N__40967),
            .in3(N__41559),
            .lcout(\CONTROL.aluOperation_12_i_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState97_i_i_o2_LC_18_21_2 .C_ON=1'b0;
    defparam \CONTROL.un1_busState97_i_i_o2_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState97_i_i_o2_LC_18_21_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \CONTROL.un1_busState97_i_i_o2_LC_18_21_2  (
            .in0(N__41558),
            .in1(N__41192),
            .in2(N__41395),
            .in3(N__44903),
            .lcout(\CONTROL.N_86_0 ),
            .ltout(\CONTROL.N_86_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_cnst_2_0__m38_i_m2_LC_18_21_3 .C_ON=1'b0;
    defparam \CONTROL.busState_cnst_2_0__m38_i_m2_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_cnst_2_0__m38_i_m2_LC_18_21_3 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \CONTROL.busState_cnst_2_0__m38_i_m2_LC_18_21_3  (
            .in0(N__41193),
            .in1(_gnd_net_),
            .in2(N__41705),
            .in3(N__41697),
            .lcout(\CONTROL.N_135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m444_am_LC_18_21_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m444_am_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m444_am_LC_18_21_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m444_am_LC_18_21_4  (
            .in0(N__64870),
            .in1(N__78712),
            .in2(_gnd_net_),
            .in3(N__75597),
            .lcout(\PROM.ROMDATA.m444_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_7_f0_163_0_o2_LC_18_21_5 .C_ON=1'b0;
    defparam \CONTROL.aluParams_7_f0_163_0_o2_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluParams_7_f0_163_0_o2_LC_18_21_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \CONTROL.aluParams_7_f0_163_0_o2_LC_18_21_5  (
            .in0(_gnd_net_),
            .in1(N__54544),
            .in2(_gnd_net_),
            .in3(N__44631),
            .lcout(\CONTROL.N_74_0 ),
            .ltout(\CONTROL.N_74_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIUBNO8E_7_LC_18_21_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIUBNO8E_7_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIUBNO8E_7_LC_18_21_6 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIUBNO8E_7_LC_18_21_6  (
            .in0(N__41476),
            .in1(N__41391),
            .in2(N__41264),
            .in3(N__44902),
            .lcout(),
            .ltout(\CONTROL.un1_busState96_1_i_i_232_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNINU4NAR_7_LC_18_21_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNINU4NAR_7_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNINU4NAR_7_LC_18_21_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNINU4NAR_7_LC_18_21_7  (
            .in0(N__41191),
            .in1(_gnd_net_),
            .in2(N__41120),
            .in3(N__47002),
            .lcout(\CONTROL.programCounter_ret_36_RNINU4NARZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_RNIT3IG_5_LC_18_22_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_RNIT3IG_5_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_19_RNIT3IG_5_LC_18_22_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \CONTROL.programCounter_ret_19_RNIT3IG_5_LC_18_22_0  (
            .in0(N__45658),
            .in1(N__64595),
            .in2(_gnd_net_),
            .in3(N__41764),
            .lcout(\CONTROL.programCounter_ret_19_RNIT3IGZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m23_LC_18_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m23_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m23_LC_18_22_1 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m23_LC_18_22_1  (
            .in0(N__77865),
            .in1(_gnd_net_),
            .in2(N__78845),
            .in3(N__77182),
            .lcout(\PROM.ROMDATA.m23 ),
            .ltout(\PROM.ROMDATA.m23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m97_LC_18_22_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m97_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m97_LC_18_22_2 .LUT_INIT=16'b1000100000001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m97_LC_18_22_2  (
            .in0(N__73997),
            .in1(N__73491),
            .in2(N__41111),
            .in3(N__75852),
            .lcout(PROM_ROMDATA_dintern_31_0__N_556_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m294_am_LC_18_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m294_am_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m294_am_LC_18_22_3 .LUT_INIT=16'b1000000001001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m294_am_LC_18_22_3  (
            .in0(N__77866),
            .in1(N__78787),
            .in2(N__75968),
            .in3(N__77183),
            .lcout(\PROM.ROMDATA.m294_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m16_LC_18_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m16_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m16_LC_18_22_4 .LUT_INIT=16'b0011010100000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m16_LC_18_22_4  (
            .in0(N__73572),
            .in1(N__73808),
            .in2(N__73719),
            .in3(N__77863),
            .lcout(\PROM.ROMDATA.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m125_e_LC_18_22_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m125_e_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m125_e_LC_18_22_5 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m125_e_LC_18_22_5  (
            .in0(N__79142),
            .in1(N__79613),
            .in2(N__76462),
            .in3(_gnd_net_),
            .lcout(m125_e),
            .ltout(m125_e_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m125_LC_18_22_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m125_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m125_LC_18_22_6 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m125_LC_18_22_6  (
            .in0(N__41846),
            .in1(N__50572),
            .in2(N__41837),
            .in3(N__75851),
            .lcout(\PROM.ROMDATA.N_557_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m77_LC_18_22_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m77_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m77_LC_18_22_7 .LUT_INIT=16'b0000101001011010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m77_LC_18_22_7  (
            .in0(N__77864),
            .in1(_gnd_net_),
            .in2(N__78844),
            .in3(N__77181),
            .lcout(\PROM.ROMDATA.m77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m93_ns_LC_18_23_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m93_ns_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m93_ns_LC_18_23_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m93_ns_LC_18_23_0  (
            .in0(N__54968),
            .in1(N__51107),
            .in2(N__79417),
            .in3(N__51047),
            .lcout(m93_ns),
            .ltout(m93_ns_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNI257R22_7_LC_18_23_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNI257R22_7_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNI257R22_7_LC_18_23_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNI257R22_7_LC_18_23_1  (
            .in0(N__74007),
            .in1(N__50561),
            .in2(N__41792),
            .in3(N__72695),
            .lcout(\CONTROL.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_5_LC_18_23_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_5_LC_18_23_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_5_LC_18_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_5_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41789),
            .lcout(\CONTROL.addrstack_reto_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73235),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI4MHF_5_LC_18_23_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI4MHF_5_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI4MHF_5_LC_18_23_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI4MHF_5_LC_18_23_3  (
            .in0(N__41716),
            .in1(N__64594),
            .in2(_gnd_net_),
            .in3(N__41763),
            .lcout(\CONTROL.programCounter_ret_1_RNI4MHFZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_5_LC_18_23_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_5_LC_18_23_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_5_LC_18_23_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_5_LC_18_23_4  (
            .in0(N__41747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73235),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_35_rep2_LC_18_23_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_35_rep2_LC_18_23_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_35_rep2_LC_18_23_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \CONTROL.programCounter_ret_35_rep2_LC_18_23_5  (
            .in0(N__50872),
            .in1(_gnd_net_),
            .in2(N__50842),
            .in3(_gnd_net_),
            .lcout(CONTROL_programCounter11_reto_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73235),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_rep1_LC_18_23_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_rep1_LC_18_23_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_18_rep1_LC_18_23_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CONTROL.programCounter_ret_18_rep1_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(N__50830),
            .in2(_gnd_net_),
            .in3(N__50871),
            .lcout(\CONTROL.un1_programCounter9_reto_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73235),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m48_LC_18_23_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m48_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m48_LC_18_23_7 .LUT_INIT=16'b0100000110010101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m48_LC_18_23_7  (
            .in0(N__78746),
            .in1(N__77995),
            .in2(N__75966),
            .in3(N__77258),
            .lcout(\PROM.ROMDATA.m48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_2_1_LC_18_24_0 .C_ON=1'b0;
    defparam \CONTROL.g0_2_1_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_2_1_LC_18_24_0 .LUT_INIT=16'b1111011101111111;
    LogicCell40 \CONTROL.g0_2_1_LC_18_24_0  (
            .in0(N__55421),
            .in1(N__72307),
            .in2(N__42262),
            .in3(N__54633),
            .lcout(\CONTROL.g0_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_4_2_LC_18_24_1 .C_ON=1'b0;
    defparam \CONTROL.g0_4_2_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_4_2_LC_18_24_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \CONTROL.g0_4_2_LC_18_24_1  (
            .in0(N__72311),
            .in1(N__42026),
            .in2(_gnd_net_),
            .in3(N__55423),
            .lcout(\CONTROL.g0_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment_0_LC_18_24_2 .C_ON=1'b0;
    defparam \CONTROL.increment_0_LC_18_24_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.increment_0_LC_18_24_2 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \CONTROL.increment_0_LC_18_24_2  (
            .in0(N__47010),
            .in1(N__42017),
            .in2(N__44713),
            .in3(N__47050),
            .lcout(\CONTROL.incrementZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.increment_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNIF0HGO91_7_LC_18_24_3 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNIF0HGO91_7_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNIF0HGO91_7_LC_18_24_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \CONTROL.addrstackptr_RNIF0HGO91_7_LC_18_24_3  (
            .in0(N__60653),
            .in1(N__42280),
            .in2(N__42011),
            .in3(N__41976),
            .lcout(\CONTROL.g1_1 ),
            .ltout(\CONTROL.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNIF61SK42_7_LC_18_24_4 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNIF61SK42_7_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNIF61SK42_7_LC_18_24_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.addrstackptr_RNIF61SK42_7_LC_18_24_4  (
            .in0(N__42334),
            .in1(N__42304),
            .in2(N__41888),
            .in3(N__41852),
            .lcout(\CONTROL.addrstackptr_N_7_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIEO2I4H_7_LC_18_24_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIEO2I4H_7_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIEO2I4H_7_LC_18_24_5 .LUT_INIT=16'b0000001001000110;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIEO2I4H_7_LC_18_24_5  (
            .in0(N__54635),
            .in1(N__42249),
            .in2(N__41864),
            .in3(N__47009),
            .lcout(\CONTROL.g0_i_m2_1 ),
            .ltout(\CONTROL.g0_i_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_7_LC_18_24_6 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_7_LC_18_24_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.addrstackptr_7_LC_18_24_6 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \CONTROL.addrstackptr_7_LC_18_24_6  (
            .in0(N__42335),
            .in1(N__42305),
            .in2(N__42296),
            .in3(N__42293),
            .lcout(\CONTROL.addrstackptrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.increment_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_2_i_1_LC_18_24_7 .C_ON=1'b0;
    defparam \CONTROL.g0_2_i_1_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_2_i_1_LC_18_24_7 .LUT_INIT=16'b1001111111111111;
    LogicCell40 \CONTROL.g0_2_i_1_LC_18_24_7  (
            .in0(N__54634),
            .in1(N__42248),
            .in2(N__72319),
            .in3(N__55422),
            .lcout(\CONTROL.g0_2_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m381_am_LC_18_25_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m381_am_LC_18_25_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m381_am_LC_18_25_0 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m381_am_LC_18_25_0  (
            .in0(N__74410),
            .in1(N__76609),
            .in2(N__47885),
            .in3(N__75856),
            .lcout(\PROM.ROMDATA.m381_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m382_ns_1_LC_18_25_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m382_ns_1_LC_18_25_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m382_ns_1_LC_18_25_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m382_ns_1_LC_18_25_5  (
            .in0(N__42131),
            .in1(N__79341),
            .in2(N__47897),
            .in3(N__79846),
            .lcout(\PROM.ROMDATA.m382_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHEO982_2_LC_19_8_0 .C_ON=1'b0;
    defparam \ALU.d_RNIHEO982_2_LC_19_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHEO982_2_LC_19_8_0 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIHEO982_2_LC_19_8_0  (
            .in0(N__60187),
            .in1(N__66240),
            .in2(N__42113),
            .in3(N__66047),
            .lcout(),
            .ltout(\ALU.N_858_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7RHUG5_2_LC_19_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNI7RHUG5_2_LC_19_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7RHUG5_2_LC_19_8_1 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.d_RNI7RHUG5_2_LC_19_8_1  (
            .in0(N__68931),
            .in1(N__42575),
            .in2(N__42095),
            .in3(N__68526),
            .lcout(),
            .ltout(\ALU.rshift_15_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0V48BA_2_LC_19_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNI0V48BA_2_LC_19_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0V48BA_2_LC_19_8_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI0V48BA_2_LC_19_8_2  (
            .in0(N__68527),
            .in1(N__56474),
            .in2(N__42092),
            .in3(N__56491),
            .lcout(\ALU.rshift_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9VEDD1_0_4_LC_19_8_4 .C_ON=1'b0;
    defparam \ALU.d_RNI9VEDD1_0_4_LC_19_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9VEDD1_0_4_LC_19_8_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.d_RNI9VEDD1_0_4_LC_19_8_4  (
            .in0(N__59637),
            .in1(N__66045),
            .in2(N__59911),
            .in3(N__66768),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5MBM92_6_LC_19_8_5 .C_ON=1'b0;
    defparam \ALU.d_RNI5MBM92_6_LC_19_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5MBM92_6_LC_19_8_5 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.d_RNI5MBM92_6_LC_19_8_5  (
            .in0(N__66046),
            .in1(N__62587),
            .in2(N__42089),
            .in3(N__62233),
            .lcout(\ALU.N_862 ),
            .ltout(\ALU.N_862_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFVCT15_6_LC_19_8_6 .C_ON=1'b0;
    defparam \ALU.d_RNIFVCT15_6_LC_19_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFVCT15_6_LC_19_8_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.d_RNIFVCT15_6_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(N__56490),
            .in2(N__42569),
            .in3(N__68930),
            .lcout(),
            .ltout(\ALU.N_922_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1AHUF8_2_LC_19_8_7 .C_ON=1'b0;
    defparam \ALU.d_RNI1AHUF8_2_LC_19_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1AHUF8_2_LC_19_8_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNI1AHUF8_2_LC_19_8_7  (
            .in0(_gnd_net_),
            .in1(N__52684),
            .in2(N__42566),
            .in3(N__42563),
            .lcout(\ALU.d_RNI1AHUF8Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_293_c_RNIOCJMD9_LC_19_9_0 .C_ON=1'b1;
    defparam \ALU.mult_293_c_RNIOCJMD9_LC_19_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_293_c_RNIOCJMD9_LC_19_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ALU.mult_293_c_RNIOCJMD9_LC_19_9_0  (
            .in0(N__42464),
            .in1(N__42710),
            .in2(N__42446),
            .in3(_gnd_net_),
            .lcout(\ALU.mult_293_c_RNIOCJMDZ0Z9 ),
            .ltout(),
            .carryin(bfn_19_9_0_),
            .carryout(\ALU.mult_21_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_464_c_RNIRCBMA3_LC_19_9_1 .C_ON=1'b1;
    defparam \ALU.mult_464_c_RNIRCBMA3_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_464_c_RNIRCBMA3_LC_19_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_464_c_RNIRCBMA3_LC_19_9_1  (
            .in0(_gnd_net_),
            .in1(N__42683),
            .in2(N__42425),
            .in3(N__42404),
            .lcout(\ALU.mult_21_11 ),
            .ltout(),
            .carryin(\ALU.mult_21_c10 ),
            .carryout(\ALU.mult_21_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_467_c_RNISOO9S3_LC_19_9_2 .C_ON=1'b1;
    defparam \ALU.mult_467_c_RNISOO9S3_LC_19_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_467_c_RNISOO9S3_LC_19_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_467_c_RNISOO9S3_LC_19_9_2  (
            .in0(_gnd_net_),
            .in1(N__42665),
            .in2(N__45902),
            .in3(N__42389),
            .lcout(\ALU.mult_21_12 ),
            .ltout(),
            .carryin(\ALU.mult_21_c11 ),
            .carryout(\ALU.mult_21_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_470_c_RNIB61LK3_LC_19_9_3 .C_ON=1'b1;
    defparam \ALU.mult_470_c_RNIB61LK3_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_470_c_RNIB61LK3_LC_19_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_470_c_RNIB61LK3_LC_19_9_3  (
            .in0(_gnd_net_),
            .in1(N__42641),
            .in2(N__45869),
            .in3(N__42380),
            .lcout(\ALU.mult_21_13 ),
            .ltout(),
            .carryin(\ALU.mult_21_c12 ),
            .carryout(\ALU.mult_21_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_473_c_RNIR822C3_LC_19_9_4 .C_ON=1'b1;
    defparam \ALU.mult_473_c_RNIR822C3_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_473_c_RNIR822C3_LC_19_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_473_c_RNIR822C3_LC_19_9_4  (
            .in0(_gnd_net_),
            .in1(N__42602),
            .in2(N__45836),
            .in3(N__42359),
            .lcout(\ALU.mult_21_14 ),
            .ltout(),
            .carryin(\ALU.mult_21_c13 ),
            .carryout(\ALU.mult_21_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_476_c_RNIFLP0O7_LC_19_9_5 .C_ON=1'b0;
    defparam \ALU.mult_476_c_RNIFLP0O7_LC_19_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_476_c_RNIFLP0O7_LC_19_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_476_c_RNIFLP0O7_LC_19_9_5  (
            .in0(N__42854),
            .in1(N__42356),
            .in2(_gnd_net_),
            .in3(N__42350),
            .lcout(\ALU.mult_476_c_RNIFLP0OZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2BV762_8_LC_19_9_6 .C_ON=1'b0;
    defparam \ALU.d_RNI2BV762_8_LC_19_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2BV762_8_LC_19_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNI2BV762_8_LC_19_9_6  (
            .in0(N__42815),
            .in1(N__42776),
            .in2(_gnd_net_),
            .in3(N__66026),
            .lcout(\ALU.N_866 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_293_c_LC_19_10_0 .C_ON=1'b1;
    defparam \ALU.mult_293_c_LC_19_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_293_c_LC_19_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_293_c_LC_19_10_0  (
            .in0(_gnd_net_),
            .in1(N__42881),
            .in2(N__42755),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_10_0_),
            .carryout(\ALU.mult_9_c9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_293_c_RNIKDLV62_LC_19_10_1 .C_ON=1'b1;
    defparam \ALU.mult_293_c_RNIKDLV62_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_293_c_RNIKDLV62_LC_19_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_293_c_RNIKDLV62_LC_19_10_1  (
            .in0(_gnd_net_),
            .in1(N__42740),
            .in2(N__42728),
            .in3(N__42704),
            .lcout(\ALU.mult_9_10 ),
            .ltout(),
            .carryin(\ALU.mult_9_c9 ),
            .carryout(\ALU.mult_9_c10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_299_c_RNIJ4OGS1_LC_19_10_2 .C_ON=1'b1;
    defparam \ALU.mult_299_c_RNIJ4OGS1_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_299_c_RNIJ4OGS1_LC_19_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_299_c_RNIJ4OGS1_LC_19_10_2  (
            .in0(_gnd_net_),
            .in1(N__42701),
            .in2(N__42695),
            .in3(N__42677),
            .lcout(\ALU.mult_9_11 ),
            .ltout(),
            .carryin(\ALU.mult_9_c10 ),
            .carryout(\ALU.mult_9_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_305_c_RNIVQ5JJ1_LC_19_10_3 .C_ON=1'b1;
    defparam \ALU.mult_305_c_RNIVQ5JJ1_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_305_c_RNIVQ5JJ1_LC_19_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_305_c_RNIVQ5JJ1_LC_19_10_3  (
            .in0(_gnd_net_),
            .in1(N__45947),
            .in2(N__42674),
            .in3(N__42659),
            .lcout(\ALU.mult_9_12 ),
            .ltout(),
            .carryin(\ALU.mult_9_c11 ),
            .carryout(\ALU.mult_9_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_311_c_RNIUDNBM1_LC_19_10_4 .C_ON=1'b1;
    defparam \ALU.mult_311_c_RNIUDNBM1_LC_19_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_311_c_RNIUDNBM1_LC_19_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_311_c_RNIUDNBM1_LC_19_10_4  (
            .in0(_gnd_net_),
            .in1(N__42848),
            .in2(N__42656),
            .in3(N__42635),
            .lcout(\ALU.mult_9_13 ),
            .ltout(),
            .carryin(\ALU.mult_9_c12 ),
            .carryout(\ALU.mult_9_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_317_c_RNID87GM1_LC_19_10_5 .C_ON=1'b1;
    defparam \ALU.mult_317_c_RNID87GM1_LC_19_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_317_c_RNID87GM1_LC_19_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_317_c_RNID87GM1_LC_19_10_5  (
            .in0(_gnd_net_),
            .in1(N__42632),
            .in2(N__42617),
            .in3(N__42596),
            .lcout(\ALU.mult_9_14 ),
            .ltout(),
            .carryin(\ALU.mult_9_c13 ),
            .carryout(\ALU.mult_9_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_323_c_RNIAA0B82_LC_19_10_6 .C_ON=1'b0;
    defparam \ALU.mult_323_c_RNIAA0B82_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_323_c_RNIAA0B82_LC_19_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_323_c_RNIAA0B82_LC_19_10_6  (
            .in0(N__42593),
            .in1(N__45821),
            .in2(N__45938),
            .in3(N__42578),
            .lcout(\ALU.mult_323_c_RNIAA0BZ0Z82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGD2441_8_LC_19_11_1 .C_ON=1'b0;
    defparam \ALU.d_RNIGD2441_8_LC_19_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGD2441_8_LC_19_11_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNIGD2441_8_LC_19_11_1  (
            .in0(N__56413),
            .in1(N__62871),
            .in2(N__62021),
            .in3(N__56259),
            .lcout(\ALU.d_RNIGD2441Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIOFVO52_4_LC_19_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNIOFVO52_4_LC_19_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIOFVO52_4_LC_19_11_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.d_RNIOFVO52_4_LC_19_11_2  (
            .in0(N__65968),
            .in1(_gnd_net_),
            .in2(N__45740),
            .in3(N__48059),
            .lcout(\ALU.N_639 ),
            .ltout(\ALU.N_639_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFVCT15_8_LC_19_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIFVCT15_8_LC_19_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFVCT15_8_LC_19_11_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.d_RNIFVCT15_8_LC_19_11_3  (
            .in0(N__68923),
            .in1(_gnd_net_),
            .in2(N__42842),
            .in3(N__46163),
            .lcout(),
            .ltout(\ALU.d_RNIFVCT15Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4U6858_2_LC_19_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNI4U6858_2_LC_19_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4U6858_2_LC_19_11_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.d_RNI4U6858_2_LC_19_11_4  (
            .in0(_gnd_net_),
            .in1(N__42839),
            .in2(N__42824),
            .in3(N__68458),
            .lcout(\ALU.lshift_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIR02AP_10_LC_19_11_5 .C_ON=1'b0;
    defparam \ALU.c_RNIR02AP_10_LC_19_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIR02AP_10_LC_19_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.c_RNIR02AP_10_LC_19_11_5  (
            .in0(N__61703),
            .in1(N__61460),
            .in2(_gnd_net_),
            .in3(N__66704),
            .lcout(\ALU.N_851 ),
            .ltout(\ALU.N_851_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINT9PO2_0_10_LC_19_11_6 .C_ON=1'b0;
    defparam \ALU.c_RNINT9PO2_0_10_LC_19_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINT9PO2_0_10_LC_19_11_6 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \ALU.c_RNINT9PO2_0_10_LC_19_11_6  (
            .in0(N__65967),
            .in1(N__62648),
            .in2(N__42797),
            .in3(N__68922),
            .lcout(\ALU.c_RNINT9PO2_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_335_c_RNO_LC_19_11_7 .C_ON=1'b0;
    defparam \ALU.mult_335_c_RNO_LC_19_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_335_c_RNO_LC_19_11_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.mult_335_c_RNO_LC_19_11_7  (
            .in0(N__61702),
            .in1(N__65966),
            .in2(N__66773),
            .in3(N__61461),
            .lcout(\ALU.mult_335_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIQ12IP_12_LC_19_12_0 .C_ON=1'b0;
    defparam \ALU.c_RNIQ12IP_12_LC_19_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIQ12IP_12_LC_19_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIQ12IP_12_LC_19_12_0  (
            .in0(N__66701),
            .in1(N__60990),
            .in2(_gnd_net_),
            .in3(N__61211),
            .lcout(\ALU.N_978 ),
            .ltout(\ALU.N_978_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIE08272_12_LC_19_12_1 .C_ON=1'b0;
    defparam \ALU.c_RNIE08272_12_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIE08272_12_LC_19_12_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.c_RNIE08272_12_LC_19_12_1  (
            .in0(_gnd_net_),
            .in1(N__62655),
            .in2(N__42779),
            .in3(N__66013),
            .lcout(\ALU.N_967 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIEOKO_1_LC_19_12_2 .C_ON=1'b0;
    defparam \ALU.d_RNIIEOKO_1_LC_19_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIEOKO_1_LC_19_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU.d_RNIIEOKO_1_LC_19_12_2  (
            .in0(N__65557),
            .in1(N__63150),
            .in2(_gnd_net_),
            .in3(N__42899),
            .lcout(\ALU.d_RNIIEOKOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI48CC42_2_LC_19_12_3 .C_ON=1'b0;
    defparam \ALU.d_RNI48CC42_2_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI48CC42_2_LC_19_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNI48CC42_2_LC_19_12_3  (
            .in0(N__45724),
            .in1(N__47978),
            .in2(_gnd_net_),
            .in3(N__66014),
            .lcout(\ALU.N_635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2HF0A9_8_LC_19_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNI2HF0A9_8_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2HF0A9_8_LC_19_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNI2HF0A9_8_LC_19_12_4  (
            .in0(N__46052),
            .in1(N__42887),
            .in2(_gnd_net_),
            .in3(N__68528),
            .lcout(\ALU.rshift_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIO8DPO_14_LC_19_12_5 .C_ON=1'b0;
    defparam \ALU.c_RNIO8DPO_14_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIO8DPO_14_LC_19_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.c_RNIO8DPO_14_LC_19_12_5  (
            .in0(N__63809),
            .in1(N__63645),
            .in2(_gnd_net_),
            .in3(N__66700),
            .lcout(\ALU.N_980 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIG8JO24_15_LC_19_13_0 .C_ON=1'b0;
    defparam \ALU.c_RNIG8JO24_15_LC_19_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIG8JO24_15_LC_19_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIG8JO24_15_LC_19_13_0  (
            .in0(N__68790),
            .in1(N__42868),
            .in2(_gnd_net_),
            .in3(N__43183),
            .lcout(\ALU.N_1026 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_293_c_RNO_0_LC_19_13_1 .C_ON=1'b0;
    defparam \ALU.mult_293_c_RNO_0_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_293_c_RNO_0_LC_19_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_293_c_RNO_0_LC_19_13_1  (
            .in0(_gnd_net_),
            .in1(N__62805),
            .in2(_gnd_net_),
            .in3(N__66718),
            .lcout(\ALU.mult_293_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIN266M_11_LC_19_13_3 .C_ON=1'b0;
    defparam \ALU.c_RNIN266M_11_LC_19_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIN266M_11_LC_19_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.c_RNIN266M_11_LC_19_13_3  (
            .in0(N__61434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68789),
            .lcout(\ALU.c_RNIN266MZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNITTCO62_10_LC_19_13_4 .C_ON=1'b0;
    defparam \ALU.c_RNITTCO62_10_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNITTCO62_10_LC_19_13_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNITTCO62_10_LC_19_13_4  (
            .in0(_gnd_net_),
            .in1(N__66080),
            .in2(N__46117),
            .in3(N__46066),
            .lcout(\ALU.N_867 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNID11991_15_LC_19_13_5 .C_ON=1'b0;
    defparam \ALU.c_RNID11991_15_LC_19_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNID11991_15_LC_19_13_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ALU.c_RNID11991_15_LC_19_13_5  (
            .in0(N__63658),
            .in1(N__66082),
            .in2(_gnd_net_),
            .in3(N__66720),
            .lcout(\ALU.N_1011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIET09P_12_LC_19_13_6 .C_ON=1'b0;
    defparam \ALU.c_RNIET09P_12_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIET09P_12_LC_19_13_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNIET09P_12_LC_19_13_6  (
            .in0(N__66719),
            .in1(N__61435),
            .in2(_gnd_net_),
            .in3(N__61212),
            .lcout(\ALU.N_852 ),
            .ltout(\ALU.N_852_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIR8GG72_12_LC_19_13_7 .C_ON=1'b0;
    defparam \ALU.c_RNIR8GG72_12_LC_19_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIR8GG72_12_LC_19_13_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ALU.c_RNIR8GG72_12_LC_19_13_7  (
            .in0(N__53332),
            .in1(_gnd_net_),
            .in2(N__43187),
            .in3(N__66081),
            .lcout(\ALU.N_966 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQQRSN_2_LC_19_14_0 .C_ON=1'b0;
    defparam \ALU.d_RNIQQRSN_2_LC_19_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQQRSN_2_LC_19_14_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ALU.d_RNIQQRSN_2_LC_19_14_0  (
            .in0(N__65565),
            .in1(_gnd_net_),
            .in2(N__66767),
            .in3(N__66287),
            .lcout(\ALU.N_766 ),
            .ltout(\ALU.N_766_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0KELT1_2_LC_19_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNI0KELT1_2_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0KELT1_2_LC_19_14_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNI0KELT1_2_LC_19_14_1  (
            .in0(N__66079),
            .in1(_gnd_net_),
            .in2(N__43169),
            .in3(N__48583),
            .lcout(\ALU.N_634 ),
            .ltout(\ALU.N_634_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILTB1L4_2_LC_19_14_2 .C_ON=1'b0;
    defparam \ALU.d_RNILTB1L4_2_LC_19_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILTB1L4_2_LC_19_14_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.d_RNILTB1L4_2_LC_19_14_2  (
            .in0(_gnd_net_),
            .in1(N__43590),
            .in2(N__43127),
            .in3(N__68921),
            .lcout(),
            .ltout(\ALU.N_811_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIK8M6K5_6_LC_19_14_3 .C_ON=1'b0;
    defparam \ALU.d_RNIK8M6K5_6_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIK8M6K5_6_LC_19_14_3 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \ALU.d_RNIK8M6K5_6_LC_19_14_3  (
            .in0(N__70197),
            .in1(N__51262),
            .in2(N__43124),
            .in3(N__68529),
            .lcout(\ALU.d_RNIK8M6K5Z0Z_6 ),
            .ltout(\ALU.d_RNIK8M6K5Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_6_LC_19_14_4 .C_ON=1'b0;
    defparam \ALU.a_6_LC_19_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.a_6_LC_19_14_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.a_6_LC_19_14_4  (
            .in0(N__43055),
            .in1(_gnd_net_),
            .in2(N__42995),
            .in3(N__42990),
            .lcout(\ALU.aZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73161),
            .ce(N__71199),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKRBVN_0_4_LC_19_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNIKRBVN_0_4_LC_19_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKRBVN_0_4_LC_19_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIKRBVN_0_4_LC_19_14_5  (
            .in0(N__60237),
            .in1(N__59849),
            .in2(_gnd_net_),
            .in3(N__66746),
            .lcout(\ALU.N_606 ),
            .ltout(\ALU.N_606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAC0J42_2_LC_19_14_6 .C_ON=1'b0;
    defparam \ALU.d_RNIAC0J42_2_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAC0J42_2_LC_19_14_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.d_RNIAC0J42_2_LC_19_14_6  (
            .in0(_gnd_net_),
            .in1(N__42908),
            .in2(N__42902),
            .in3(N__66077),
            .lcout(\ALU.N_636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDBRC52_4_LC_19_14_7 .C_ON=1'b0;
    defparam \ALU.d_RNIDBRC52_4_LC_19_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDBRC52_4_LC_19_14_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNIDBRC52_4_LC_19_14_7  (
            .in0(N__66078),
            .in1(N__48672),
            .in2(_gnd_net_),
            .in3(N__43610),
            .lcout(\ALU.N_638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m0_am_2_LC_19_15_0 .C_ON=1'b0;
    defparam \ALU.a_15_m0_am_2_LC_19_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m0_am_2_LC_19_15_0 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \ALU.a_15_m0_am_2_LC_19_15_0  (
            .in0(N__43531),
            .in1(N__49830),
            .in2(_gnd_net_),
            .in3(N__43507),
            .lcout(\ALU.a_15_m0_amZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGE45L7_9_LC_19_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIGE45L7_9_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGE45L7_9_LC_19_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIGE45L7_9_LC_19_15_1  (
            .in0(N__51437),
            .in1(N__48002),
            .in2(_gnd_net_),
            .in3(N__70117),
            .lcout(\ALU.a_15_m1_9 ),
            .ltout(\ALU.a_15_m1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_9_LC_19_15_2 .C_ON=1'b0;
    defparam \ALU.a_9_LC_19_15_2 .SEQ_MODE=4'b1000;
    defparam \ALU.a_9_LC_19_15_2 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \ALU.a_9_LC_19_15_2  (
            .in0(N__66844),
            .in1(N__58552),
            .in2(N__43556),
            .in3(N__52805),
            .lcout(\ALU.aZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73172),
            .ce(N__71198),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIV0F38_0_LC_19_15_3 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIV0F38_0_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIV0F38_0_LC_19_15_3 .LUT_INIT=16'b0111001001110010;
    LogicCell40 \CONTROL.busState_1_RNIV0F38_0_LC_19_15_3  (
            .in0(N__49831),
            .in1(N__43532),
            .in2(N__43511),
            .in3(_gnd_net_),
            .lcout(bus_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI5FSP_4_LC_19_15_4 .C_ON=1'b0;
    defparam \ALU.b_RNI5FSP_4_LC_19_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI5FSP_4_LC_19_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_RNI5FSP_4_LC_19_15_4  (
            .in0(N__46897),
            .in1(N__44139),
            .in2(_gnd_net_),
            .in3(N__43444),
            .lcout(\ALU.b_RNI5FSPZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIHV2S_9_LC_19_15_5 .C_ON=1'b0;
    defparam \ALU.c_RNIHV2S_9_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIHV2S_9_LC_19_15_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIHV2S_9_LC_19_15_5  (
            .in0(N__72348),
            .in1(N__46654),
            .in2(_gnd_net_),
            .in3(N__46898),
            .lcout(\ALU.c_RNIHV2SZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9R8E_4_LC_19_15_6 .C_ON=1'b0;
    defparam \ALU.d_RNI9R8E_4_LC_19_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9R8E_4_LC_19_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNI9R8E_4_LC_19_15_6  (
            .in0(N__46896),
            .in1(N__43402),
            .in2(_gnd_net_),
            .in3(N__43349),
            .lcout(\ALU.d_RNI9R8EZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI83KC1_14_LC_19_15_7 .C_ON=1'b0;
    defparam \ALU.b_RNI83KC1_14_LC_19_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI83KC1_14_LC_19_15_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.b_RNI83KC1_14_LC_19_15_7  (
            .in0(N__57582),
            .in1(N__67964),
            .in2(_gnd_net_),
            .in3(N__43303),
            .lcout(\ALU.b_RNI83KC1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_7_LC_19_16_0 .C_ON=1'b0;
    defparam \ALU.h_7_LC_19_16_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_7_LC_19_16_0 .LUT_INIT=16'b0101110101011000;
    LogicCell40 \ALU.h_7_LC_19_16_0  (
            .in0(N__58886),
            .in1(N__51931),
            .in2(N__67242),
            .in3(N__51853),
            .lcout(h_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73183),
            .ce(N__69449),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIO7K62_7_LC_19_16_1 .C_ON=1'b0;
    defparam \ALU.c_RNIO7K62_7_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIO7K62_7_LC_19_16_1 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \ALU.c_RNIO7K62_7_LC_19_16_1  (
            .in0(N__46402),
            .in1(N__43937),
            .in2(N__48867),
            .in3(N__46780),
            .lcout(\ALU.N_1204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISJ0R1_7_LC_19_16_2 .C_ON=1'b0;
    defparam \ALU.d_RNISJ0R1_7_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISJ0R1_7_LC_19_16_2 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \ALU.d_RNISJ0R1_7_LC_19_16_2  (
            .in0(N__46781),
            .in1(N__51806),
            .in2(N__43822),
            .in3(N__43616),
            .lcout(),
            .ltout(\ALU.N_1252_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO5IF4_7_LC_19_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNIO5IF4_7_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO5IF4_7_LC_19_16_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIO5IF4_7_LC_19_16_3  (
            .in0(_gnd_net_),
            .in1(N__53889),
            .in2(N__43649),
            .in3(N__43646),
            .lcout(),
            .ltout(\ALU.d_RNIO5IF4Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIM3JB6_7_LC_19_16_4 .C_ON=1'b0;
    defparam \ALU.d_RNIM3JB6_7_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIM3JB6_7_LC_19_16_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIM3JB6_7_LC_19_16_4  (
            .in0(_gnd_net_),
            .in1(N__71436),
            .in2(N__43640),
            .in3(N__43637),
            .lcout(),
            .ltout(\ALU.d_RNIM3JB6Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3GMNC_7_LC_19_16_5 .C_ON=1'b0;
    defparam \ALU.d_RNI3GMNC_7_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3GMNC_7_LC_19_16_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ALU.d_RNI3GMNC_7_LC_19_16_5  (
            .in0(N__53305),
            .in1(N__49580),
            .in2(N__43622),
            .in3(N__43759),
            .lcout(\ALU.status_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIB0OT_7_LC_19_17_0 .C_ON=1'b0;
    defparam \ALU.e_RNIB0OT_7_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIB0OT_7_LC_19_17_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.e_RNIB0OT_7_LC_19_17_0  (
            .in0(N__46610),
            .in1(N__43915),
            .in2(N__46298),
            .in3(N__47273),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIN3QQ1_7_LC_19_17_1 .C_ON=1'b0;
    defparam \ALU.c_RNIN3QQ1_7_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIN3QQ1_7_LC_19_17_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.c_RNIN3QQ1_7_LC_19_17_1  (
            .in0(N__46403),
            .in1(N__48871),
            .in2(N__43619),
            .in3(N__47190),
            .lcout(\ALU.N_1092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNID4971_7_LC_19_17_2 .C_ON=1'b0;
    defparam \ALU.b_RNID4971_7_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNID4971_7_LC_19_17_2 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.b_RNID4971_7_LC_19_17_2  (
            .in0(N__53401),
            .in1(N__48346),
            .in2(N__49081),
            .in3(N__43979),
            .lcout(\ALU.operand2_6_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIBU251_7_LC_19_17_3 .C_ON=1'b0;
    defparam \ALU.e_RNIBU251_7_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIBU251_7_LC_19_17_3 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.e_RNIBU251_7_LC_19_17_3  (
            .in0(N__43980),
            .in1(N__46294),
            .in2(N__46609),
            .in3(N__53400),
            .lcout(\ALU.operand2_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNID6UV_7_LC_19_17_4 .C_ON=1'b0;
    defparam \ALU.b_RNID6UV_7_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNID6UV_7_LC_19_17_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.b_RNID6UV_7_LC_19_17_4  (
            .in0(N__48347),
            .in1(N__43914),
            .in2(N__49080),
            .in3(N__47272),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRF6F1_7_LC_19_17_5 .C_ON=1'b0;
    defparam \ALU.d_RNIRF6F1_7_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRF6F1_7_LC_19_17_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIRF6F1_7_LC_19_17_5  (
            .in0(N__43815),
            .in1(N__51805),
            .in2(N__43799),
            .in3(N__47191),
            .lcout(),
            .ltout(\ALU.N_1140_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILNEJ3_7_LC_19_17_6 .C_ON=1'b0;
    defparam \ALU.d_RNILNEJ3_7_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILNEJ3_7_LC_19_17_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNILNEJ3_7_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(N__54118),
            .in2(N__43796),
            .in3(N__43793),
            .lcout(aluOut_7),
            .ltout(aluOut_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIG8VE5_1_LC_19_17_7 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIG8VE5_1_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIG8VE5_1_LC_19_17_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \CONTROL.busState_1_RNIG8VE5_1_LC_19_17_7  (
            .in0(N__50305),
            .in1(N__43787),
            .in2(N__43772),
            .in3(N__50213),
            .lcout(N_200),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m267_LC_19_18_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m267_LC_19_18_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m267_LC_19_18_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m267_LC_19_18_0  (
            .in0(N__78769),
            .in1(N__78026),
            .in2(N__75993),
            .in3(N__77295),
            .lcout(),
            .ltout(\PROM.ROMDATA.m267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m442_LC_19_18_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m442_LC_19_18_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m442_LC_19_18_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m442_LC_19_18_1  (
            .in0(N__44307),
            .in1(N__79788),
            .in2(N__43748),
            .in3(N__76585),
            .lcout(\PROM.ROMDATA.m442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m282_LC_19_18_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m282_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m282_LC_19_18_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m282_LC_19_18_2  (
            .in0(N__78766),
            .in1(N__78023),
            .in2(N__75990),
            .in3(N__77292),
            .lcout(\PROM.ROMDATA.m282 ),
            .ltout(\PROM.ROMDATA.m282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.dout_13_LC_19_18_3 .C_ON=1'b0;
    defparam \CONTROL.dout_13_LC_19_18_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.dout_13_LC_19_18_3 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \CONTROL.dout_13_LC_19_18_3  (
            .in0(N__44308),
            .in1(N__43703),
            .in2(N__43679),
            .in3(N__76586),
            .lcout(\CONTROL.ctrlOut_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.dout_13C_net ),
            .ce(N__44397),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m444_bm_LC_19_18_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m444_bm_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m444_bm_LC_19_18_4 .LUT_INIT=16'b0001000000000111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m444_bm_LC_19_18_4  (
            .in0(N__78767),
            .in1(N__78024),
            .in2(N__75991),
            .in3(N__77293),
            .lcout(),
            .ltout(\PROM.ROMDATA.m444_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m447_ns_1_LC_19_18_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m447_ns_1_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m447_ns_1_LC_19_18_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m447_ns_1_LC_19_18_5  (
            .in0(N__44336),
            .in1(N__79787),
            .in2(N__44327),
            .in3(N__76584),
            .lcout(\PROM.ROMDATA.m447_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m289_LC_19_18_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m289_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m289_LC_19_18_6 .LUT_INIT=16'b0000000100001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m289_LC_19_18_6  (
            .in0(N__78768),
            .in1(N__78025),
            .in2(N__75992),
            .in3(N__77294),
            .lcout(\PROM.ROMDATA.m289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m418_ns_LC_19_19_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m418_ns_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m418_ns_LC_19_19_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m418_ns_LC_19_19_1  (
            .in0(N__64169),
            .in1(N__72684),
            .in2(N__44294),
            .in3(N__79300),
            .lcout(PROM_ROMDATA_dintern_19ro),
            .ltout(PROM_ROMDATA_dintern_19ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_19dflt_LC_19_19_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_19dflt_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_19dflt_LC_19_19_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_19dflt_LC_19_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44258),
            .in3(N__72256),
            .lcout(controlWord_19),
            .ltout(controlWord_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_3_LC_19_19_3 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_3_LC_19_19_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_3_LC_19_19_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \CONTROL.ramAddReg_3_LC_19_19_3  (
            .in0(N__70549),
            .in1(N__44243),
            .in2(N__44195),
            .in3(N__70790),
            .lcout(A3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_3C_net ),
            .ce(N__70330),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_4_LC_19_19_4 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_4_LC_19_19_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_4_LC_19_19_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.ramAddReg_4_LC_19_19_4  (
            .in0(N__44192),
            .in1(N__70789),
            .in2(N__44162),
            .in3(N__70551),
            .lcout(A4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_3C_net ),
            .ce(N__70330),
            .sr(_gnd_net_));
    defparam \RAM.un1_WR_105_0_7_LC_19_19_5 .C_ON=1'b0;
    defparam \RAM.un1_WR_105_0_7_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \RAM.un1_WR_105_0_7_LC_19_19_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RAM.un1_WR_105_0_7_LC_19_19_5  (
            .in0(N__44101),
            .in1(N__44059),
            .in2(N__44962),
            .in3(N__44032),
            .lcout(\RAM.un1_WR_105_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_15_LC_19_19_6 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_15_LC_19_19_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_15_LC_19_19_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.ramAddReg_15_LC_19_19_6  (
            .in0(N__45020),
            .in1(N__70788),
            .in2(N__53534),
            .in3(N__70550),
            .lcout(A15_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_3C_net ),
            .ce(N__70330),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m266_LC_19_20_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m266_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m266_LC_19_20_0 .LUT_INIT=16'b0111111011111111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m266_LC_19_20_0  (
            .in0(N__78731),
            .in1(N__77199),
            .in2(N__75614),
            .in3(N__77909),
            .lcout(\PROM.ROMDATA.m266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m446_bm_LC_19_20_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m446_bm_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m446_bm_LC_19_20_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m446_bm_LC_19_20_1  (
            .in0(N__64007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__75304),
            .lcout(\PROM.ROMDATA.m446_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m157_LC_19_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m157_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m157_LC_19_20_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m157_LC_19_20_2  (
            .in0(N__78732),
            .in1(N__77200),
            .in2(_gnd_net_),
            .in3(N__77910),
            .lcout(\PROM.ROMDATA.m157 ),
            .ltout(\PROM.ROMDATA.m157_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m268_LC_19_20_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m268_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m268_LC_19_20_3 .LUT_INIT=16'b1101000100010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m268_LC_19_20_3  (
            .in0(N__44945),
            .in1(N__76603),
            .in2(N__44939),
            .in3(N__75299),
            .lcout(\PROM.ROMDATA.m268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m265_LC_19_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m265_LC_19_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m265_LC_19_20_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m265_LC_19_20_4  (
            .in0(N__78733),
            .in1(N__77201),
            .in2(N__75615),
            .in3(N__77911),
            .lcout(),
            .ltout(\PROM.ROMDATA.m265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m270_bm_LC_19_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m270_bm_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m270_bm_LC_19_20_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m270_bm_LC_19_20_5  (
            .in0(N__79714),
            .in1(_gnd_net_),
            .in2(N__44936),
            .in3(N__44933),
            .lcout(\PROM.ROMDATA.m270_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_6_LC_19_20_6 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_6_LC_19_20_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_6_LC_19_20_6 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \CONTROL.aluOperation_6_LC_19_20_6  (
            .in0(N__44909),
            .in1(N__44900),
            .in2(N__44774),
            .in3(N__44704),
            .lcout(aluOperation_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.aluOperation_6C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m278_LC_19_20_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m278_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m278_LC_19_20_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m278_LC_19_20_7  (
            .in0(N__64235),
            .in1(N__76604),
            .in2(N__79830),
            .in3(N__75303),
            .lcout(\PROM.ROMDATA.N_544_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_RNIUD971_LC_19_21_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_RNIUD971_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_18_RNIUD971_LC_19_21_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.programCounter_ret_18_RNIUD971_LC_19_21_0  (
            .in0(N__45144),
            .in1(N__45641),
            .in2(_gnd_net_),
            .in3(N__45296),
            .lcout(progRomAddress_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m258_bm_LC_19_21_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m258_bm_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m258_bm_LC_19_21_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m258_bm_LC_19_21_1  (
            .in0(N__75306),
            .in1(N__64105),
            .in2(N__76579),
            .in3(N__47708),
            .lcout(\PROM.ROMDATA.m258_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_1_LC_19_21_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_1_LC_19_21_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_1_LC_19_21_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_1_LC_19_21_2  (
            .in0(N__45187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73224),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_RNIQ9971_LC_19_21_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_RNIQ9971_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_18_RNIQ9971_LC_19_21_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CONTROL.programCounter_ret_18_RNIQ9971_LC_19_21_3  (
            .in0(N__45161),
            .in1(N__45155),
            .in2(_gnd_net_),
            .in3(N__45143),
            .lcout(progRomAddress_5),
            .ltout(progRomAddress_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m243_1_LC_19_21_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m243_1_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m243_1_LC_19_21_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m243_1_LC_19_21_4  (
            .in0(N__79248),
            .in1(N__76463),
            .in2(N__45098),
            .in3(N__75305),
            .lcout(\PROM.ROMDATA.m243_1 ),
            .ltout(\PROM.ROMDATA.m243_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_1_1_LC_19_21_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_1_1_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m244_ns_1_1_LC_19_21_5 .LUT_INIT=16'b0001101110111011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m244_ns_1_1_LC_19_21_5  (
            .in0(N__72648),
            .in1(N__79751),
            .in2(N__45095),
            .in3(N__64106),
            .lcout(\PROM.ROMDATA.m244_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_0_LC_19_21_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_0_LC_19_21_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_0_LC_19_21_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_19_0_LC_19_21_6  (
            .in0(N__45080),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.dout_reto_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73224),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m260_1_LC_19_21_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m260_1_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m260_1_LC_19_21_7 .LUT_INIT=16'b0101001111110011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m260_1_LC_19_21_7  (
            .in0(N__45065),
            .in1(N__79249),
            .in2(N__72725),
            .in3(N__64107),
            .lcout(\PROM.ROMDATA.m260_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNILC5J_2_LC_19_22_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNILC5J_2_LC_19_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNILC5J_2_LC_19_22_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.programCounter_ret_1_RNILC5J_2_LC_19_22_0  (
            .in0(N__55077),
            .in1(N__54803),
            .in2(_gnd_net_),
            .in3(N__47564),
            .lcout(N_417),
            .ltout(N_417_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m27_LC_19_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m27_LC_19_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m27_LC_19_22_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m27_LC_19_22_1  (
            .in0(N__64597),
            .in1(N__64694),
            .in2(N__45326),
            .in3(N__77175),
            .lcout(\PROM.ROMDATA.N_28_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_2_LC_19_22_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_2_LC_19_22_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_2_LC_19_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_2_LC_19_22_2  (
            .in0(N__45323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73236),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNI6OHF_6_LC_19_22_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNI6OHF_6_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNI6OHF_6_LC_19_22_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \CONTROL.programCounter_ret_1_RNI6OHF_6_LC_19_22_3  (
            .in0(N__64596),
            .in1(_gnd_net_),
            .in2(N__47816),
            .in3(N__45614),
            .lcout(\CONTROL.programCounter_ret_1_RNI6OHFZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_3_LC_19_22_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_3_LC_19_22_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_3_LC_19_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_3_LC_19_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45290),
            .lcout(\CONTROL.dout_reto_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73236),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_4_LC_19_22_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_4_LC_19_22_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_4_LC_19_22_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_4_LC_19_22_5  (
            .in0(N__45266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73236),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_N_2L1_LC_19_22_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_N_2L1_LC_19_22_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_N_2L1_LC_19_22_6 .LUT_INIT=16'b0111011101011111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m215_ns_1_N_2L1_LC_19_22_6  (
            .in0(N__75307),
            .in1(N__78943),
            .in2(N__64871),
            .in3(N__78634),
            .lcout(),
            .ltout(\PROM.ROMDATA.m215_ns_1_N_2L1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_LC_19_22_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_LC_19_22_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_LC_19_22_7 .LUT_INIT=16'b0100010001110010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m215_ns_1_LC_19_22_7  (
            .in0(N__79207),
            .in1(N__47714),
            .in2(N__45242),
            .in3(N__76500),
            .lcout(\PROM.ROMDATA.m215_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_3_i_a7_1_LC_19_23_0 .C_ON=1'b0;
    defparam \CONTROL.g0_3_i_a7_1_LC_19_23_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_3_i_a7_1_LC_19_23_0 .LUT_INIT=16'b0111000001110111;
    LogicCell40 \CONTROL.g0_3_i_a7_1_LC_19_23_0  (
            .in0(N__53718),
            .in1(N__53666),
            .in2(N__45523),
            .in3(N__45402),
            .lcout(\CONTROL.g0_3_i_a7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_2_LC_19_23_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_2_LC_19_23_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_2_LC_19_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_2_LC_19_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45206),
            .lcout(CONTROL_addrstack_reto_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73246),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m36_LC_19_23_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m36_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m36_LC_19_23_2 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m36_LC_19_23_2  (
            .in0(N__47570),
            .in1(N__54935),
            .in2(_gnd_net_),
            .in3(N__79286),
            .lcout(\PROM.ROMDATA.m36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m235_LC_19_23_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m235_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m235_LC_19_23_3 .LUT_INIT=16'b0000111001011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m235_LC_19_23_3  (
            .in0(N__77185),
            .in1(N__78806),
            .in2(N__75914),
            .in3(N__77878),
            .lcout(),
            .ltout(\PROM.ROMDATA.N_526_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m238_bm_LC_19_23_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m238_bm_LC_19_23_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m238_bm_LC_19_23_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m238_bm_LC_19_23_4  (
            .in0(N__76534),
            .in1(N__64108),
            .in2(N__45542),
            .in3(N__75736),
            .lcout(\PROM.ROMDATA.m238_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m30_LC_19_23_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m30_LC_19_23_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m30_LC_19_23_5 .LUT_INIT=16'b0100111011111100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m30_LC_19_23_5  (
            .in0(N__77186),
            .in1(N__78807),
            .in2(N__75915),
            .in3(N__77879),
            .lcout(\PROM.ROMDATA.m30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g0_5_0_LC_19_23_6 .C_ON=1'b0;
    defparam \CONTROL.g0_5_0_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g0_5_0_LC_19_23_6 .LUT_INIT=16'b0111000001110111;
    LogicCell40 \CONTROL.g0_5_0_LC_19_23_6  (
            .in0(N__53719),
            .in1(N__53667),
            .in2(N__45524),
            .in3(N__45403),
            .lcout(\CONTROL.g0_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m258_am_LC_19_23_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m258_am_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m258_am_LC_19_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m258_am_LC_19_23_7  (
            .in0(N__47687),
            .in1(N__47693),
            .in2(_gnd_net_),
            .in3(N__76535),
            .lcout(\PROM.ROMDATA.m258_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNINE5J_3_LC_19_24_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNINE5J_3_LC_19_24_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNINE5J_3_LC_19_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.programCounter_ret_1_RNINE5J_3_LC_19_24_0  (
            .in0(N__55078),
            .in1(N__51125),
            .in2(_gnd_net_),
            .in3(N__47639),
            .lcout(N_418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m69_LC_19_24_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m69_LC_19_24_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m69_LC_19_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m69_LC_19_24_1  (
            .in0(_gnd_net_),
            .in1(N__64340),
            .in2(_gnd_net_),
            .in3(N__74023),
            .lcout(PROM_ROMDATA_dintern_31_0__N_555_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m53_am_LC_19_24_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m53_am_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m53_am_LC_19_24_2 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m53_am_LC_19_24_2  (
            .in0(N__45566),
            .in1(N__51368),
            .in2(_gnd_net_),
            .in3(N__76605),
            .lcout(\PROM.ROMDATA.m53_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_5_LC_19_24_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_5_LC_19_24_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_5_LC_19_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_5_LC_19_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45680),
            .lcout(\CONTROL.dout_reto_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73256),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_RNIV5IG_6_LC_19_24_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_RNIV5IG_6_LC_19_24_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_19_RNIV5IG_6_LC_19_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_19_RNIV5IG_6_LC_19_24_4  (
            .in0(N__45572),
            .in1(N__45613),
            .in2(_gnd_net_),
            .in3(N__64598),
            .lcout(\CONTROL.programCounter_ret_19_RNIV5IGZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_6_LC_19_24_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_6_LC_19_24_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_6_LC_19_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_6_LC_19_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45632),
            .lcout(\CONTROL.addrstack_reto_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73256),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m53_bm_LC_19_24_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m53_bm_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m53_bm_LC_19_24_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m53_bm_LC_19_24_6  (
            .in0(N__47804),
            .in1(N__45599),
            .in2(_gnd_net_),
            .in3(N__76606),
            .lcout(\PROM.ROMDATA.m53_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_6_LC_19_24_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_6_LC_19_24_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_6_LC_19_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_6_LC_19_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45593),
            .lcout(\CONTROL.dout_reto_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73256),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m7_LC_19_25_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m7_LC_19_25_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m7_LC_19_25_0 .LUT_INIT=16'b0101010001100001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m7_LC_19_25_0  (
            .in0(N__77875),
            .in1(N__78831),
            .in2(N__75916),
            .in3(N__77187),
            .lcout(\PROM.ROMDATA.m7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m392_bm_LC_19_25_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m392_bm_LC_19_25_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m392_bm_LC_19_25_1 .LUT_INIT=16'b0001000000001001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m392_bm_LC_19_25_1  (
            .in0(N__77188),
            .in1(N__78808),
            .in2(N__76002),
            .in3(N__77876),
            .lcout(),
            .ltout(\PROM.ROMDATA.m392_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m392_ns_LC_19_25_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m392_ns_LC_19_25_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m392_ns_LC_19_25_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m392_ns_LC_19_25_2  (
            .in0(_gnd_net_),
            .in1(N__47552),
            .in2(N__45560),
            .in3(N__76607),
            .lcout(),
            .ltout(\PROM.ROMDATA.m392_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m401_ns_1_LC_19_25_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m401_ns_1_LC_19_25_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m401_ns_1_LC_19_25_3 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m401_ns_1_LC_19_25_3  (
            .in0(N__79418),
            .in1(N__47855),
            .in2(N__45557),
            .in3(N__79808),
            .lcout(\PROM.ROMDATA.m401_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m396_bm_LC_19_25_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m396_bm_LC_19_25_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m396_bm_LC_19_25_4 .LUT_INIT=16'b0001010001000010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m396_bm_LC_19_25_4  (
            .in0(N__77877),
            .in1(N__78832),
            .in2(N__75917),
            .in3(N__77189),
            .lcout(\PROM.ROMDATA.m396_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m396_am_LC_19_25_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m396_am_LC_19_25_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m396_am_LC_19_25_5 .LUT_INIT=16'b1100110000100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m396_am_LC_19_25_5  (
            .in0(N__78995),
            .in1(N__45809),
            .in2(_gnd_net_),
            .in3(N__75746),
            .lcout(),
            .ltout(\PROM.ROMDATA.m396_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m396_ns_LC_19_25_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m396_ns_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m396_ns_LC_19_25_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m396_ns_LC_19_25_6  (
            .in0(_gnd_net_),
            .in1(N__45785),
            .in2(N__45779),
            .in3(N__76608),
            .lcout(),
            .ltout(\PROM.ROMDATA.m396_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m401_ns_LC_19_25_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m401_ns_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m401_ns_LC_19_25_7 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m401_ns_LC_19_25_7  (
            .in0(N__79419),
            .in1(N__47771),
            .in2(N__45776),
            .in3(N__45773),
            .lcout(\PROM.ROMDATA.m401_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBQSTO_11_LC_20_9_0 .C_ON=1'b0;
    defparam \ALU.c_RNIBQSTO_11_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBQSTO_11_LC_20_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.c_RNIBQSTO_11_LC_20_9_0  (
            .in0(_gnd_net_),
            .in1(N__61470),
            .in2(_gnd_net_),
            .in3(N__66049),
            .lcout(\ALU.c_RNIBQSTOZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID9MMO_4_LC_20_9_1 .C_ON=1'b0;
    defparam \ALU.d_RNID9MMO_4_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID9MMO_4_LC_20_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNID9MMO_4_LC_20_9_1  (
            .in0(N__59910),
            .in1(N__59638),
            .in2(_gnd_net_),
            .in3(N__66763),
            .lcout(\ALU.N_607 ),
            .ltout(\ALU.N_607_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4DGL42_4_LC_20_9_2 .C_ON=1'b0;
    defparam \ALU.d_RNI4DGL42_4_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4DGL42_4_LC_20_9_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.d_RNI4DGL42_4_LC_20_9_2  (
            .in0(_gnd_net_),
            .in1(N__45728),
            .in2(N__45683),
            .in3(N__66050),
            .lcout(\ALU.N_637 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIG5G6F1_10_LC_20_9_3 .C_ON=1'b0;
    defparam \ALU.c_RNIG5G6F1_10_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIG5G6F1_10_LC_20_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.c_RNIG5G6F1_10_LC_20_9_3  (
            .in0(N__61471),
            .in1(N__61636),
            .in2(N__66083),
            .in3(N__68909),
            .lcout(\ALU.c_RNIG5G6F1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIT73F71_10_LC_20_9_4 .C_ON=1'b0;
    defparam \ALU.c_RNIT73F71_10_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIT73F71_10_LC_20_9_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.c_RNIT73F71_10_LC_20_9_4  (
            .in0(N__68910),
            .in1(N__61472),
            .in2(N__61675),
            .in3(N__68507),
            .lcout(\ALU.c_RNIT73F71Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFHB5A2_8_LC_20_9_5 .C_ON=1'b0;
    defparam \ALU.d_RNIFHB5A2_8_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFHB5A2_8_LC_20_9_5 .LUT_INIT=16'b1011100100110001;
    LogicCell40 \ALU.d_RNIFHB5A2_8_LC_20_9_5  (
            .in0(N__66051),
            .in1(N__45962),
            .in2(N__62026),
            .in3(N__62883),
            .lcout(\ALU.N_643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4N3K21_8_LC_20_9_6 .C_ON=1'b0;
    defparam \ALU.d_RNI4N3K21_8_LC_20_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4N3K21_8_LC_20_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI4N3K21_8_LC_20_9_6  (
            .in0(N__62884),
            .in1(N__56416),
            .in2(N__68530),
            .in3(N__62010),
            .lcout(\ALU.d_RNI4N3K21Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIH8D821_8_LC_20_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNIH8D821_8_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIH8D821_8_LC_20_9_7 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.d_RNIH8D821_8_LC_20_9_7  (
            .in0(N__55949),
            .in1(N__62882),
            .in2(N__62025),
            .in3(N__56120),
            .lcout(\ALU.d_RNIH8D821Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_335_c_LC_20_10_0 .C_ON=1'b1;
    defparam \ALU.mult_335_c_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_335_c_LC_20_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_335_c_LC_20_10_0  (
            .in0(_gnd_net_),
            .in1(N__46127),
            .in2(N__45929),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_10_0_),
            .carryout(\ALU.mult_11_c11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_335_c_RNI96NH82_LC_20_10_1 .C_ON=1'b1;
    defparam \ALU.mult_335_c_RNI96NH82_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_335_c_RNI96NH82_LC_20_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_335_c_RNI96NH82_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__45917),
            .in2(N__45911),
            .in3(N__45893),
            .lcout(\ALU.mult_11_12 ),
            .ltout(),
            .carryin(\ALU.mult_11_c11 ),
            .carryout(\ALU.mult_11_c12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_341_c_RNIVBI3U1_LC_20_10_2 .C_ON=1'b1;
    defparam \ALU.mult_341_c_RNIVBI3U1_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_341_c_RNIVBI3U1_LC_20_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_341_c_RNIVBI3U1_LC_20_10_2  (
            .in0(_gnd_net_),
            .in1(N__45890),
            .in2(N__45878),
            .in3(N__45860),
            .lcout(\ALU.mult_11_13 ),
            .ltout(),
            .carryin(\ALU.mult_11_c12 ),
            .carryout(\ALU.mult_11_c13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_347_c_RNITD0CL1_LC_20_10_3 .C_ON=1'b1;
    defparam \ALU.mult_347_c_RNITD0CL1_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_347_c_RNITD0CL1_LC_20_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_347_c_RNITD0CL1_LC_20_10_3  (
            .in0(_gnd_net_),
            .in1(N__45815),
            .in2(N__45857),
            .in3(N__45827),
            .lcout(\ALU.mult_11_14 ),
            .ltout(),
            .carryin(\ALU.mult_11_c13 ),
            .carryout(\ALU.mult_11_c14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_11_c14_THRU_LUT4_0_LC_20_10_4 .C_ON=1'b0;
    defparam \ALU.mult_11_c14_THRU_LUT4_0_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_11_c14_THRU_LUT4_0_LC_20_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.mult_11_c14_THRU_LUT4_0_LC_20_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45824),
            .lcout(\ALU.mult_11_c14_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIOSF6H_11_LC_20_10_7 .C_ON=1'b0;
    defparam \ALU.c_RNIOSF6H_11_LC_20_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIOSF6H_11_LC_20_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.c_RNIOSF6H_11_LC_20_10_7  (
            .in0(N__61473),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__68395),
            .lcout(\ALU.c_RNIOSF6HZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_335_c_RNO_0_LC_20_11_0 .C_ON=1'b0;
    defparam \ALU.mult_335_c_RNO_0_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_335_c_RNO_0_LC_20_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_335_c_RNO_0_LC_20_11_0  (
            .in0(_gnd_net_),
            .in1(N__61446),
            .in2(_gnd_net_),
            .in3(N__66702),
            .lcout(\ALU.mult_335_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPTT4O_8_LC_20_11_1 .C_ON=1'b0;
    defparam \ALU.d_RNIPTT4O_8_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPTT4O_8_LC_20_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIPTT4O_8_LC_20_11_1  (
            .in0(N__66703),
            .in1(N__62017),
            .in2(_gnd_net_),
            .in3(N__62209),
            .lcout(\ALU.N_835 ),
            .ltout(\ALU.N_835_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGSBJN2_8_LC_20_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNIGSBJN2_8_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGSBJN2_8_LC_20_11_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.d_RNIGSBJN2_8_LC_20_11_2  (
            .in0(N__66059),
            .in1(N__68929),
            .in2(N__46121),
            .in3(N__46075),
            .lcout(),
            .ltout(\ALU.rshift_7_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIND5CS4_12_LC_20_11_3 .C_ON=1'b0;
    defparam \ALU.c_RNIND5CS4_12_LC_20_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIND5CS4_12_LC_20_11_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.c_RNIND5CS4_12_LC_20_11_3  (
            .in0(N__46118),
            .in1(N__53333),
            .in2(N__46100),
            .in3(N__68926),
            .lcout(),
            .ltout(\ALU.N_925_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIEPHJC7_12_LC_20_11_4 .C_ON=1'b0;
    defparam \ALU.c_RNIEPHJC7_12_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIEPHJC7_12_LC_20_11_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNIEPHJC7_12_LC_20_11_4  (
            .in0(_gnd_net_),
            .in1(N__52685),
            .in2(N__46097),
            .in3(N__45968),
            .lcout(\ALU.a_15_m0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIL9TBN2_6_LC_20_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNIL9TBN2_6_LC_20_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIL9TBN2_6_LC_20_11_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.d_RNIL9TBN2_6_LC_20_11_5  (
            .in0(N__65276),
            .in1(N__68924),
            .in2(N__46094),
            .in3(N__66058),
            .lcout(),
            .ltout(\ALU.rshift_7_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9GG8Q4_8_LC_20_11_6 .C_ON=1'b0;
    defparam \ALU.d_RNI9GG8Q4_8_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9GG8Q4_8_LC_20_11_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI9GG8Q4_8_LC_20_11_6  (
            .in0(N__68925),
            .in1(N__46076),
            .in2(N__46055),
            .in3(N__52705),
            .lcout(\ALU.N_921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI08R632_15_LC_20_11_7 .C_ON=1'b0;
    defparam \ALU.c_RNI08R632_15_LC_20_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI08R632_15_LC_20_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNI08R632_15_LC_20_11_7  (
            .in0(N__70007),
            .in1(N__46032),
            .in2(_gnd_net_),
            .in3(N__45983),
            .lcout(\ALU.c_RNI08R632Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_1_LC_20_12_0 .C_ON=1'b0;
    defparam \ALU.e_1_LC_20_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.e_1_LC_20_12_0 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.e_1_LC_20_12_0  (
            .in0(N__59290),
            .in1(N__69748),
            .in2(N__52246),
            .in3(N__69012),
            .lcout(\ALU.eZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73156),
            .ce(N__69243),
            .sr(_gnd_net_));
    defparam \ALU.e_0_LC_20_12_1 .C_ON=1'b0;
    defparam \ALU.e_0_LC_20_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.e_0_LC_20_12_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.e_0_LC_20_12_1  (
            .in0(N__69170),
            .in1(N__52123),
            .in2(N__69752),
            .in3(N__52033),
            .lcout(\ALU.eZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73156),
            .ce(N__69243),
            .sr(_gnd_net_));
    defparam \ALU.e_7_LC_20_12_2 .C_ON=1'b0;
    defparam \ALU.e_7_LC_20_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.e_7_LC_20_12_2 .LUT_INIT=16'b0101110101011000;
    LogicCell40 \ALU.e_7_LC_20_12_2  (
            .in0(N__58877),
            .in1(N__51904),
            .in2(N__67266),
            .in3(N__51858),
            .lcout(\ALU.eZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73156),
            .ce(N__69243),
            .sr(_gnd_net_));
    defparam \ALU.e_8_LC_20_12_3 .C_ON=1'b0;
    defparam \ALU.e_8_LC_20_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.e_8_LC_20_12_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \ALU.e_8_LC_20_12_3  (
            .in0(N__51727),
            .in1(N__67226),
            .in2(N__51788),
            .in3(N__51638),
            .lcout(\ALU.eZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73156),
            .ce(N__69243),
            .sr(_gnd_net_));
    defparam \ALU.e_15_LC_20_12_4 .C_ON=1'b0;
    defparam \ALU.e_15_LC_20_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.e_15_LC_20_12_4 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.e_15_LC_20_12_4  (
            .in0(N__67225),
            .in1(N__52933),
            .in2(N__59176),
            .in3(N__53006),
            .lcout(\ALU.eZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73156),
            .ce(N__69243),
            .sr(_gnd_net_));
    defparam \ALU.e_9_LC_20_12_5 .C_ON=1'b0;
    defparam \ALU.e_9_LC_20_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.e_9_LC_20_12_5 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \ALU.e_9_LC_20_12_5  (
            .in0(N__52871),
            .in1(N__66843),
            .in2(N__58547),
            .in3(N__52787),
            .lcout(\ALU.eZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73156),
            .ce(N__69243),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIIM1475_12_LC_20_13_0 .C_ON=1'b0;
    defparam \ALU.c_RNIIM1475_12_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIIM1475_12_LC_20_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNIIM1475_12_LC_20_13_0  (
            .in0(N__68812),
            .in1(N__46178),
            .in2(_gnd_net_),
            .in3(N__46159),
            .lcout(\ALU.N_707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_14_c_RNI134CV5_0_LC_20_13_1 .C_ON=1'b0;
    defparam \ALU.addsub_cry_14_c_RNI134CV5_0_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_14_c_RNI134CV5_0_LC_20_13_1 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \ALU.addsub_cry_14_c_RNI134CV5_0_LC_20_13_1  (
            .in0(N__46523),
            .in1(N__63524),
            .in2(N__67255),
            .in3(N__68483),
            .lcout(),
            .ltout(\ALU.addsub_cry_14_c_RNI134CV5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_14_c_RNIKS9S5H_LC_20_13_2 .C_ON=1'b0;
    defparam \ALU.addsub_cry_14_c_RNIKS9S5H_LC_20_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_14_c_RNIKS9S5H_LC_20_13_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.addsub_cry_14_c_RNIKS9S5H_LC_20_13_2  (
            .in0(_gnd_net_),
            .in1(N__46139),
            .in2(N__46133),
            .in3(N__46514),
            .lcout(),
            .ltout(\ALU.addsub_cry_14_c_RNIKS9S5HZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3NTFTL_15_LC_20_13_3 .C_ON=1'b0;
    defparam \ALU.c_RNI3NTFTL_15_LC_20_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3NTFTL_15_LC_20_13_3 .LUT_INIT=16'b0000111000011111;
    LogicCell40 \ALU.c_RNI3NTFTL_15_LC_20_13_3  (
            .in0(N__59338),
            .in1(N__67219),
            .in2(N__46130),
            .in3(N__46565),
            .lcout(\ALU.a_15_1_15 ),
            .ltout(\ALU.a_15_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_LC_20_13_4 .C_ON=1'b0;
    defparam \ALU.a_15_LC_20_13_4 .SEQ_MODE=4'b1000;
    defparam \ALU.a_15_LC_20_13_4 .LUT_INIT=16'b0010111100001101;
    LogicCell40 \ALU.a_15_LC_20_13_4  (
            .in0(N__59169),
            .in1(N__67212),
            .in2(N__46553),
            .in3(N__52987),
            .lcout(\ALU.aZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73162),
            .ce(N__71207),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4MD4S4_2_LC_20_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNI4MD4S4_2_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4MD4S4_2_LC_20_13_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNI4MD4S4_2_LC_20_13_5  (
            .in0(N__46477),
            .in1(N__46500),
            .in2(_gnd_net_),
            .in3(N__68810),
            .lcout(\ALU.N_812 ),
            .ltout(\ALU.N_812_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_14_c_RNI134CV5_LC_20_13_6 .C_ON=1'b0;
    defparam \ALU.addsub_cry_14_c_RNI134CV5_LC_20_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_14_c_RNI134CV5_LC_20_13_6 .LUT_INIT=16'b1100110011110101;
    LogicCell40 \ALU.addsub_cry_14_c_RNI134CV5_LC_20_13_6  (
            .in0(N__68482),
            .in1(N__63523),
            .in2(N__46517),
            .in3(N__67208),
            .lcout(\ALU.addsub_cry_14_c_RNI134CVZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDEP395_2_LC_20_13_7 .C_ON=1'b0;
    defparam \ALU.d_RNIDEP395_2_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDEP395_2_LC_20_13_7 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \ALU.d_RNIDEP395_2_LC_20_13_7  (
            .in0(N__46501),
            .in1(N__68481),
            .in2(N__46481),
            .in3(N__68811),
            .lcout(\ALU.lshift_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_1_LC_20_14_0 .C_ON=1'b0;
    defparam \ALU.c_1_LC_20_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.c_1_LC_20_14_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.c_1_LC_20_14_0  (
            .in0(N__59248),
            .in1(N__52236),
            .in2(N__69678),
            .in3(N__69009),
            .lcout(\ALU.cZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73173),
            .ce(N__71558),
            .sr(_gnd_net_));
    defparam \ALU.c_0_LC_20_14_1 .C_ON=1'b0;
    defparam \ALU.c_0_LC_20_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.c_0_LC_20_14_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.c_0_LC_20_14_1  (
            .in0(N__69149),
            .in1(N__52122),
            .in2(N__69747),
            .in3(N__52049),
            .lcout(\ALU.cZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73173),
            .ce(N__71558),
            .sr(_gnd_net_));
    defparam \ALU.c_7_LC_20_14_2 .C_ON=1'b0;
    defparam \ALU.c_7_LC_20_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.c_7_LC_20_14_2 .LUT_INIT=16'b0111010101100100;
    LogicCell40 \ALU.c_7_LC_20_14_2  (
            .in0(N__58889),
            .in1(N__67273),
            .in2(N__51933),
            .in3(N__51851),
            .lcout(\ALU.cZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73173),
            .ce(N__71558),
            .sr(_gnd_net_));
    defparam \ALU.c_8_LC_20_14_3 .C_ON=1'b0;
    defparam \ALU.c_8_LC_20_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.c_8_LC_20_14_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \ALU.c_8_LC_20_14_3  (
            .in0(N__67271),
            .in1(N__51776),
            .in2(N__51728),
            .in3(N__51633),
            .lcout(\ALU.cZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73173),
            .ce(N__71558),
            .sr(_gnd_net_));
    defparam \ALU.c_15_LC_20_14_4 .C_ON=1'b0;
    defparam \ALU.c_15_LC_20_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.c_15_LC_20_14_4 .LUT_INIT=16'b0111010101000101;
    LogicCell40 \ALU.c_15_LC_20_14_4  (
            .in0(N__52931),
            .in1(N__67272),
            .in2(N__59177),
            .in3(N__53009),
            .lcout(\ALU.cZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73173),
            .ce(N__71558),
            .sr(_gnd_net_));
    defparam \ALU.c_9_LC_20_14_5 .C_ON=1'b0;
    defparam \ALU.c_9_LC_20_14_5 .SEQ_MODE=4'b1000;
    defparam \ALU.c_9_LC_20_14_5 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \ALU.c_9_LC_20_14_5  (
            .in0(N__58524),
            .in1(N__52879),
            .in2(N__52807),
            .in3(N__66833),
            .lcout(\ALU.cZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73173),
            .ce(N__71558),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI500DG_7_LC_20_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNI500DG_7_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI500DG_7_LC_20_15_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ALU.d_RNI500DG_7_LC_20_15_0  (
            .in0(N__55886),
            .in1(N__63217),
            .in2(_gnd_net_),
            .in3(N__62158),
            .lcout(\ALU.d_RNI500DGZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5KAEG_7_LC_20_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNI5KAEG_7_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5KAEG_7_LC_20_15_1 .LUT_INIT=16'b0011011011101000;
    LogicCell40 \ALU.d_RNI5KAEG_7_LC_20_15_1  (
            .in0(N__62157),
            .in1(N__74778),
            .in2(N__63273),
            .in3(N__55887),
            .lcout(\ALU.log_1_7 ),
            .ltout(\ALU.log_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_492_c_RNIQ5B457_LC_20_15_2 .C_ON=1'b0;
    defparam \ALU.mult_492_c_RNIQ5B457_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_492_c_RNIQ5B457_LC_20_15_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.mult_492_c_RNIQ5B457_LC_20_15_2  (
            .in0(_gnd_net_),
            .in1(N__59100),
            .in2(N__46643),
            .in3(N__46640),
            .lcout(),
            .ltout(\ALU.mult_492_c_RNIQ5BZ0Z457_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_492_c_RNIGN2JEC_LC_20_15_3 .C_ON=1'b0;
    defparam \ALU.mult_492_c_RNIGN2JEC_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_492_c_RNIGN2JEC_LC_20_15_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \ALU.mult_492_c_RNIGN2JEC_LC_20_15_3  (
            .in0(N__59101),
            .in1(N__70096),
            .in2(N__46625),
            .in3(N__46622),
            .lcout(\ALU.mult_492_c_RNIGN2JECZ0 ),
            .ltout(\ALU.mult_492_c_RNIGN2JECZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_7_LC_20_15_4 .C_ON=1'b0;
    defparam \ALU.a_7_LC_20_15_4 .SEQ_MODE=4'b1000;
    defparam \ALU.a_7_LC_20_15_4 .LUT_INIT=16'b0111011000110010;
    LogicCell40 \ALU.a_7_LC_20_15_4  (
            .in0(N__67230),
            .in1(N__58887),
            .in2(N__46613),
            .in3(N__51932),
            .lcout(\ALU.aZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73184),
            .ce(N__71176),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO75BG_7_LC_20_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNIO75BG_7_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO75BG_7_LC_20_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIO75BG_7_LC_20_15_5  (
            .in0(N__62156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55885),
            .lcout(\ALU.d_RNIO75BGZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_d_d_s_0_LC_20_15_6 .C_ON=1'b0;
    defparam \ALU.a_15_m2_d_d_s_0_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_d_d_s_0_LC_20_15_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \ALU.a_15_m2_d_d_s_0_LC_20_15_6  (
            .in0(N__70095),
            .in1(N__69790),
            .in2(_gnd_net_),
            .in3(N__63218),
            .lcout(\ALU.a_15_m2_d_d_sZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2s2_i_LC_20_15_7 .C_ON=1'b0;
    defparam \ALU.a_15_m2s2_i_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2s2_i_LC_20_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.a_15_m2s2_i_LC_20_15_7  (
            .in0(_gnd_net_),
            .in1(N__69789),
            .in2(_gnd_net_),
            .in3(N__70094),
            .lcout(\ALU.a_15_sm0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI9SHF_14_LC_20_16_0 .C_ON=1'b0;
    defparam \ALU.c_RNI9SHF_14_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI9SHF_14_LC_20_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNI9SHF_14_LC_20_16_0  (
            .in0(N__52291),
            .in1(N__67312),
            .in2(_gnd_net_),
            .in3(N__46923),
            .lcout(\ALU.c_RNI9SHFZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_s_1_LC_20_16_1 .C_ON=1'b0;
    defparam \ALU.a_15_m2_s_1_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_s_1_LC_20_16_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ALU.a_15_m2_s_1_LC_20_16_1  (
            .in0(N__69972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59262),
            .lcout(\ALU.a_15_m2_sZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPNGFE_14_LC_20_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNIPNGFE_14_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPNGFE_14_LC_20_16_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \ALU.d_RNIPNGFE_14_LC_20_16_3  (
            .in0(N__53306),
            .in1(N__47062),
            .in2(N__46697),
            .in3(N__49581),
            .lcout(\ALU.status_19_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI5CPU_14_LC_20_16_4 .C_ON=1'b0;
    defparam \ALU.a_RNI5CPU_14_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI5CPU_14_LC_20_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.a_RNI5CPU_14_LC_20_16_4  (
            .in0(N__52447),
            .in1(N__57454),
            .in2(_gnd_net_),
            .in3(N__46924),
            .lcout(),
            .ltout(\ALU.a_RNI5CPUZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINT5A2_14_LC_20_16_5 .C_ON=1'b0;
    defparam \ALU.c_RNINT5A2_14_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINT5A2_14_LC_20_16_5 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.c_RNINT5A2_14_LC_20_16_5  (
            .in0(N__46850),
            .in1(N__53938),
            .in2(N__46844),
            .in3(N__46827),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFU325_14_LC_20_16_6 .C_ON=1'b0;
    defparam \ALU.d_RNIFU325_14_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFU325_14_LC_20_16_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIFU325_14_LC_20_16_6  (
            .in0(N__53939),
            .in1(N__46733),
            .in2(N__46724),
            .in3(N__46721),
            .lcout(),
            .ltout(\ALU.operand2_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINISC7_14_LC_20_16_7 .C_ON=1'b0;
    defparam \ALU.d_RNINISC7_14_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINISC7_14_LC_20_16_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.d_RNINISC7_14_LC_20_16_7  (
            .in0(_gnd_net_),
            .in1(N__46712),
            .in2(N__46700),
            .in3(N__71454),
            .lcout(\ALU.d_RNINISC7Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI80U51_14_LC_20_17_0 .C_ON=1'b0;
    defparam \ALU.a_RNI80U51_14_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI80U51_14_LC_20_17_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.a_RNI80U51_14_LC_20_17_0  (
            .in0(N__57458),
            .in1(N__47275),
            .in2(N__52451),
            .in3(N__54298),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIG4FM1_14_LC_20_17_1 .C_ON=1'b0;
    defparam \ALU.c_RNIG4FM1_14_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIG4FM1_14_LC_20_17_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.c_RNIG4FM1_14_LC_20_17_1  (
            .in0(N__67313),
            .in1(N__52284),
            .in2(N__46688),
            .in3(N__47192),
            .lcout(\ALU.N_1099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIA8AE1_14_LC_20_17_2 .C_ON=1'b0;
    defparam \ALU.b_RNIA8AE1_14_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIA8AE1_14_LC_20_17_2 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNIA8AE1_14_LC_20_17_2  (
            .in0(N__67963),
            .in1(N__47274),
            .in2(N__57586),
            .in3(N__54299),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKK772_14_LC_20_17_3 .C_ON=1'b0;
    defparam \ALU.d_RNIKK772_14_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKK772_14_LC_20_17_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.d_RNIKK772_14_LC_20_17_3  (
            .in0(N__67784),
            .in1(N__57859),
            .in2(N__47216),
            .in3(N__47193),
            .lcout(),
            .ltout(\ALU.N_1147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI7T474_14_LC_20_17_4 .C_ON=1'b0;
    defparam \ALU.c_RNI7T474_14_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI7T474_14_LC_20_17_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.c_RNI7T474_14_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(N__47099),
            .in2(N__47093),
            .in3(N__54139),
            .lcout(aluOut_14),
            .ltout(aluOut_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI51G56_1_LC_20_17_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI51G56_1_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI51G56_1_LC_20_17_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \CONTROL.busState_1_RNI51G56_1_LC_20_17_5  (
            .in0(N__47090),
            .in1(N__50325),
            .in2(N__47075),
            .in3(N__50214),
            .lcout(N_207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.increment_1_LC_20_18_0 .C_ON=1'b0;
    defparam \CONTROL.increment_1_LC_20_18_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.increment_1_LC_20_18_0 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \CONTROL.increment_1_LC_20_18_0  (
            .in0(N__47051),
            .in1(N__47011),
            .in2(N__46964),
            .in3(N__54686),
            .lcout(\CONTROL.incrementZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.increment_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIH85J_0_LC_20_18_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIH85J_0_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIH85J_0_LC_20_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIH85J_0_LC_20_18_1  (
            .in0(N__55079),
            .in1(N__50990),
            .in2(_gnd_net_),
            .in3(N__47615),
            .lcout(N_415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m399_bm_LC_20_18_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m399_bm_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m399_bm_LC_20_18_2 .LUT_INIT=16'b0010000000000100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m399_bm_LC_20_18_2  (
            .in0(N__78027),
            .in1(N__78823),
            .in2(N__75994),
            .in3(N__77296),
            .lcout(\PROM.ROMDATA.m399_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m422_am_LC_20_18_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m422_am_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m422_am_LC_20_18_3 .LUT_INIT=16'b0011100000100100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m422_am_LC_20_18_3  (
            .in0(N__77297),
            .in1(N__75938),
            .in2(N__78862),
            .in3(N__78028),
            .lcout(\PROM.ROMDATA.m422_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m422_bm_LC_20_18_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m422_bm_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m422_bm_LC_20_18_4 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m422_bm_LC_20_18_4  (
            .in0(N__75939),
            .in1(N__64863),
            .in2(_gnd_net_),
            .in3(N__78827),
            .lcout(),
            .ltout(\PROM.ROMDATA.m422_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m422_ns_LC_20_18_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m422_ns_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m422_ns_LC_20_18_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m422_ns_LC_20_18_5  (
            .in0(_gnd_net_),
            .in1(N__47372),
            .in2(N__47366),
            .in3(N__76587),
            .lcout(\PROM.ROMDATA.m422_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m381_bm_LC_20_18_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m381_bm_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m381_bm_LC_20_18_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m381_bm_LC_20_18_6  (
            .in0(N__75940),
            .in1(N__50447),
            .in2(N__76623),
            .in3(N__64254),
            .lcout(\PROM.ROMDATA.m381_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m482_LC_20_18_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m482_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m482_LC_20_18_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m482_LC_20_18_7  (
            .in0(N__78828),
            .in1(N__47514),
            .in2(N__64875),
            .in3(N__75941),
            .lcout(\PROM.ROMDATA.N_551_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m298_ns_LC_20_19_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m298_ns_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m298_ns_LC_20_19_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m298_ns_LC_20_19_0  (
            .in0(N__47345),
            .in1(N__64031),
            .in2(_gnd_net_),
            .in3(N__76483),
            .lcout(\PROM.ROMDATA.m298_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_RNIMGJ31_4_LC_20_19_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_RNIMGJ31_4_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_36_RNIMGJ31_4_LC_20_19_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \CONTROL.programCounter_ret_36_RNIMGJ31_4_LC_20_19_1  (
            .in0(N__73721),
            .in1(_gnd_net_),
            .in2(N__47681),
            .in3(N__55168),
            .lcout(\CONTROL.programCounter_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m35_1_LC_20_19_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m35_1_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m35_1_LC_20_19_3 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m35_1_LC_20_19_3  (
            .in0(N__76482),
            .in1(N__47726),
            .in2(N__50645),
            .in3(N__79761),
            .lcout(\PROM.ROMDATA.m35_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m498_bm_LC_20_19_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m498_bm_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m498_bm_LC_20_19_4 .LUT_INIT=16'b0101110011010111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m498_bm_LC_20_19_4  (
            .in0(N__78830),
            .in1(N__77932),
            .in2(N__77314),
            .in3(N__75934),
            .lcout(\PROM.ROMDATA.m498_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m124_e_LC_20_19_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m124_e_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m124_e_LC_20_19_5 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m124_e_LC_20_19_5  (
            .in0(N__73720),
            .in1(N__79762),
            .in2(N__47680),
            .in3(N__55167),
            .lcout(\PROM.ROMDATA.N_543_mux_2 ),
            .ltout(\PROM.ROMDATA.N_543_mux_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m176_LC_20_19_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m176_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m176_LC_20_19_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m176_LC_20_19_6  (
            .in0(N__64323),
            .in1(N__79293),
            .in2(N__47312),
            .in3(N__75932),
            .lcout(\PROM.ROMDATA.N_559_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m392_am_LC_20_19_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m392_am_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m392_am_LC_20_19_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m392_am_LC_20_19_7  (
            .in0(N__75933),
            .in1(N__78829),
            .in2(N__64324),
            .in3(N__78980),
            .lcout(\PROM.ROMDATA.m392_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m163_LC_20_20_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m163_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m163_LC_20_20_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m163_LC_20_20_0  (
            .in0(N__77198),
            .in1(_gnd_net_),
            .in2(N__77994),
            .in3(N__78730),
            .lcout(\PROM.ROMDATA.m163 ),
            .ltout(\PROM.ROMDATA.m163_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m176_x_LC_20_20_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m176_x_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m176_x_LC_20_20_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m176_x_LC_20_20_1  (
            .in0(N__75247),
            .in1(_gnd_net_),
            .in2(N__47540),
            .in3(N__79208),
            .lcout(\PROM.ROMDATA.m176_x ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m474_LC_20_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m474_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m474_LC_20_20_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m474_LC_20_20_2  (
            .in0(N__79209),
            .in1(N__75248),
            .in2(N__47523),
            .in3(N__64965),
            .lcout(\PROM.ROMDATA.N_569_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m109_am_1_LC_20_20_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m109_am_1_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m109_am_1_LC_20_20_3 .LUT_INIT=16'b0011000101000110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m109_am_1_LC_20_20_3  (
            .in0(N__78727),
            .in1(N__77842),
            .in2(N__75539),
            .in3(N__77196),
            .lcout(),
            .ltout(\PROM.ROMDATA.m109_am_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m109_am_LC_20_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m109_am_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m109_am_LC_20_20_4 .LUT_INIT=16'b0100111101101111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m109_am_LC_20_20_4  (
            .in0(N__76479),
            .in1(N__75243),
            .in2(N__47429),
            .in3(N__78729),
            .lcout(\PROM.ROMDATA.m109_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m11_am_LC_20_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m11_am_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m11_am_LC_20_20_5 .LUT_INIT=16'b1100110110011110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m11_am_LC_20_20_5  (
            .in0(N__78728),
            .in1(N__77843),
            .in2(N__75540),
            .in3(N__77197),
            .lcout(\PROM.ROMDATA.m11_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_0_LC_20_20_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_0_LC_20_20_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_0_LC_20_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_0_LC_20_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47426),
            .lcout(CONTROL_addrstack_reto_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73225),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_0_LC_20_20_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_0_LC_20_20_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_0_LC_20_20_7 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \CONTROL.programCounter_ret_1_0_LC_20_20_7  (
            .in0(N__47403),
            .in1(N__73712),
            .in2(_gnd_net_),
            .in3(N__50955),
            .lcout(\CONTROL.programCounter_1_reto_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73225),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIPG5J_4_LC_20_21_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIPG5J_4_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIPG5J_4_LC_20_21_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIPG5J_4_LC_20_21_0  (
            .in0(N__55057),
            .in1(N__55183),
            .in2(_gnd_net_),
            .in3(N__55301),
            .lcout(N_419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_1_LC_20_21_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_1_LC_20_21_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_1_LC_20_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_1_LC_20_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47660),
            .lcout(CONTROL_addrstack_reto_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73237),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_RNIEO8J_3_LC_20_21_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_RNIEO8J_3_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_19_RNIEO8J_3_LC_20_21_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.programCounter_ret_19_RNIEO8J_3_LC_20_21_2  (
            .in0(N__55120),
            .in1(N__47635),
            .in2(_gnd_net_),
            .in3(N__64465),
            .lcout(\CONTROL.programCounter_ret_19_RNIEO8JZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNILA8I_3_LC_20_21_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNILA8I_3_LC_20_21_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNILA8I_3_LC_20_21_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CONTROL.programCounter_ret_1_RNILA8I_3_LC_20_21_3  (
            .in0(N__64466),
            .in1(N__51121),
            .in2(_gnd_net_),
            .in3(N__55119),
            .lcout(),
            .ltout(\CONTROL.programCounter_ret_1_RNILA8IZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_fast_RNI93CH1_LC_20_21_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_fast_RNI93CH1_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_18_fast_RNI93CH1_LC_20_21_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \CONTROL.programCounter_ret_18_fast_RNI93CH1_LC_20_21_4  (
            .in0(N__55056),
            .in1(_gnd_net_),
            .in2(N__47624),
            .in3(N__47621),
            .lcout(progRomAddress_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIF48I_0_LC_20_21_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIF48I_0_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIF48I_0_LC_20_21_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIF48I_0_LC_20_21_5  (
            .in0(N__47611),
            .in1(N__55118),
            .in2(_gnd_net_),
            .in3(N__50947),
            .lcout(\CONTROL.programCounter_ret_1_RNIF48IZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_3_LC_20_21_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_3_LC_20_21_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_3_LC_20_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_3_LC_20_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47600),
            .lcout(CONTROL_addrstack_reto_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73237),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m35_LC_20_22_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m35_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m35_LC_20_22_0 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m35_LC_20_22_0  (
            .in0(N__47588),
            .in1(N__47582),
            .in2(N__54923),
            .in3(N__79715),
            .lcout(\PROM.ROMDATA.m35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIJ88I_2_LC_20_22_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIJ88I_2_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIJ88I_2_LC_20_22_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIJ88I_2_LC_20_22_1  (
            .in0(N__47563),
            .in1(N__64692),
            .in2(_gnd_net_),
            .in3(N__55123),
            .lcout(\CONTROL.programCounter_ret_1_RNIJ88IZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_1_LC_20_22_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_1_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_1_LC_20_22_2 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_1_LC_20_22_2  (
            .in0(N__75291),
            .in1(N__78625),
            .in2(_gnd_net_),
            .in3(N__77613),
            .lcout(),
            .ltout(\PROM.ROMDATA.m215_ns_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_LC_20_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_LC_20_22_3 .LUT_INIT=16'b0010111101111001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_LC_20_22_3  (
            .in0(N__77114),
            .in1(N__76499),
            .in2(N__47717),
            .in3(N__75292),
            .lcout(\PROM.ROMDATA.m215_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m178_LC_20_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m178_LC_20_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m178_LC_20_22_4 .LUT_INIT=16'b0001000110001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m178_LC_20_22_4  (
            .in0(N__78636),
            .in1(N__77615),
            .in2(_gnd_net_),
            .in3(N__77116),
            .lcout(\PROM.ROMDATA.m178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_RNICM8J_2_LC_20_22_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_RNICM8J_2_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_19_RNICM8J_2_LC_20_22_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_19_RNICM8J_2_LC_20_22_5  (
            .in0(N__54802),
            .in1(N__64693),
            .in2(_gnd_net_),
            .in3(N__55124),
            .lcout(\CONTROL.programCounter_ret_19_RNICM8JZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m256_LC_20_22_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m256_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m256_LC_20_22_6 .LUT_INIT=16'b0000100000110010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m256_LC_20_22_6  (
            .in0(N__78635),
            .in1(N__77614),
            .in2(N__75613),
            .in3(N__77115),
            .lcout(\PROM.ROMDATA.m256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_35_fast_LC_20_22_7 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_35_fast_LC_20_22_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_35_fast_LC_20_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \CONTROL.programCounter_ret_35_fast_LC_20_22_7  (
            .in0(_gnd_net_),
            .in1(N__50834),
            .in2(_gnd_net_),
            .in3(N__50898),
            .lcout(\CONTROL.programCounter11_reto_fast ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73247),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m38_LC_20_23_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m38_LC_20_23_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m38_LC_20_23_0 .LUT_INIT=16'b0111101101101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m38_LC_20_23_0  (
            .in0(N__77620),
            .in1(N__78688),
            .in2(N__75919),
            .in3(N__76937),
            .lcout(\PROM.ROMDATA.m38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m251_LC_20_23_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m251_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m251_LC_20_23_1 .LUT_INIT=16'b0100010100111000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m251_LC_20_23_1  (
            .in0(N__76933),
            .in1(N__78692),
            .in2(N__75912),
            .in3(N__77618),
            .lcout(\PROM.ROMDATA.m251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m253_LC_20_23_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m253_LC_20_23_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m253_LC_20_23_2 .LUT_INIT=16'b0100101000101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m253_LC_20_23_2  (
            .in0(N__77617),
            .in1(N__75726),
            .in2(N__78833),
            .in3(N__76934),
            .lcout(\PROM.ROMDATA.m253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m389_bm_LC_20_23_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m389_bm_LC_20_23_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m389_bm_LC_20_23_3 .LUT_INIT=16'b0000010000000010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m389_bm_LC_20_23_3  (
            .in0(N__76936),
            .in1(N__78693),
            .in2(N__75913),
            .in3(N__77619),
            .lcout(\PROM.ROMDATA.m389_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m20_LC_20_23_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m20_LC_20_23_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m20_LC_20_23_4 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m20_LC_20_23_4  (
            .in0(N__64741),
            .in1(N__64698),
            .in2(N__64641),
            .in3(N__76932),
            .lcout(\PROM.ROMDATA.m20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_6_LC_20_23_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_6_LC_20_23_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_6_LC_20_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_1_6_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47846),
            .lcout(\CONTROL.programCounter_1_reto_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73257),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m51_LC_20_23_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m51_LC_20_23_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m51_LC_20_23_6 .LUT_INIT=16'b0010011110110001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m51_LC_20_23_6  (
            .in0(N__77616),
            .in1(N__78687),
            .in2(N__75918),
            .in3(N__76935),
            .lcout(\PROM.ROMDATA.m51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m433_am_LC_20_23_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m433_am_LC_20_23_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m433_am_LC_20_23_7 .LUT_INIT=16'b0101000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m433_am_LC_20_23_7  (
            .in0(N__76528),
            .in1(N__74447),
            .in2(N__73373),
            .in3(N__75750),
            .lcout(\PROM.ROMDATA.m433_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m399_am_LC_20_24_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m399_am_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m399_am_LC_20_24_0 .LUT_INIT=16'b0000000011010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m399_am_LC_20_24_0  (
            .in0(N__77874),
            .in1(N__75383),
            .in2(N__64861),
            .in3(N__78639),
            .lcout(),
            .ltout(\PROM.ROMDATA.m399_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m399_ns_LC_20_24_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m399_ns_LC_20_24_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m399_ns_LC_20_24_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m399_ns_LC_20_24_1  (
            .in0(_gnd_net_),
            .in1(N__76529),
            .in2(N__47786),
            .in3(N__47783),
            .lcout(\PROM.ROMDATA.m399_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m461_ns_1_LC_20_24_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m461_ns_1_LC_20_24_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m461_ns_1_LC_20_24_2 .LUT_INIT=16'b0111011101000111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m461_ns_1_LC_20_24_2  (
            .in0(N__64199),
            .in1(N__79391),
            .in2(N__47906),
            .in3(N__79850),
            .lcout(\PROM.ROMDATA.m461_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_36_4_LC_20_24_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_36_4_LC_20_24_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_36_4_LC_20_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_36_4_LC_20_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47744),
            .lcout(CONTROL_addrstack_reto_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73266),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m22_LC_20_24_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m22_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m22_LC_20_24_5 .LUT_INIT=16'b0101110000010011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m22_LC_20_24_5  (
            .in0(N__78638),
            .in1(N__77873),
            .in2(N__75676),
            .in3(N__77184),
            .lcout(\PROM.ROMDATA.m22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m451_bm_LC_20_24_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m451_bm_LC_20_24_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m451_bm_LC_20_24_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m451_bm_LC_20_24_6  (
            .in0(N__64837),
            .in1(N__75384),
            .in2(N__73892),
            .in3(N__78640),
            .lcout(),
            .ltout(\PROM.ROMDATA.m451_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m451_ns_LC_20_24_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m451_ns_LC_20_24_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m451_ns_LC_20_24_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m451_ns_LC_20_24_7  (
            .in0(_gnd_net_),
            .in1(N__76530),
            .in2(N__47918),
            .in3(N__47915),
            .lcout(\PROM.ROMDATA.m451_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m375_bm_LC_20_25_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m375_bm_LC_20_25_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m375_bm_LC_20_25_0 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m375_bm_LC_20_25_0  (
            .in0(N__47873),
            .in1(N__76527),
            .in2(N__74285),
            .in3(N__75790),
            .lcout(\PROM.ROMDATA.m375_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m280_LC_20_25_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m280_LC_20_25_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m280_LC_20_25_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m280_LC_20_25_1  (
            .in0(N__78994),
            .in1(N__75791),
            .in2(N__76602),
            .in3(N__78695),
            .lcout(\PROM.ROMDATA.m280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m376_LC_20_25_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m376_LC_20_25_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m376_LC_20_25_2 .LUT_INIT=16'b0001001010010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m376_LC_20_25_2  (
            .in0(N__77882),
            .in1(N__75789),
            .in2(N__78835),
            .in3(N__77192),
            .lcout(\PROM.ROMDATA.m376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m255_LC_20_25_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m255_LC_20_25_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m255_LC_20_25_4 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m255_LC_20_25_4  (
            .in0(N__77881),
            .in1(_gnd_net_),
            .in2(N__78834),
            .in3(N__77190),
            .lcout(\PROM.ROMDATA.N_256_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m389_am_LC_20_25_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m389_am_LC_20_25_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m389_am_LC_20_25_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m389_am_LC_20_25_5  (
            .in0(N__78993),
            .in1(N__78696),
            .in2(N__75950),
            .in3(N__77880),
            .lcout(),
            .ltout(\PROM.ROMDATA.m389_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m389_ns_LC_20_25_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m389_ns_LC_20_25_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m389_ns_LC_20_25_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m389_ns_LC_20_25_6  (
            .in0(_gnd_net_),
            .in1(N__47867),
            .in2(N__47858),
            .in3(N__76526),
            .lcout(\PROM.ROMDATA.m389_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m103_LC_20_25_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m103_LC_20_25_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m103_LC_20_25_7 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m103_LC_20_25_7  (
            .in0(N__77191),
            .in1(N__78700),
            .in2(_gnd_net_),
            .in3(N__77883),
            .lcout(\PROM.ROMDATA.m103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIMNQ8E1_0_12_LC_21_9_0 .C_ON=1'b0;
    defparam \ALU.c_RNIMNQ8E1_0_12_LC_21_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIMNQ8E1_0_12_LC_21_9_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.c_RNIMNQ8E1_0_12_LC_21_9_0  (
            .in0(N__61010),
            .in1(N__66063),
            .in2(N__61225),
            .in3(N__66757),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIUU8GB2_10_LC_21_9_1 .C_ON=1'b0;
    defparam \ALU.c_RNIUU8GB2_10_LC_21_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIUU8GB2_10_LC_21_9_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNIUU8GB2_10_LC_21_9_1  (
            .in0(N__66064),
            .in1(N__61640),
            .in2(N__48092),
            .in3(N__61474),
            .lcout(),
            .ltout(\ALU.N_645_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI5G4OF5_10_LC_21_9_2 .C_ON=1'b0;
    defparam \ALU.c_RNI5G4OF5_10_LC_21_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI5G4OF5_10_LC_21_9_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.c_RNI5G4OF5_10_LC_21_9_2  (
            .in0(N__68918),
            .in1(N__68511),
            .in2(N__48089),
            .in3(N__48032),
            .lcout(),
            .ltout(\ALU.a_15_m1_am_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRFBHE9_0_LC_21_9_3 .C_ON=1'b0;
    defparam \ALU.d_RNIRFBHE9_0_LC_21_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRFBHE9_0_LC_21_9_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.d_RNIRFBHE9_0_LC_21_9_3  (
            .in0(N__48016),
            .in1(N__48086),
            .in2(N__48065),
            .in3(N__68510),
            .lcout(\ALU.d_RNIRFBHE9Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBK47O_0_8_LC_21_9_4 .C_ON=1'b0;
    defparam \ALU.d_RNIBK47O_0_8_LC_21_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBK47O_0_8_LC_21_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIBK47O_0_8_LC_21_9_4  (
            .in0(N__62023),
            .in1(N__62885),
            .in2(_gnd_net_),
            .in3(N__66756),
            .lcout(),
            .ltout(\ALU.N_611_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMQD952_8_LC_21_9_5 .C_ON=1'b0;
    defparam \ALU.d_RNIMQD952_8_LC_21_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMQD952_8_LC_21_9_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNIMQD952_8_LC_21_9_5  (
            .in0(N__66062),
            .in1(_gnd_net_),
            .in2(N__48062),
            .in3(N__48058),
            .lcout(\ALU.N_641 ),
            .ltout(\ALU.N_641_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITG2137_0_LC_21_9_6 .C_ON=1'b0;
    defparam \ALU.d_RNITG2137_0_LC_21_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITG2137_0_LC_21_9_6 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \ALU.d_RNITG2137_0_LC_21_9_6  (
            .in0(N__68509),
            .in1(N__47942),
            .in2(N__48026),
            .in3(N__48015),
            .lcout(\ALU.d_RNITG2137Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQGO2C2_0_LC_21_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNIQGO2C2_0_LC_21_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQGO2C2_0_LC_21_9_7 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \ALU.d_RNIQGO2C2_0_LC_21_9_7  (
            .in0(N__66061),
            .in1(N__68508),
            .in2(N__47990),
            .in3(N__68917),
            .lcout(\ALU.a_15_m1_am_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0OR9G_3_LC_21_10_5 .C_ON=1'b0;
    defparam \ALU.d_RNI0OR9G_3_LC_21_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0OR9G_3_LC_21_10_5 .LUT_INIT=16'b1110000100010111;
    LogicCell40 \ALU.d_RNI0OR9G_3_LC_21_10_5  (
            .in0(N__63253),
            .in1(N__60260),
            .in2(N__74816),
            .in3(N__68490),
            .lcout(\ALU.a_15_m3_d_d_0_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBRG4Q9_0_12_LC_21_11_0 .C_ON=1'b0;
    defparam \ALU.c_RNIBRG4Q9_0_12_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBRG4Q9_0_12_LC_21_11_0 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \ALU.c_RNIBRG4Q9_0_12_LC_21_11_0  (
            .in0(N__58497),
            .in1(N__70171),
            .in2(N__48188),
            .in3(N__48175),
            .lcout(\ALU.c_RNIBRG4Q9_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_555_c_RNIJF56AM_LC_21_11_1 .C_ON=1'b0;
    defparam \ALU.mult_555_c_RNIJF56AM_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_555_c_RNIJF56AM_LC_21_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.mult_555_c_RNIJF56AM_LC_21_11_1  (
            .in0(N__69640),
            .in1(N__48290),
            .in2(_gnd_net_),
            .in3(N__48506),
            .lcout(\ALU.mult_555_c_RNIJF56AMZ0 ),
            .ltout(\ALU.mult_555_c_RNIJF56AMZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_12_LC_21_11_2 .C_ON=1'b0;
    defparam \ALU.a_12_LC_21_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.a_12_LC_21_11_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \ALU.a_12_LC_21_11_2  (
            .in0(_gnd_net_),
            .in1(N__67742),
            .in2(N__48272),
            .in3(N__67654),
            .lcout(\ALU.aZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73157),
            .ce(N__71197),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI5SENO2_12_LC_21_11_3 .C_ON=1'b0;
    defparam \ALU.c_RNI5SENO2_12_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI5SENO2_12_LC_21_11_3 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.c_RNI5SENO2_12_LC_21_11_3  (
            .in0(N__48236),
            .in1(N__68927),
            .in2(N__48212),
            .in3(N__66060),
            .lcout(),
            .ltout(\ALU.lshift_7_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3I5IR4_8_LC_21_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNI3I5IR4_8_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3I5IR4_8_LC_21_11_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI3I5IR4_8_LC_21_11_4  (
            .in0(N__68928),
            .in1(N__48677),
            .in2(N__48194),
            .in3(N__48710),
            .lcout(),
            .ltout(\ALU.N_704_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGNBT49_8_LC_21_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNIGNBT49_8_LC_21_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGNBT49_8_LC_21_11_5 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \ALU.d_RNIGNBT49_8_LC_21_11_5  (
            .in0(N__70169),
            .in1(N__48535),
            .in2(N__48191),
            .in3(N__68484),
            .lcout(\ALU.d_RNIGNBT49Z0Z_8 ),
            .ltout(\ALU.d_RNIGNBT49Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBRG4Q9_12_LC_21_11_6 .C_ON=1'b0;
    defparam \ALU.c_RNIBRG4Q9_12_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBRG4Q9_12_LC_21_11_6 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \ALU.c_RNIBRG4Q9_12_LC_21_11_6  (
            .in0(N__58496),
            .in1(N__70170),
            .in2(N__48179),
            .in3(N__48174),
            .lcout(\ALU.c_RNIBRG4Q9Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_8_LC_21_12_0 .C_ON=1'b0;
    defparam \ALU.h_8_LC_21_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_8_LC_21_12_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \ALU.h_8_LC_21_12_0  (
            .in0(N__67231),
            .in1(N__51784),
            .in2(N__51723),
            .in3(N__51637),
            .lcout(h_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73163),
            .ce(N__69452),
            .sr(_gnd_net_));
    defparam \ALU.h_15_LC_21_12_1 .C_ON=1'b0;
    defparam \ALU.h_15_LC_21_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.h_15_LC_21_12_1 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.h_15_LC_21_12_1  (
            .in0(N__67207),
            .in1(N__52934),
            .in2(N__59140),
            .in3(N__53012),
            .lcout(h_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73163),
            .ce(N__69452),
            .sr(_gnd_net_));
    defparam \ALU.mult_555_c_RNI5VJUOI_LC_21_12_2 .C_ON=1'b0;
    defparam \ALU.mult_555_c_RNI5VJUOI_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_555_c_RNI5VJUOI_LC_21_12_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.mult_555_c_RNI5VJUOI_LC_21_12_2  (
            .in0(N__61042),
            .in1(N__67205),
            .in2(_gnd_net_),
            .in3(N__48518),
            .lcout(\ALU.mult_555_c_RNI5VJUOIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_546_c_RNIJOT4J8_LC_21_12_4 .C_ON=1'b0;
    defparam \ALU.mult_546_c_RNIJOT4J8_LC_21_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_546_c_RNIJOT4J8_LC_21_12_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ALU.mult_546_c_RNIJOT4J8_LC_21_12_4  (
            .in0(N__66896),
            .in1(N__67206),
            .in2(_gnd_net_),
            .in3(N__48500),
            .lcout(\ALU.mult_546_c_RNIJOT4JZ0Z8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_3_0_LC_21_12_5 .C_ON=1'b0;
    defparam \ALU.status_RNO_3_0_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_3_0_LC_21_12_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ALU.status_RNO_3_0_LC_21_12_5  (
            .in0(N__61277),
            .in1(N__60839),
            .in2(N__53360),
            .in3(N__61043),
            .lcout(),
            .ltout(\ALU.status_14_12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_1_0_LC_21_12_6 .C_ON=1'b0;
    defparam \ALU.status_RNO_1_0_LC_21_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_1_0_LC_21_12_6 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \ALU.status_RNO_1_0_LC_21_12_6  (
            .in0(N__69512),
            .in1(N__48487),
            .in2(N__48428),
            .in3(N__53342),
            .lcout(\ALU.status_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_1_LC_21_13_0 .C_ON=1'b0;
    defparam \ALU.b_1_LC_21_13_0 .SEQ_MODE=4'b1000;
    defparam \ALU.b_1_LC_21_13_0 .LUT_INIT=16'b0100111000001111;
    LogicCell40 \ALU.b_1_LC_21_13_0  (
            .in0(N__59306),
            .in1(N__69002),
            .in2(N__52245),
            .in3(N__69729),
            .lcout(\ALU.bZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73174),
            .ce(N__67931),
            .sr(_gnd_net_));
    defparam \ALU.b_0_LC_21_13_1 .C_ON=1'b0;
    defparam \ALU.b_0_LC_21_13_1 .SEQ_MODE=4'b1000;
    defparam \ALU.b_0_LC_21_13_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.b_0_LC_21_13_1  (
            .in0(N__69169),
            .in1(N__52118),
            .in2(N__69744),
            .in3(N__52050),
            .lcout(\ALU.bZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73174),
            .ce(N__67931),
            .sr(_gnd_net_));
    defparam \ALU.b_7_LC_21_13_2 .C_ON=1'b0;
    defparam \ALU.b_7_LC_21_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.b_7_LC_21_13_2 .LUT_INIT=16'b0111011001010100;
    LogicCell40 \ALU.b_7_LC_21_13_2  (
            .in0(N__58888),
            .in1(N__67218),
            .in2(N__51863),
            .in3(N__51930),
            .lcout(\ALU.bZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73174),
            .ce(N__67931),
            .sr(_gnd_net_));
    defparam \ALU.b_8_LC_21_13_3 .C_ON=1'b0;
    defparam \ALU.b_8_LC_21_13_3 .SEQ_MODE=4'b1000;
    defparam \ALU.b_8_LC_21_13_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \ALU.b_8_LC_21_13_3  (
            .in0(N__67217),
            .in1(N__51775),
            .in2(N__51720),
            .in3(N__51632),
            .lcout(\ALU.bZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73174),
            .ce(N__67931),
            .sr(_gnd_net_));
    defparam \ALU.b_15_LC_21_13_4 .C_ON=1'b0;
    defparam \ALU.b_15_LC_21_13_4 .SEQ_MODE=4'b1000;
    defparam \ALU.b_15_LC_21_13_4 .LUT_INIT=16'b0011001110100011;
    LogicCell40 \ALU.b_15_LC_21_13_4  (
            .in0(N__53007),
            .in1(N__52932),
            .in2(N__59141),
            .in3(N__67216),
            .lcout(\ALU.bZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73174),
            .ce(N__67931),
            .sr(_gnd_net_));
    defparam \ALU.b_9_LC_21_13_5 .C_ON=1'b0;
    defparam \ALU.b_9_LC_21_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.b_9_LC_21_13_5 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \ALU.b_9_LC_21_13_5  (
            .in0(N__52878),
            .in1(N__66827),
            .in2(N__58565),
            .in3(N__52786),
            .lcout(\ALU.bZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73174),
            .ce(N__67931),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIS1QRR6_0_LC_21_14_0 .C_ON=1'b0;
    defparam \ALU.d_RNIS1QRR6_0_LC_21_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIS1QRR6_0_LC_21_14_0 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \ALU.d_RNIS1QRR6_0_LC_21_14_0  (
            .in0(N__68480),
            .in1(N__48626),
            .in2(N__48719),
            .in3(N__48611),
            .lcout(\ALU.lshift_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_495_c_RNIKOB51J_LC_21_14_1 .C_ON=1'b0;
    defparam \ALU.mult_495_c_RNIKOB51J_LC_21_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_495_c_RNIKOB51J_LC_21_14_1 .LUT_INIT=16'b1100101010101100;
    LogicCell40 \ALU.mult_495_c_RNIKOB51J_LC_21_14_1  (
            .in0(N__57065),
            .in1(N__57134),
            .in2(N__48806),
            .in3(N__48779),
            .lcout(\ALU.mult_495_c_RNIKOB51JZ0 ),
            .ltout(\ALU.mult_495_c_RNIKOB51JZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_8_LC_21_14_2 .C_ON=1'b0;
    defparam \ALU.a_8_LC_21_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.a_8_LC_21_14_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \ALU.a_8_LC_21_14_2  (
            .in0(N__67214),
            .in1(N__51704),
            .in2(N__48755),
            .in3(N__51779),
            .lcout(\ALU.aZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73185),
            .ce(N__71163),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINF0N42_0_LC_21_14_3 .C_ON=1'b0;
    defparam \ALU.d_RNINF0N42_0_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINF0N42_0_LC_21_14_3 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \ALU.d_RNINF0N42_0_LC_21_14_3  (
            .in0(N__66066),
            .in1(N__68479),
            .in2(N__48596),
            .in3(N__68895),
            .lcout(\ALU.lshift_15_ns_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIDDI52_8_LC_21_14_4 .C_ON=1'b0;
    defparam \ALU.d_RNIIDDI52_8_LC_21_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIDDI52_8_LC_21_14_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNIIDDI52_8_LC_21_14_4  (
            .in0(N__48709),
            .in1(N__48673),
            .in2(_gnd_net_),
            .in3(N__66067),
            .lcout(\ALU.N_640 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_7_c_RNIDLTN71_LC_21_14_5 .C_ON=1'b0;
    defparam \ALU.addsub_cry_7_c_RNIDLTN71_LC_21_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_7_c_RNIDLTN71_LC_21_14_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.addsub_cry_7_c_RNIDLTN71_LC_21_14_5  (
            .in0(N__61760),
            .in1(N__67213),
            .in2(_gnd_net_),
            .in3(N__51238),
            .lcout(),
            .ltout(\ALU.addsub_cry_7_c_RNIDLTNZ0Z71_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_7_c_RNIHPLU38_LC_21_14_6 .C_ON=1'b0;
    defparam \ALU.addsub_cry_7_c_RNIHPLU38_LC_21_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_7_c_RNIHPLU38_LC_21_14_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \ALU.addsub_cry_7_c_RNIHPLU38_LC_21_14_6  (
            .in0(N__70159),
            .in1(N__67215),
            .in2(N__48620),
            .in3(N__48617),
            .lcout(\ALU.addsub_cry_7_c_RNIHPLUZ0Z38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO3LAS3_0_LC_21_14_7 .C_ON=1'b0;
    defparam \ALU.d_RNIO3LAS3_0_LC_21_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO3LAS3_0_LC_21_14_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ALU.d_RNIO3LAS3_0_LC_21_14_7  (
            .in0(N__66065),
            .in1(N__48610),
            .in2(N__48595),
            .in3(N__68894),
            .lcout(\ALU.N_809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_1_LC_21_15_0 .C_ON=1'b0;
    defparam \ALU.f_1_LC_21_15_0 .SEQ_MODE=4'b1000;
    defparam \ALU.f_1_LC_21_15_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.f_1_LC_21_15_0  (
            .in0(N__59249),
            .in1(N__52241),
            .in2(N__69698),
            .in3(N__69010),
            .lcout(f_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73192),
            .ce(N__67860),
            .sr(_gnd_net_));
    defparam \ALU.f_0_LC_21_15_1 .C_ON=1'b0;
    defparam \ALU.f_0_LC_21_15_1 .SEQ_MODE=4'b1000;
    defparam \ALU.f_0_LC_21_15_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.f_0_LC_21_15_1  (
            .in0(N__69117),
            .in1(N__52096),
            .in2(N__69699),
            .in3(N__52051),
            .lcout(f_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73192),
            .ce(N__67860),
            .sr(_gnd_net_));
    defparam \ALU.f_7_LC_21_15_2 .C_ON=1'b0;
    defparam \ALU.f_7_LC_21_15_2 .SEQ_MODE=4'b1000;
    defparam \ALU.f_7_LC_21_15_2 .LUT_INIT=16'b0101110101011000;
    LogicCell40 \ALU.f_7_LC_21_15_2  (
            .in0(N__58884),
            .in1(N__51929),
            .in2(N__67286),
            .in3(N__51857),
            .lcout(f_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73192),
            .ce(N__67860),
            .sr(_gnd_net_));
    defparam \ALU.f_8_LC_21_15_3 .C_ON=1'b0;
    defparam \ALU.f_8_LC_21_15_3 .SEQ_MODE=4'b1000;
    defparam \ALU.f_8_LC_21_15_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \ALU.f_8_LC_21_15_3  (
            .in0(N__67269),
            .in1(N__51777),
            .in2(N__51721),
            .in3(N__51634),
            .lcout(f_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73192),
            .ce(N__67860),
            .sr(_gnd_net_));
    defparam \ALU.f_15_LC_21_15_4 .C_ON=1'b0;
    defparam \ALU.f_15_LC_21_15_4 .SEQ_MODE=4'b1000;
    defparam \ALU.f_15_LC_21_15_4 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.f_15_LC_21_15_4  (
            .in0(N__67282),
            .in1(N__52936),
            .in2(N__59143),
            .in3(N__53010),
            .lcout(f_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73192),
            .ce(N__67860),
            .sr(_gnd_net_));
    defparam \ALU.f_9_LC_21_15_5 .C_ON=1'b0;
    defparam \ALU.f_9_LC_21_15_5 .SEQ_MODE=4'b1000;
    defparam \ALU.f_9_LC_21_15_5 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \ALU.f_9_LC_21_15_5  (
            .in0(N__52856),
            .in1(N__66831),
            .in2(N__58563),
            .in3(N__52801),
            .lcout(f_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73192),
            .ce(N__67860),
            .sr(_gnd_net_));
    defparam \ALU.g_1_LC_21_16_0 .C_ON=1'b0;
    defparam \ALU.g_1_LC_21_16_0 .SEQ_MODE=4'b1000;
    defparam \ALU.g_1_LC_21_16_0 .LUT_INIT=16'b0111010101000101;
    LogicCell40 \ALU.g_1_LC_21_16_0  (
            .in0(N__52240),
            .in1(N__59291),
            .in2(N__69746),
            .in3(N__69011),
            .lcout(g_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73199),
            .ce(N__70986),
            .sr(_gnd_net_));
    defparam \ALU.g_0_LC_21_16_1 .C_ON=1'b0;
    defparam \ALU.g_0_LC_21_16_1 .SEQ_MODE=4'b1000;
    defparam \ALU.g_0_LC_21_16_1 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \ALU.g_0_LC_21_16_1  (
            .in0(N__52117),
            .in1(N__69106),
            .in2(N__69745),
            .in3(N__52052),
            .lcout(g_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73199),
            .ce(N__70986),
            .sr(_gnd_net_));
    defparam \ALU.g_7_LC_21_16_2 .C_ON=1'b0;
    defparam \ALU.g_7_LC_21_16_2 .SEQ_MODE=4'b1000;
    defparam \ALU.g_7_LC_21_16_2 .LUT_INIT=16'b0101110101011000;
    LogicCell40 \ALU.g_7_LC_21_16_2  (
            .in0(N__58885),
            .in1(N__51937),
            .in2(N__67267),
            .in3(N__51852),
            .lcout(g_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73199),
            .ce(N__70986),
            .sr(_gnd_net_));
    defparam \ALU.g_8_LC_21_16_3 .C_ON=1'b0;
    defparam \ALU.g_8_LC_21_16_3 .SEQ_MODE=4'b1000;
    defparam \ALU.g_8_LC_21_16_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \ALU.g_8_LC_21_16_3  (
            .in0(N__51703),
            .in1(N__51783),
            .in2(N__67268),
            .in3(N__51636),
            .lcout(g_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73199),
            .ce(N__70986),
            .sr(_gnd_net_));
    defparam \ALU.g_15_LC_21_16_4 .C_ON=1'b0;
    defparam \ALU.g_15_LC_21_16_4 .SEQ_MODE=4'b1000;
    defparam \ALU.g_15_LC_21_16_4 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.g_15_LC_21_16_4  (
            .in0(N__67232),
            .in1(N__52937),
            .in2(N__59120),
            .in3(N__53011),
            .lcout(g_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73199),
            .ce(N__70986),
            .sr(_gnd_net_));
    defparam \ALU.g_9_LC_21_16_5 .C_ON=1'b0;
    defparam \ALU.g_9_LC_21_16_5 .SEQ_MODE=4'b1000;
    defparam \ALU.g_9_LC_21_16_5 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \ALU.g_9_LC_21_16_5  (
            .in0(N__52866),
            .in1(N__66832),
            .in2(N__58551),
            .in3(N__52806),
            .lcout(g_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73199),
            .ce(N__70986),
            .sr(_gnd_net_));
    defparam \ALU.c_RNID85GQ_0_15_LC_21_17_0 .C_ON=1'b0;
    defparam \ALU.c_RNID85GQ_0_15_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNID85GQ_0_15_LC_21_17_0 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \ALU.c_RNID85GQ_0_15_LC_21_17_0  (
            .in0(N__59267),
            .in1(N__49194),
            .in2(N__50543),
            .in3(N__50513),
            .lcout(),
            .ltout(\ALU.c_RNID85GQ_0Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI9DCRE2_15_LC_21_17_1 .C_ON=1'b0;
    defparam \ALU.c_RNI9DCRE2_15_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI9DCRE2_15_LC_21_17_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.c_RNI9DCRE2_15_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(N__74524),
            .in2(N__50354),
            .in3(N__50504),
            .lcout(\ALU.c_RNI9DCRE2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNI117N5_1_LC_21_17_2 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNI117N5_1_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNI117N5_1_LC_21_17_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \CONTROL.busState_1_RNI117N5_1_LC_21_17_2  (
            .in0(N__63592),
            .in1(N__50326),
            .in2(N__50243),
            .in3(N__50215),
            .lcout(N_208),
            .ltout(N_208_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIH202E_15_LC_21_17_3 .C_ON=1'b0;
    defparam \ALU.c_RNIH202E_15_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIH202E_15_LC_21_17_3 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \ALU.c_RNIH202E_15_LC_21_17_3  (
            .in0(N__53757),
            .in1(N__53299),
            .in2(N__49844),
            .in3(N__49592),
            .lcout(\ALU.status_19_14 ),
            .ltout(\ALU.status_19_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJI6SH_15_LC_21_17_4 .C_ON=1'b0;
    defparam \ALU.c_RNIJI6SH_15_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJI6SH_15_LC_21_17_4 .LUT_INIT=16'b0101101010100000;
    LogicCell40 \ALU.c_RNIJI6SH_15_LC_21_17_4  (
            .in0(N__63594),
            .in1(_gnd_net_),
            .in2(N__49841),
            .in3(N__74833),
            .lcout(\ALU.c_RNIJI6SHZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_RNIRLED8_0_LC_21_17_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_RNIRLED8_0_LC_21_17_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.busState_1_RNIRLED8_0_LC_21_17_5 .LUT_INIT=16'b0000001110001011;
    LogicCell40 \CONTROL.busState_1_RNIRLED8_0_LC_21_17_5  (
            .in0(N__49838),
            .in1(N__49832),
            .in2(N__49628),
            .in3(N__49593),
            .lcout(bus_15),
            .ltout(bus_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNID85GQ_15_LC_21_17_6 .C_ON=1'b0;
    defparam \ALU.c_RNID85GQ_15_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNID85GQ_15_LC_21_17_6 .LUT_INIT=16'b1111111001010100;
    LogicCell40 \ALU.c_RNID85GQ_15_LC_21_17_6  (
            .in0(N__50537),
            .in1(N__59266),
            .in2(N__50516),
            .in3(N__50512),
            .lcout(\ALU.c_RNID85GQZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIU5NNB_15_LC_21_17_7 .C_ON=1'b0;
    defparam \ALU.c_RNIU5NNB_15_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIU5NNB_15_LC_21_17_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \ALU.c_RNIU5NNB_15_LC_21_17_7  (
            .in0(N__53758),
            .in1(N__63593),
            .in2(_gnd_net_),
            .in3(N__53300),
            .lcout(\ALU.un14_log_0_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m248_ns_LC_21_18_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m248_ns_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m248_ns_LC_21_18_0 .LUT_INIT=16'b0011101000001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m248_ns_LC_21_18_0  (
            .in0(N__55221),
            .in1(N__76648),
            .in2(N__50921),
            .in3(N__76471),
            .lcout(),
            .ltout(\PROM.ROMDATA.m248_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m249_LC_21_18_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m249_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m249_LC_21_18_1 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m249_LC_21_18_1  (
            .in0(N__76472),
            .in1(N__79873),
            .in2(N__50498),
            .in3(N__50591),
            .lcout(\PROM.ROMDATA.m249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m410_am_LC_21_18_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m410_am_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m410_am_LC_21_18_2 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m410_am_LC_21_18_2  (
            .in0(N__77956),
            .in1(N__78818),
            .in2(N__75814),
            .in3(N__77273),
            .lcout(\PROM.ROMDATA.m410_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m359_LC_21_18_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m359_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m359_LC_21_18_3 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m359_LC_21_18_3  (
            .in0(N__77272),
            .in1(_gnd_net_),
            .in2(N__78860),
            .in3(N__77955),
            .lcout(\PROM.ROMDATA.m359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m304_LC_21_18_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m304_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m304_LC_21_18_5 .LUT_INIT=16'b0001101000001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m304_LC_21_18_5  (
            .in0(N__77274),
            .in1(N__75534),
            .in2(N__78861),
            .in3(N__77957),
            .lcout(\PROM.ROMDATA.m304 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m71_LC_21_18_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m71_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m71_LC_21_18_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m71_LC_21_18_6  (
            .in0(N__77954),
            .in1(N__78814),
            .in2(_gnd_net_),
            .in3(N__77271),
            .lcout(\PROM.ROMDATA.N_72_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m413_bm_LC_21_18_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m413_bm_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m413_bm_LC_21_18_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m413_bm_LC_21_18_7  (
            .in0(N__78819),
            .in1(N__75533),
            .in2(_gnd_net_),
            .in3(N__78984),
            .lcout(\PROM.ROMDATA.m413_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m150_LC_21_19_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m150_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m150_LC_21_19_0 .LUT_INIT=16'b0101101011111010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m150_LC_21_19_0  (
            .in0(N__77142),
            .in1(_gnd_net_),
            .in2(N__78038),
            .in3(N__78810),
            .lcout(\PROM.ROMDATA.m150 ),
            .ltout(\PROM.ROMDATA.m150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m195_am_LC_21_19_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m195_am_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m195_am_LC_21_19_1 .LUT_INIT=16'b0011001100000101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m195_am_LC_21_19_1  (
            .in0(N__75529),
            .in1(N__50693),
            .in2(N__50651),
            .in3(N__76480),
            .lcout(\PROM.ROMDATA.m195_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m228_am_LC_21_19_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m228_am_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m228_am_LC_21_19_2 .LUT_INIT=16'b1010001100001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m228_am_LC_21_19_2  (
            .in0(N__77143),
            .in1(N__75528),
            .in2(N__78040),
            .in3(N__78812),
            .lcout(),
            .ltout(\PROM.ROMDATA.m228_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m229_1_LC_21_19_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m229_1_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m229_1_LC_21_19_3 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m229_1_LC_21_19_3  (
            .in0(N__50590),
            .in1(_gnd_net_),
            .in2(N__50648),
            .in3(N__76481),
            .lcout(\PROM.ROMDATA.m229_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m25_LC_21_19_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m25_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m25_LC_21_19_4 .LUT_INIT=16'b0000011100001001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m25_LC_21_19_4  (
            .in0(N__77140),
            .in1(N__75526),
            .in2(N__78037),
            .in3(N__78809),
            .lcout(\PROM.ROMDATA.m25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m438_LC_21_19_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m438_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m438_LC_21_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m438_LC_21_19_5  (
            .in0(N__54863),
            .in1(N__50633),
            .in2(_gnd_net_),
            .in3(N__79843),
            .lcout(\PROM.ROMDATA.m438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m173_LC_21_19_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m173_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m173_LC_21_19_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m173_LC_21_19_6  (
            .in0(N__77141),
            .in1(N__75527),
            .in2(N__78039),
            .in3(N__78811),
            .lcout(\PROM.ROMDATA.m173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m246_LC_21_19_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m246_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m246_LC_21_19_7 .LUT_INIT=16'b0110011011011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m246_LC_21_19_7  (
            .in0(N__78813),
            .in1(N__77953),
            .in2(_gnd_net_),
            .in3(N__77144),
            .lcout(\PROM.ROMDATA.m246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__g1_LC_21_20_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__g1_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__g1_LC_21_20_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__g1_LC_21_20_0  (
            .in0(N__75659),
            .in1(N__73503),
            .in2(_gnd_net_),
            .in3(N__50579),
            .lcout(PROM_ROMDATA_dintern_31_0__g1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m145_LC_21_20_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m145_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m145_LC_21_20_1 .LUT_INIT=16'b0010111010001001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m145_LC_21_20_1  (
            .in0(N__77805),
            .in1(N__75653),
            .in2(N__78543),
            .in3(N__77123),
            .lcout(\PROM.ROMDATA.m145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m169_LC_21_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m169_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m169_LC_21_20_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m169_LC_21_20_2  (
            .in0(N__77125),
            .in1(N__78320),
            .in2(N__75890),
            .in3(N__77808),
            .lcout(),
            .ltout(\PROM.ROMDATA.m169_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m270_am_LC_21_20_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m270_am_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m270_am_LC_21_20_3 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m270_am_LC_21_20_3  (
            .in0(N__76485),
            .in1(N__79862),
            .in2(N__50723),
            .in3(N__50678),
            .lcout(\PROM.ROMDATA.m270_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m13_LC_21_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m13_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m13_LC_21_20_4 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m13_LC_21_20_4  (
            .in0(N__77124),
            .in1(N__78319),
            .in2(_gnd_net_),
            .in3(N__77806),
            .lcout(\PROM.ROMDATA.m13 ),
            .ltout(\PROM.ROMDATA.m13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m18_am_LC_21_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m18_am_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m18_am_LC_21_20_5 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m18_am_LC_21_20_5  (
            .in0(N__77807),
            .in1(N__75654),
            .in2(N__50696),
            .in3(N__78362),
            .lcout(\PROM.ROMDATA.m18_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m188_LC_21_20_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m188_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m188_LC_21_20_6 .LUT_INIT=16'b0111111101001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m188_LC_21_20_6  (
            .in0(N__77122),
            .in1(N__78315),
            .in2(N__75889),
            .in3(N__77804),
            .lcout(\PROM.ROMDATA.m188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m263_LC_21_20_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m263_LC_21_20_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m263_LC_21_20_7 .LUT_INIT=16'b0110001001000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m263_LC_21_20_7  (
            .in0(N__76484),
            .in1(N__75655),
            .in2(N__50687),
            .in3(N__64964),
            .lcout(\PROM.ROMDATA.m263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_RNIAK8J_1_LC_21_21_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_RNIAK8J_1_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_19_RNIAK8J_1_LC_21_21_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_19_RNIAK8J_1_LC_21_21_0  (
            .in0(N__54901),
            .in1(N__73766),
            .in2(_gnd_net_),
            .in3(N__55122),
            .lcout(\CONTROL.programCounter_ret_19_RNIAK8JZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_1_LC_21_21_1 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_1_LC_21_21_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_1_LC_21_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_1_LC_21_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50672),
            .lcout(\CONTROL.dout_reto_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73248),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_RNI8I8J_0_LC_21_21_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_RNI8I8J_0_LC_21_21_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_19_RNI8I8J_0_LC_21_21_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \CONTROL.programCounter_ret_19_RNI8I8J_0_LC_21_21_2  (
            .in0(N__50986),
            .in1(N__55121),
            .in2(_gnd_net_),
            .in3(N__50948),
            .lcout(\CONTROL.programCounter_ret_19_RNI8I8JZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m74_LC_21_21_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m74_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m74_LC_21_21_3 .LUT_INIT=16'b0100000001111001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m74_LC_21_21_3  (
            .in0(N__77611),
            .in1(N__76966),
            .in2(N__75611),
            .in3(N__78468),
            .lcout(\PROM.ROMDATA.m74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m248_ns_1_LC_21_21_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m248_ns_1_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m248_ns_1_LC_21_21_4 .LUT_INIT=16'b0011011100111101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m248_ns_1_LC_21_21_4  (
            .in0(N__78472),
            .in1(N__75287),
            .in2(N__76454),
            .in3(N__77612),
            .lcout(\PROM.ROMDATA.m248_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_fast_LC_21_21_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_fast_LC_21_21_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_18_fast_LC_21_21_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \CONTROL.programCounter_ret_18_fast_LC_21_21_5  (
            .in0(N__50899),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50835),
            .lcout(\CONTROL.un1_programCounter9_reto_fast ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73248),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m104_ns_1_LC_21_21_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m104_ns_1_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m104_ns_1_LC_21_21_6 .LUT_INIT=16'b0001100000011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m104_ns_1_LC_21_21_6  (
            .in0(N__76965),
            .in1(N__75283),
            .in2(N__78704),
            .in3(_gnd_net_),
            .lcout(\PROM.ROMDATA.m104_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m284_1_LC_21_21_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m284_1_LC_21_21_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m284_1_LC_21_21_7 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m284_1_LC_21_21_7  (
            .in0(N__78569),
            .in1(N__79747),
            .in2(N__75612),
            .in3(N__76268),
            .lcout(\PROM.ROMDATA.m284_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_fast_RNITMBH1_LC_21_22_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_fast_RNITMBH1_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_18_fast_RNITMBH1_LC_21_22_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.programCounter_ret_18_fast_RNITMBH1_LC_21_22_0  (
            .in0(N__55053),
            .in1(N__50747),
            .in2(_gnd_net_),
            .in3(N__50741),
            .lcout(progRomAddress_0),
            .ltout(progRomAddress_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m143_LC_21_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m143_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m143_LC_21_22_1 .LUT_INIT=16'b0100001111010010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m143_LC_21_22_1  (
            .in0(N__77688),
            .in1(N__75236),
            .in2(N__50735),
            .in3(N__78327),
            .lcout(\PROM.ROMDATA.m143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m72_LC_21_22_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m72_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m72_LC_21_22_2 .LUT_INIT=16'b0111111011111001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m72_LC_21_22_2  (
            .in0(N__78328),
            .in1(N__77689),
            .in2(N__75538),
            .in3(N__76927),
            .lcout(),
            .ltout(\PROM.ROMDATA.m72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m80_am_LC_21_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m80_am_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m80_am_LC_21_22_3 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m80_am_LC_21_22_3  (
            .in0(_gnd_net_),
            .in1(N__76273),
            .in2(N__50732),
            .in3(N__50729),
            .lcout(),
            .ltout(\PROM.ROMDATA.m80_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m93_ns_1_LC_21_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m93_ns_1_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m93_ns_1_LC_21_22_4 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m93_ns_1_LC_21_22_4  (
            .in0(N__79314),
            .in1(N__79839),
            .in2(N__51050),
            .in3(N__64757),
            .lcout(\PROM.ROMDATA.m93_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m179_LC_21_22_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m179_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m179_LC_21_22_5 .LUT_INIT=16'b0100000000111001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m179_LC_21_22_5  (
            .in0(N__76925),
            .in1(N__75234),
            .in2(N__77893),
            .in3(N__78325),
            .lcout(\PROM.ROMDATA.m179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_fast_RNI5VBH1_LC_21_22_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_fast_RNI5VBH1_LC_21_22_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_18_fast_RNI5VBH1_LC_21_22_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \CONTROL.programCounter_ret_18_fast_RNI5VBH1_LC_21_22_6  (
            .in0(N__55054),
            .in1(N__51035),
            .in2(_gnd_net_),
            .in3(N__51029),
            .lcout(progRomAddress_2),
            .ltout(progRomAddress_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m127_LC_21_22_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m127_LC_21_22_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m127_LC_21_22_7 .LUT_INIT=16'b0000111101011011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m127_LC_21_22_7  (
            .in0(N__76926),
            .in1(N__75235),
            .in2(N__51023),
            .in3(N__78326),
            .lcout(\PROM.ROMDATA.m127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m196_ns_1_LC_21_23_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m196_ns_1_LC_21_23_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m196_ns_1_LC_21_23_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m196_ns_1_LC_21_23_0  (
            .in0(N__79844),
            .in1(N__55253),
            .in2(N__79413),
            .in3(N__50996),
            .lcout(),
            .ltout(\PROM.ROMDATA.m196_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m196_ns_LC_21_23_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m196_ns_LC_21_23_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m196_ns_LC_21_23_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m196_ns_LC_21_23_1  (
            .in0(N__51164),
            .in1(N__51020),
            .in2(N__51008),
            .in3(N__79318),
            .lcout(\PROM.ROMDATA.m196_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m185_am_LC_21_23_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m185_am_LC_21_23_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m185_am_LC_21_23_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m185_am_LC_21_23_2  (
            .in0(N__51005),
            .in1(N__76269),
            .in2(_gnd_net_),
            .in3(N__74185),
            .lcout(\PROM.ROMDATA.m185_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m193_LC_21_23_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m193_LC_21_23_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m193_LC_21_23_3 .LUT_INIT=16'b0010100000000001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m193_LC_21_23_3  (
            .in0(N__77608),
            .in1(N__76977),
            .in2(N__75886),
            .in3(N__78677),
            .lcout(\PROM.ROMDATA.m193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m191_LC_21_23_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m191_LC_21_23_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m191_LC_21_23_4 .LUT_INIT=16'b0110111011111010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m191_LC_21_23_4  (
            .in0(N__76978),
            .in1(N__78679),
            .in2(N__75960),
            .in3(N__77609),
            .lcout(),
            .ltout(\PROM.ROMDATA.m191_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m195_bm_LC_21_23_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m195_bm_LC_21_23_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m195_bm_LC_21_23_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m195_bm_LC_21_23_5  (
            .in0(N__76270),
            .in1(_gnd_net_),
            .in2(N__51173),
            .in3(N__51170),
            .lcout(\PROM.ROMDATA.m195_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_3_LC_21_23_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_3_LC_21_23_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_3_LC_21_23_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \CONTROL.programCounter_ret_1_3_LC_21_23_6  (
            .in0(_gnd_net_),
            .in1(N__51158),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.programCounter_1_reto_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73267),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m92_am_LC_21_23_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m92_am_LC_21_23_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m92_am_LC_21_23_7 .LUT_INIT=16'b1100000110100001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m92_am_LC_21_23_7  (
            .in0(N__77610),
            .in1(N__75821),
            .in2(N__55205),
            .in3(N__78678),
            .lcout(\PROM.ROMDATA.m92_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m62_LC_21_24_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m62_LC_21_24_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m62_LC_21_24_0 .LUT_INIT=16'b0100001011011100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m62_LC_21_24_0  (
            .in0(N__77794),
            .in1(N__78694),
            .in2(N__75903),
            .in3(N__77151),
            .lcout(),
            .ltout(\PROM.ROMDATA.m62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m64_bm_LC_21_24_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m64_bm_LC_21_24_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m64_bm_LC_21_24_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m64_bm_LC_21_24_1  (
            .in0(N__54922),
            .in1(_gnd_net_),
            .in2(N__51098),
            .in3(N__76322),
            .lcout(\PROM.ROMDATA.m64_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m65_ns_1_LC_21_24_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m65_ns_1_LC_21_24_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m65_ns_1_LC_21_24_2 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m65_ns_1_LC_21_24_2  (
            .in0(N__79319),
            .in1(N__51095),
            .in2(N__51086),
            .in3(N__79840),
            .lcout(),
            .ltout(\PROM.ROMDATA.m65_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m65_ns_LC_21_24_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m65_ns_LC_21_24_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m65_ns_LC_21_24_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m65_ns_LC_21_24_3  (
            .in0(N__51074),
            .in1(N__51374),
            .in2(N__51068),
            .in3(N__79320),
            .lcout(m65_ns),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_RNIGQ8J_4_LC_21_24_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_RNIGQ8J_4_LC_21_24_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_19_RNIGQ8J_4_LC_21_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_19_RNIGQ8J_4_LC_21_24_4  (
            .in0(N__55294),
            .in1(N__55155),
            .in2(_gnd_net_),
            .in3(N__55138),
            .lcout(\CONTROL.programCounter_ret_19_RNIGQ8JZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m58_LC_21_24_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m58_LC_21_24_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m58_LC_21_24_5 .LUT_INIT=16'b0001001001101101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m58_LC_21_24_5  (
            .in0(N__77150),
            .in1(N__78686),
            .in2(N__75962),
            .in3(N__77795),
            .lcout(),
            .ltout(\PROM.ROMDATA.m58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m64_am_LC_21_24_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m64_am_LC_21_24_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m64_am_LC_21_24_6 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m64_am_LC_21_24_6  (
            .in0(N__76321),
            .in1(_gnd_net_),
            .in2(N__51377),
            .in3(N__55196),
            .lcout(\PROM.ROMDATA.m64_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m45_LC_21_24_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m45_LC_21_24_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m45_LC_21_24_7 .LUT_INIT=16'b0101001101110001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m45_LC_21_24_7  (
            .in0(N__77149),
            .in1(N__78685),
            .in2(N__75961),
            .in3(N__77793),
            .lcout(\PROM.ROMDATA.m45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNID1RPI_14_LC_22_9_0 .C_ON=1'b0;
    defparam \ALU.c_RNID1RPI_14_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNID1RPI_14_LC_22_9_0 .LUT_INIT=16'b0011011011101000;
    LogicCell40 \ALU.c_RNID1RPI_14_LC_22_9_0  (
            .in0(N__63116),
            .in1(N__74860),
            .in2(N__63848),
            .in3(N__56741),
            .lcout(\ALU.log_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_20_0_LC_22_9_1 .C_ON=1'b0;
    defparam \ALU.status_RNO_20_0_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_20_0_LC_22_9_1 .LUT_INIT=16'b0001111011101000;
    LogicCell40 \ALU.status_RNO_20_0_LC_22_9_1  (
            .in0(N__63114),
            .in1(N__66314),
            .in2(N__74886),
            .in3(N__68943),
            .lcout(\ALU.status_8_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_14_0_LC_22_9_2 .C_ON=1'b0;
    defparam \ALU.status_RNO_14_0_LC_22_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_14_0_LC_22_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALU.status_RNO_14_0_LC_22_9_2  (
            .in0(N__51359),
            .in1(N__51344),
            .in2(N__51323),
            .in3(N__51295),
            .lcout(),
            .ltout(\ALU.status_8_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_7_0_LC_22_9_3 .C_ON=1'b0;
    defparam \ALU.status_RNO_7_0_LC_22_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_7_0_LC_22_9_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ALU.status_RNO_7_0_LC_22_9_3  (
            .in0(N__51263),
            .in1(N__51242),
            .in2(N__51206),
            .in3(N__51179),
            .lcout(\ALU.status_8_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_19_0_LC_22_9_5 .C_ON=1'b0;
    defparam \ALU.status_RNO_19_0_LC_22_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_19_0_LC_22_9_5 .LUT_INIT=16'b0100101110110010;
    LogicCell40 \ALU.status_RNO_19_0_LC_22_9_5  (
            .in0(N__63115),
            .in1(N__53048),
            .in2(N__74887),
            .in3(N__74607),
            .lcout(),
            .ltout(\ALU.log_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_15_0_LC_22_9_6 .C_ON=1'b0;
    defparam \ALU.status_RNO_15_0_LC_22_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_15_0_LC_22_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALU.status_RNO_15_0_LC_22_9_6  (
            .in0(N__57248),
            .in1(N__51188),
            .in2(N__51182),
            .in3(N__57514),
            .lcout(\ALU.status_8_13_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIV5AOK_13_LC_22_10_0 .C_ON=1'b0;
    defparam \ALU.c_RNIV5AOK_13_LC_22_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIV5AOK_13_LC_22_10_0 .LUT_INIT=16'b0001111011101000;
    LogicCell40 \ALU.c_RNIV5AOK_13_LC_22_10_0  (
            .in0(N__63301),
            .in1(N__61009),
            .in2(N__74826),
            .in3(N__56829),
            .lcout(\ALU.c_RNIV5AOKZ0Z_13 ),
            .ltout(\ALU.c_RNIV5AOKZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIO5N04A_0_13_LC_22_10_1 .C_ON=1'b0;
    defparam \ALU.c_RNIO5N04A_0_13_LC_22_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIO5N04A_0_13_LC_22_10_1 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \ALU.c_RNIO5N04A_0_13_LC_22_10_1  (
            .in0(N__70198),
            .in1(N__58533),
            .in2(N__51554),
            .in3(N__51502),
            .lcout(\ALU.c_RNIO5N04A_0Z0Z_13 ),
            .ltout(\ALU.c_RNIO5N04A_0Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_13_LC_22_10_2 .C_ON=1'b0;
    defparam \ALU.b_13_LC_22_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.b_13_LC_22_10_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.b_13_LC_22_10_2  (
            .in0(_gnd_net_),
            .in1(N__67432),
            .in2(N__51551),
            .in3(N__67388),
            .lcout(\ALU.bZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73158),
            .ce(N__67942),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIO5N04A_13_LC_22_10_3 .C_ON=1'b0;
    defparam \ALU.c_RNIO5N04A_13_LC_22_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIO5N04A_13_LC_22_10_3 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \ALU.c_RNIO5N04A_13_LC_22_10_3  (
            .in0(N__70199),
            .in1(N__51515),
            .in2(N__51509),
            .in3(N__58534),
            .lcout(\ALU.c_RNIO5N04AZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_13_0_LC_22_10_4 .C_ON=1'b0;
    defparam \ALU.status_RNO_13_0_LC_22_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_13_0_LC_22_10_4 .LUT_INIT=16'b0001111011101000;
    LogicCell40 \ALU.status_RNO_13_0_LC_22_10_4  (
            .in0(N__63299),
            .in1(N__61008),
            .in2(N__74825),
            .in3(N__56828),
            .lcout(),
            .ltout(\ALU.N_16_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_6_0_LC_22_10_5 .C_ON=1'b0;
    defparam \ALU.status_RNO_6_0_LC_22_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_6_0_LC_22_10_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \ALU.status_RNO_6_0_LC_22_10_5  (
            .in0(N__51490),
            .in1(_gnd_net_),
            .in2(N__51461),
            .in3(N__51443),
            .lcout(\ALU.status_8_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_12_0_LC_22_10_6 .C_ON=1'b0;
    defparam \ALU.status_RNO_12_0_LC_22_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_12_0_LC_22_10_6 .LUT_INIT=16'b1100101110010010;
    LogicCell40 \ALU.status_RNO_12_0_LC_22_10_6  (
            .in0(N__63298),
            .in1(N__62939),
            .in2(N__74824),
            .in3(N__62887),
            .lcout(\ALU.log_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7KS2I_9_LC_22_10_7 .C_ON=1'b0;
    defparam \ALU.d_RNI7KS2I_9_LC_22_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7KS2I_9_LC_22_10_7 .LUT_INIT=16'b1110001110000110;
    LogicCell40 \ALU.d_RNI7KS2I_9_LC_22_10_7  (
            .in0(N__62888),
            .in1(N__74771),
            .in2(N__62949),
            .in3(N__63300),
            .lcout(\ALU.d_RNI7KS2IZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_12_LC_22_11_0 .C_ON=1'b0;
    defparam \ALU.e_12_LC_22_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.e_12_LC_22_11_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \ALU.e_12_LC_22_11_0  (
            .in0(_gnd_net_),
            .in1(N__67743),
            .in2(N__67602),
            .in3(N__67655),
            .lcout(\ALU.eZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73164),
            .ce(N__69245),
            .sr(_gnd_net_));
    defparam \ALU.e_13_LC_22_11_1 .C_ON=1'b0;
    defparam \ALU.e_13_LC_22_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.e_13_LC_22_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.e_13_LC_22_11_1  (
            .in0(N__67494),
            .in1(N__67442),
            .in2(_gnd_net_),
            .in3(N__67392),
            .lcout(\ALU.eZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73164),
            .ce(N__69245),
            .sr(_gnd_net_));
    defparam \ALU.e_14_LC_22_11_2 .C_ON=1'b0;
    defparam \ALU.e_14_LC_22_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.e_14_LC_22_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_14_LC_22_11_2  (
            .in0(N__68137),
            .in1(N__68057),
            .in2(_gnd_net_),
            .in3(N__68004),
            .lcout(\ALU.eZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73164),
            .ce(N__69245),
            .sr(_gnd_net_));
    defparam \ALU.g_12_LC_22_12_0 .C_ON=1'b0;
    defparam \ALU.g_12_LC_22_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.g_12_LC_22_12_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.g_12_LC_22_12_0  (
            .in0(N__67741),
            .in1(N__67668),
            .in2(_gnd_net_),
            .in3(N__67595),
            .lcout(g_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73175),
            .ce(N__70993),
            .sr(_gnd_net_));
    defparam \ALU.g_13_LC_22_12_1 .C_ON=1'b0;
    defparam \ALU.g_13_LC_22_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.g_13_LC_22_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.g_13_LC_22_12_1  (
            .in0(N__67455),
            .in1(N__67512),
            .in2(_gnd_net_),
            .in3(N__67400),
            .lcout(g_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73175),
            .ce(N__70993),
            .sr(_gnd_net_));
    defparam \ALU.g_14_LC_22_12_2 .C_ON=1'b0;
    defparam \ALU.g_14_LC_22_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.g_14_LC_22_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_14_LC_22_12_2  (
            .in0(N__68138),
            .in1(N__68086),
            .in2(_gnd_net_),
            .in3(N__68001),
            .lcout(g_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73175),
            .ce(N__70993),
            .sr(_gnd_net_));
    defparam \ALU.d_1_LC_22_13_0 .C_ON=1'b0;
    defparam \ALU.d_1_LC_22_13_0 .SEQ_MODE=4'b1000;
    defparam \ALU.d_1_LC_22_13_0 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.d_1_LC_22_13_0  (
            .in0(N__59305),
            .in1(N__69690),
            .in2(N__52247),
            .in3(N__68989),
            .lcout(\ALU.dZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73186),
            .ce(N__70250),
            .sr(_gnd_net_));
    defparam \ALU.d_0_LC_22_13_1 .C_ON=1'b0;
    defparam \ALU.d_0_LC_22_13_1 .SEQ_MODE=4'b1000;
    defparam \ALU.d_0_LC_22_13_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ALU.d_0_LC_22_13_1  (
            .in0(N__69156),
            .in1(N__52124),
            .in2(N__69715),
            .in3(N__52053),
            .lcout(\ALU.dZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73186),
            .ce(N__70250),
            .sr(_gnd_net_));
    defparam \ALU.d_7_LC_22_13_2 .C_ON=1'b0;
    defparam \ALU.d_7_LC_22_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.d_7_LC_22_13_2 .LUT_INIT=16'b0111010101100100;
    LogicCell40 \ALU.d_7_LC_22_13_2  (
            .in0(N__58864),
            .in1(N__67254),
            .in2(N__51938),
            .in3(N__51862),
            .lcout(\ALU.dZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73186),
            .ce(N__70250),
            .sr(_gnd_net_));
    defparam \ALU.d_8_LC_22_13_3 .C_ON=1'b0;
    defparam \ALU.d_8_LC_22_13_3 .SEQ_MODE=4'b1000;
    defparam \ALU.d_8_LC_22_13_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \ALU.d_8_LC_22_13_3  (
            .in0(N__67252),
            .in1(N__51778),
            .in2(N__51722),
            .in3(N__51635),
            .lcout(\ALU.dZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73186),
            .ce(N__70250),
            .sr(_gnd_net_));
    defparam \ALU.d_15_LC_22_13_4 .C_ON=1'b0;
    defparam \ALU.d_15_LC_22_13_4 .SEQ_MODE=4'b1000;
    defparam \ALU.d_15_LC_22_13_4 .LUT_INIT=16'b0010000011101111;
    LogicCell40 \ALU.d_15_LC_22_13_4  (
            .in0(N__53008),
            .in1(N__67253),
            .in2(N__59142),
            .in3(N__52935),
            .lcout(\ALU.dZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73186),
            .ce(N__70250),
            .sr(_gnd_net_));
    defparam \ALU.d_9_LC_22_13_5 .C_ON=1'b0;
    defparam \ALU.d_9_LC_22_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.d_9_LC_22_13_5 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \ALU.d_9_LC_22_13_5  (
            .in0(N__52870),
            .in1(N__66806),
            .in2(N__58564),
            .in3(N__52788),
            .lcout(\ALU.dZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73186),
            .ce(N__70250),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPFFDD1_0_6_LC_22_14_0 .C_ON=1'b0;
    defparam \ALU.d_RNIPFFDD1_0_6_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPFFDD1_0_6_LC_22_14_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ALU.d_RNIPFFDD1_0_6_LC_22_14_0  (
            .in0(N__66766),
            .in1(N__62583),
            .in2(N__59645),
            .in3(N__66074),
            .lcout(),
            .ltout(\ALU.d_RNIPFFDD1_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBTSVI3_6_LC_22_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNIBTSVI3_6_LC_22_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBTSVI3_6_LC_22_14_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNIBTSVI3_6_LC_22_14_1  (
            .in0(N__52709),
            .in1(_gnd_net_),
            .in2(N__52691),
            .in3(N__52493),
            .lcout(\ALU.N_863 ),
            .ltout(\ALU.N_863_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGPBNB6_2_LC_22_14_2 .C_ON=1'b0;
    defparam \ALU.d_RNIGPBNB6_2_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGPBNB6_2_LC_22_14_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNIGPBNB6_2_LC_22_14_2  (
            .in0(N__68935),
            .in1(_gnd_net_),
            .in2(N__52688),
            .in3(N__68174),
            .lcout(),
            .ltout(\ALU.d_RNIGPBNB6Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIUDSOL9_2_LC_22_14_3 .C_ON=1'b0;
    defparam \ALU.d_RNIUDSOL9_2_LC_22_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIUDSOL9_2_LC_22_14_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIUDSOL9_2_LC_22_14_3  (
            .in0(_gnd_net_),
            .in1(N__52683),
            .in2(N__52640),
            .in3(N__52499),
            .lcout(\ALU.a_15_m0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINGV0T2_15_LC_22_14_4 .C_ON=1'b0;
    defparam \ALU.c_RNINGV0T2_15_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINGV0T2_15_LC_22_14_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ALU.c_RNINGV0T2_15_LC_22_14_4  (
            .in0(N__68934),
            .in1(N__69973),
            .in2(N__68556),
            .in3(N__52527),
            .lcout(\ALU.c_RNINGV0T2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPFFDD1_6_LC_22_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNIPFFDD1_6_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPFFDD1_6_LC_22_14_5 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \ALU.d_RNIPFFDD1_6_LC_22_14_5  (
            .in0(N__66073),
            .in1(N__59640),
            .in2(N__62588),
            .in3(N__66765),
            .lcout(\ALU.d_RNIPFFDD1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_16_0_LC_22_14_6 .C_ON=1'b0;
    defparam \ALU.status_RNO_16_0_LC_22_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_16_0_LC_22_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ALU.status_RNO_16_0_LC_22_14_6  (
            .in0(_gnd_net_),
            .in1(N__60358),
            .in2(_gnd_net_),
            .in3(N__60319),
            .lcout(),
            .ltout(\ALU.status_14_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_8_0_LC_22_14_7 .C_ON=1'b0;
    defparam \ALU.status_RNO_8_0_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_8_0_LC_22_14_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ALU.status_RNO_8_0_LC_22_14_7  (
            .in0(N__60280),
            .in1(N__59929),
            .in2(N__53363),
            .in3(N__61753),
            .lcout(\ALU.status_14_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_10_0_LC_22_15_0 .C_ON=1'b0;
    defparam \ALU.status_RNO_10_0_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_10_0_LC_22_15_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ALU.status_RNO_10_0_LC_22_15_0  (
            .in0(N__62338),
            .in1(N__62047),
            .in2(_gnd_net_),
            .in3(N__61492),
            .lcout(),
            .ltout(\ALU.status_14_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_4_0_LC_22_15_1 .C_ON=1'b0;
    defparam \ALU.status_RNO_4_0_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_4_0_LC_22_15_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.status_RNO_4_0_LC_22_15_1  (
            .in0(N__53036),
            .in1(N__63699),
            .in2(N__53345),
            .in3(N__63512),
            .lcout(\ALU.status_14_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIHLMGP_14_LC_22_15_2 .C_ON=1'b0;
    defparam \ALU.c_RNIHLMGP_14_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIHLMGP_14_LC_22_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.c_RNIHLMGP_14_LC_22_15_2  (
            .in0(N__61014),
            .in1(N__63774),
            .in2(_gnd_net_),
            .in3(N__66736),
            .lcout(\ALU.N_979 ),
            .ltout(\ALU.N_979_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIUMNP22_15_LC_22_15_3 .C_ON=1'b0;
    defparam \ALU.c_RNIUMNP22_15_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIUMNP22_15_LC_22_15_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ALU.c_RNIUMNP22_15_LC_22_15_3  (
            .in0(N__63639),
            .in1(N__66742),
            .in2(N__53309),
            .in3(N__66076),
            .lcout(\ALU.N_968 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_22_0_LC_22_15_4 .C_ON=1'b0;
    defparam \ALU.status_RNO_22_0_LC_22_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_22_0_LC_22_15_4 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \ALU.status_RNO_22_0_LC_22_15_4  (
            .in0(N__53762),
            .in1(N__63638),
            .in2(N__63274),
            .in3(N__53177),
            .lcout(\ALU.status_RNO_22Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_9_0_LC_22_15_5 .C_ON=1'b0;
    defparam \ALU.status_RNO_9_0_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_9_0_LC_22_15_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ALU.status_RNO_9_0_LC_22_15_5  (
            .in0(N__59665),
            .in1(N__59353),
            .in2(_gnd_net_),
            .in3(N__66856),
            .lcout(\ALU.status_14_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIVHVMK_13_LC_22_15_6 .C_ON=1'b0;
    defparam \ALU.c_RNIVHVMK_13_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIVHVMK_13_LC_22_15_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \ALU.c_RNIVHVMK_13_LC_22_15_6  (
            .in0(N__63225),
            .in1(N__61018),
            .in2(N__56839),
            .in3(_gnd_net_),
            .lcout(\ALU.c_RNIVHVMKZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_17_I_21_c_RNO_LC_22_16_0 .C_ON=1'b0;
    defparam \ALU.status_17_I_21_c_RNO_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_17_I_21_c_RNO_LC_22_16_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \ALU.status_17_I_21_c_RNO_LC_22_16_0  (
            .in0(N__56719),
            .in1(N__63778),
            .in2(N__63613),
            .in3(N__74570),
            .lcout(\ALU.status_17_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIDDGOI_14_LC_22_16_1 .C_ON=1'b0;
    defparam \ALU.c_RNIDDGOI_14_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIDDGOI_14_LC_22_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.c_RNIDDGOI_14_LC_22_16_1  (
            .in0(N__63779),
            .in1(N__63240),
            .in2(_gnd_net_),
            .in3(N__56718),
            .lcout(\ALU.c_RNIDDGOIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_e_0_RNO_0_2_LC_22_16_2 .C_ON=1'b0;
    defparam \ALU.status_e_0_RNO_0_2_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_e_0_RNO_0_2_LC_22_16_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.status_e_0_RNO_0_2_LC_22_16_2  (
            .in0(N__69519),
            .in1(N__53690),
            .in2(_gnd_net_),
            .in3(N__63516),
            .lcout(),
            .ltout(\ALU.status_e_0_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_e_0_2_LC_22_16_3 .C_ON=1'b0;
    defparam \ALU.status_e_0_2_LC_22_16_3 .SEQ_MODE=4'b1000;
    defparam \ALU.status_e_0_2_LC_22_16_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.status_e_0_2_LC_22_16_3  (
            .in0(_gnd_net_),
            .in1(N__56543),
            .in2(N__53732),
            .in3(N__53726),
            .lcout(aluStatus_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73208),
            .ce(N__56603),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI0NMSH_15_LC_22_16_4 .C_ON=1'b0;
    defparam \ALU.c_RNI0NMSH_15_LC_22_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI0NMSH_15_LC_22_16_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.c_RNI0NMSH_15_LC_22_16_4  (
            .in0(N__63241),
            .in1(_gnd_net_),
            .in2(N__63614),
            .in3(N__74569),
            .lcout(\ALU.c_RNI0NMSHZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_e_0_RNO_2_2_LC_22_16_5 .C_ON=1'b0;
    defparam \ALU.status_e_0_RNO_2_2_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_e_0_RNO_2_2_LC_22_16_5 .LUT_INIT=16'b0110011010001000;
    LogicCell40 \ALU.status_e_0_RNO_2_2_LC_22_16_5  (
            .in0(N__74571),
            .in1(N__74856),
            .in2(_gnd_net_),
            .in3(N__63582),
            .lcout(),
            .ltout(\ALU.N_570_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_e_0_RNO_1_2_LC_22_16_6 .C_ON=1'b0;
    defparam \ALU.status_e_0_RNO_1_2_LC_22_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_e_0_RNO_1_2_LC_22_16_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.status_e_0_RNO_1_2_LC_22_16_6  (
            .in0(N__63242),
            .in1(_gnd_net_),
            .in2(N__53729),
            .in3(N__74528),
            .lcout(\ALU.status_e_0_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.g3_0_LC_22_16_7 .C_ON=1'b0;
    defparam \CONTROL.g3_0_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.g3_0_LC_22_16_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \CONTROL.g3_0_LC_22_16_7  (
            .in0(N__53689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53669),
            .lcout(\CONTROL.g3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI9NEO1_15_LC_22_17_0 .C_ON=1'b0;
    defparam \ALU.b_RNI9NEO1_15_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI9NEO1_15_LC_22_17_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.b_RNI9NEO1_15_LC_22_17_0  (
            .in0(N__53611),
            .in1(N__53588),
            .in2(N__53517),
            .in3(N__53478),
            .lcout(),
            .ltout(\ALU.operand2_6_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKIDM2_15_LC_22_17_1 .C_ON=1'b0;
    defparam \ALU.d_RNIKIDM2_15_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKIDM2_15_LC_22_17_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIKIDM2_15_LC_22_17_1  (
            .in0(N__54186),
            .in1(N__54328),
            .in2(N__53438),
            .in3(N__53434),
            .lcout(\ALU.N_1260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIILK02_15_LC_22_17_2 .C_ON=1'b0;
    defparam \ALU.d_RNIILK02_15_LC_22_17_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIILK02_15_LC_22_17_2 .LUT_INIT=16'b1011001110000011;
    LogicCell40 \ALU.d_RNIILK02_15_LC_22_17_2  (
            .in0(N__54329),
            .in1(N__54317),
            .in2(N__54308),
            .in3(N__54187),
            .lcout(),
            .ltout(\ALU.N_1148_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI2SRO3_15_LC_22_17_3 .C_ON=1'b0;
    defparam \ALU.c_RNI2SRO3_15_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI2SRO3_15_LC_22_17_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.c_RNI2SRO3_15_LC_22_17_3  (
            .in0(_gnd_net_),
            .in1(N__54161),
            .in2(N__54146),
            .in3(N__54140),
            .lcout(aluOut_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI8VV95_15_LC_22_17_4 .C_ON=1'b0;
    defparam \ALU.c_RNI8VV95_15_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI8VV95_15_LC_22_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNI8VV95_15_LC_22_17_4  (
            .in0(N__53990),
            .in1(N__53984),
            .in2(_gnd_net_),
            .in3(N__53968),
            .lcout(),
            .ltout(\ALU.c_RNI8VV95Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJTKD7_15_LC_22_17_5 .C_ON=1'b0;
    defparam \ALU.c_RNIJTKD7_15_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJTKD7_15_LC_22_17_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.c_RNIJTKD7_15_LC_22_17_5  (
            .in0(_gnd_net_),
            .in1(N__53783),
            .in2(N__53765),
            .in3(N__71463),
            .lcout(\ALU.c_RNIJTKD7Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m320_bm_LC_22_18_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m320_bm_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m320_bm_LC_22_18_0 .LUT_INIT=16'b0100100010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m320_bm_LC_22_18_0  (
            .in0(N__78776),
            .in1(N__77993),
            .in2(N__75965),
            .in3(N__77304),
            .lcout(),
            .ltout(\PROM.ROMDATA.m320_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m320_ns_LC_22_18_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m320_ns_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m320_ns_LC_22_18_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m320_ns_LC_22_18_1  (
            .in0(_gnd_net_),
            .in1(N__54401),
            .in2(N__53744),
            .in3(N__76475),
            .lcout(\PROM.ROMDATA.m320_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m413_am_LC_22_18_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m413_am_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m413_am_LC_22_18_2 .LUT_INIT=16'b0000000001000011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m413_am_LC_22_18_2  (
            .in0(N__78774),
            .in1(N__77989),
            .in2(N__75964),
            .in3(N__77302),
            .lcout(),
            .ltout(\PROM.ROMDATA.m413_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m414_ns_1_LC_22_18_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m414_ns_1_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m414_ns_1_LC_22_18_3 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m414_ns_1_LC_22_18_3  (
            .in0(N__79874),
            .in1(N__53741),
            .in2(N__53735),
            .in3(N__76474),
            .lcout(\PROM.ROMDATA.m414_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_2_LC_22_18_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_2_LC_22_18_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_2_LC_22_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.programCounter_ret_19_2_LC_22_18_4  (
            .in0(N__54821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\CONTROL.dout_reto_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73226),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.un1_busState97_i_i_LC_22_18_5 .C_ON=1'b0;
    defparam \CONTROL.un1_busState97_i_i_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.un1_busState97_i_i_LC_22_18_5 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \CONTROL.un1_busState97_i_i_LC_22_18_5  (
            .in0(N__54782),
            .in1(N__54770),
            .in2(N__54752),
            .in3(N__54685),
            .lcout(\CONTROL.N_45_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m139_LC_22_18_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m139_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m139_LC_22_18_6 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m139_LC_22_18_6  (
            .in0(N__78773),
            .in1(N__77988),
            .in2(_gnd_net_),
            .in3(N__77301),
            .lcout(\PROM.ROMDATA.m139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m320_am_LC_22_18_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m320_am_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m320_am_LC_22_18_7 .LUT_INIT=16'b0001111000110010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m320_am_LC_22_18_7  (
            .in0(N__77303),
            .in1(N__75839),
            .in2(N__78054),
            .in3(N__78775),
            .lcout(\PROM.ROMDATA.m320_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m154_LC_22_19_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m154_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m154_LC_22_19_1 .LUT_INIT=16'b1000110100000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m154_LC_22_19_1  (
            .in0(N__75831),
            .in1(N__54395),
            .in2(N__64286),
            .in3(N__74061),
            .lcout(\PROM.ROMDATA.N_558_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m323_bm_LC_22_19_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m323_bm_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m323_bm_LC_22_19_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m323_bm_LC_22_19_2  (
            .in0(N__78736),
            .in1(N__75832),
            .in2(N__79048),
            .in3(N__77982),
            .lcout(\PROM.ROMDATA.m323_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m49_LC_22_19_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m49_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m49_LC_22_19_3 .LUT_INIT=16'b0000101010101111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m49_LC_22_19_3  (
            .in0(N__77165),
            .in1(_gnd_net_),
            .in2(N__78049),
            .in3(N__78735),
            .lcout(),
            .ltout(\PROM.ROMDATA.m49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m228_bm_LC_22_19_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m228_bm_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m228_bm_LC_22_19_4 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m228_bm_LC_22_19_4  (
            .in0(_gnd_net_),
            .in1(N__55222),
            .in2(N__54374),
            .in3(N__75830),
            .lcout(),
            .ltout(\PROM.ROMDATA.m228_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m229_LC_22_19_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m229_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m229_LC_22_19_5 .LUT_INIT=16'b1011000100100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m229_LC_22_19_5  (
            .in0(N__79842),
            .in1(N__54371),
            .in2(N__54365),
            .in3(N__76473),
            .lcout(\PROM.ROMDATA.m229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m226_LC_22_19_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m226_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m226_LC_22_19_6 .LUT_INIT=16'b0110011000100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m226_LC_22_19_6  (
            .in0(N__78734),
            .in1(N__77977),
            .in2(_gnd_net_),
            .in3(N__77164),
            .lcout(\PROM.ROMDATA.m226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m312_bm_LC_22_19_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m312_bm_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m312_bm_LC_22_19_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m312_bm_LC_22_19_7  (
            .in0(N__77981),
            .in1(N__73905),
            .in2(N__75963),
            .in3(N__78737),
            .lcout(\PROM.ROMDATA.m312_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m437_ns_LC_22_20_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m437_ns_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m437_ns_LC_22_20_0 .LUT_INIT=16'b0010001011010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m437_ns_LC_22_20_0  (
            .in0(N__54836),
            .in1(N__76460),
            .in2(N__64442),
            .in3(N__77121),
            .lcout(\PROM.ROMDATA.m437_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m11_bm_LC_22_20_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m11_bm_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m11_bm_LC_22_20_1 .LUT_INIT=16'b0100010101111001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m11_bm_LC_22_20_1  (
            .in0(N__77118),
            .in1(N__75645),
            .in2(N__77973),
            .in3(N__78330),
            .lcout(\PROM.ROMDATA.m11_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m118_LC_22_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m118_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m118_LC_22_20_2 .LUT_INIT=16'b0110101100011110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m118_LC_22_20_2  (
            .in0(N__78329),
            .in1(N__77796),
            .in2(N__75887),
            .in3(N__77117),
            .lcout(\PROM.ROMDATA.m118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m312_ns_LC_22_20_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m312_ns_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m312_ns_LC_22_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m312_ns_LC_22_20_3  (
            .in0(N__76461),
            .in1(N__54857),
            .in2(_gnd_net_),
            .in3(N__54851),
            .lcout(\PROM.ROMDATA.m312_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m437_ns_1_LC_22_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m437_ns_1_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m437_ns_1_LC_22_20_4 .LUT_INIT=16'b0000100001111101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m437_ns_1_LC_22_20_4  (
            .in0(N__78332),
            .in1(N__77803),
            .in2(N__75888),
            .in3(N__77120),
            .lcout(\PROM.ROMDATA.m437_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m18_bm_LC_22_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m18_bm_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m18_bm_LC_22_20_5 .LUT_INIT=16'b0000001011100001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m18_bm_LC_22_20_5  (
            .in0(N__77119),
            .in1(N__75646),
            .in2(N__77974),
            .in3(N__78331),
            .lcout(),
            .ltout(\PROM.ROMDATA.m18_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m19_ns_1_LC_22_20_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m19_ns_1_LC_22_20_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m19_ns_1_LC_22_20_6 .LUT_INIT=16'b0001110100110011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m19_ns_1_LC_22_20_6  (
            .in0(N__54830),
            .in1(N__79841),
            .in2(N__54824),
            .in3(N__76458),
            .lcout(),
            .ltout(\PROM.ROMDATA.m19_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m19_ns_LC_22_20_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m19_ns_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m19_ns_LC_22_20_7 .LUT_INIT=16'b0100111101001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m19_ns_LC_22_20_7  (
            .in0(N__76459),
            .in1(N__54956),
            .in2(N__54944),
            .in3(N__54941),
            .lcout(\PROM.ROMDATA.m19_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m111_LC_22_21_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m111_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m111_LC_22_21_0 .LUT_INIT=16'b0101001101011010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m111_LC_22_21_0  (
            .in0(N__76911),
            .in1(N__78323),
            .in2(N__77838),
            .in3(N__75423),
            .lcout(\PROM.ROMDATA.m111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m117_LC_22_21_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m117_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m117_LC_22_21_1 .LUT_INIT=16'b0110001111001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m117_LC_22_21_1  (
            .in0(N__78321),
            .in1(N__77575),
            .in2(N__75709),
            .in3(N__76909),
            .lcout(\PROM.ROMDATA.m117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m33_LC_22_21_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m33_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m33_LC_22_21_2 .LUT_INIT=16'b0011001000110110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m33_LC_22_21_2  (
            .in0(N__76913),
            .in1(N__78324),
            .in2(N__77839),
            .in3(N__75424),
            .lcout(\PROM.ROMDATA.m33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m211_ns_N_2L1_LC_22_21_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m211_ns_N_2L1_LC_22_21_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m211_ns_N_2L1_LC_22_21_3 .LUT_INIT=16'b0011100100011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m211_ns_N_2L1_LC_22_21_3  (
            .in0(N__78322),
            .in1(N__76173),
            .in2(N__75710),
            .in3(N__76910),
            .lcout(\PROM.ROMDATA.m211_ns_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIJA5J_1_LC_22_21_4 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIJA5J_1_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIJA5J_1_LC_22_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIJA5J_1_LC_22_21_4  (
            .in0(N__55064),
            .in1(N__54902),
            .in2(_gnd_net_),
            .in3(N__54890),
            .lcout(N_416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNIH68I_1_LC_22_21_5 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNIH68I_1_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNIH68I_1_LC_22_21_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNIH68I_1_LC_22_21_5  (
            .in0(N__54889),
            .in1(N__73787),
            .in2(_gnd_net_),
            .in3(N__55139),
            .lcout(),
            .ltout(\CONTROL.programCounter_ret_1_RNIH68IZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_fast_RNI1RBH1_LC_22_21_6 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_fast_RNI1RBH1_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_18_fast_RNI1RBH1_LC_22_21_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \CONTROL.programCounter_ret_18_fast_RNI1RBH1_LC_22_21_6  (
            .in0(_gnd_net_),
            .in1(N__55055),
            .in2(N__54875),
            .in3(N__54872),
            .lcout(progRomAddress_1),
            .ltout(progRomAddress_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m114_LC_22_21_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m114_LC_22_21_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m114_LC_22_21_7 .LUT_INIT=16'b0100100111010101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m114_LC_22_21_7  (
            .in0(N__75422),
            .in1(N__77576),
            .in2(N__54866),
            .in3(N__76912),
            .lcout(\PROM.ROMDATA.m114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m492_am_LC_22_22_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m492_am_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m492_am_LC_22_22_0 .LUT_INIT=16'b0011010100000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m492_am_LC_22_22_0  (
            .in0(N__73542),
            .in1(N__73811),
            .in2(N__73741),
            .in3(N__77700),
            .lcout(\PROM.ROMDATA.m492_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m55_LC_22_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m55_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m55_LC_22_22_1 .LUT_INIT=16'b0101111000010010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m55_LC_22_22_1  (
            .in0(N__77073),
            .in1(N__75817),
            .in2(N__77895),
            .in3(N__78339),
            .lcout(\PROM.ROMDATA.m55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_RNINC8I_4_LC_22_22_2 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_RNINC8I_4_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_1_RNINC8I_4_LC_22_22_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \CONTROL.programCounter_ret_1_RNINC8I_4_LC_22_22_2  (
            .in0(N__55184),
            .in1(N__55169),
            .in2(_gnd_net_),
            .in3(N__55137),
            .lcout(),
            .ltout(\CONTROL.programCounter_ret_1_RNINC8IZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_18_fast_RNID7CH1_LC_22_22_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_18_fast_RNID7CH1_LC_22_22_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.programCounter_ret_18_fast_RNID7CH1_LC_22_22_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \CONTROL.programCounter_ret_18_fast_RNID7CH1_LC_22_22_3  (
            .in0(_gnd_net_),
            .in1(N__55058),
            .in2(N__55013),
            .in3(N__55010),
            .lcout(progRomAddress_4),
            .ltout(progRomAddress_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m147_bm_LC_22_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m147_bm_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m147_bm_LC_22_22_4 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m147_bm_LC_22_22_4  (
            .in0(_gnd_net_),
            .in1(N__54998),
            .in2(N__54992),
            .in3(N__54989),
            .lcout(\PROM.ROMDATA.m147_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m140_LC_22_22_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m140_LC_22_22_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m140_LC_22_22_5 .LUT_INIT=16'b0111000111101001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m140_LC_22_22_5  (
            .in0(N__77072),
            .in1(N__75816),
            .in2(N__77894),
            .in3(N__78338),
            .lcout(\PROM.ROMDATA.m140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m156_LC_22_22_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m156_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m156_LC_22_22_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m156_LC_22_22_6  (
            .in0(N__78337),
            .in1(N__77693),
            .in2(_gnd_net_),
            .in3(N__77071),
            .lcout(\PROM.ROMDATA.m156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m92_bm_LC_22_22_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m92_bm_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m92_bm_LC_22_22_7 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m92_bm_LC_22_22_7  (
            .in0(N__54980),
            .in1(N__65183),
            .in2(_gnd_net_),
            .in3(N__76286),
            .lcout(\PROM.ROMDATA.m92_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m183_LC_22_23_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m183_LC_22_23_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m183_LC_22_23_0 .LUT_INIT=16'b0011011010011100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m183_LC_22_23_0  (
            .in0(N__64642),
            .in1(N__76264),
            .in2(N__64531),
            .in3(N__64485),
            .lcout(\PROM.ROMDATA.m183 ),
            .ltout(\PROM.ROMDATA.m183_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m185_bm_LC_22_23_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m185_bm_LC_22_23_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m185_bm_LC_22_23_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m185_bm_LC_22_23_1  (
            .in0(_gnd_net_),
            .in1(N__55244),
            .in2(N__55256),
            .in3(N__64919),
            .lcout(\PROM.ROMDATA.m185_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m166_LC_22_23_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m166_LC_22_23_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m166_LC_22_23_2 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m166_LC_22_23_2  (
            .in0(N__76930),
            .in1(N__78790),
            .in2(N__77841),
            .in3(N__75631),
            .lcout(\PROM.ROMDATA.N_525_mux ),
            .ltout(\PROM.ROMDATA.N_525_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m427_bm_LC_22_23_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m427_bm_LC_22_23_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m427_bm_LC_22_23_3 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m427_bm_LC_22_23_3  (
            .in0(N__75635),
            .in1(N__64017),
            .in2(N__55247),
            .in3(N__76287),
            .lcout(\PROM.ROMDATA.m427_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m164_LC_22_23_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m164_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m164_LC_22_23_4 .LUT_INIT=16'b0100000000000001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m164_LC_22_23_4  (
            .in0(N__76929),
            .in1(N__78789),
            .in2(N__77840),
            .in3(N__75630),
            .lcout(\PROM.ROMDATA.m164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m132_LC_22_23_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m132_LC_22_23_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m132_LC_22_23_5 .LUT_INIT=16'b0010010000101111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m132_LC_22_23_5  (
            .in0(N__78791),
            .in1(N__77590),
            .in2(N__75885),
            .in3(N__76931),
            .lcout(\PROM.ROMDATA.m132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m492_bm_LC_22_23_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m492_bm_LC_22_23_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m492_bm_LC_22_23_6 .LUT_INIT=16'b0000000100110001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m492_bm_LC_22_23_6  (
            .in0(N__73553),
            .in1(N__64862),
            .in2(N__73742),
            .in3(N__73810),
            .lcout(\PROM.ROMDATA.m492_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m133_LC_22_23_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m133_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m133_LC_22_23_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m133_LC_22_23_7  (
            .in0(N__78788),
            .in1(N__77583),
            .in2(_gnd_net_),
            .in3(N__76928),
            .lcout(\PROM.ROMDATA.m133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m182_LC_22_24_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m182_LC_22_24_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m182_LC_22_24_0 .LUT_INIT=16'b0000000001000010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m182_LC_22_24_0  (
            .in0(N__77145),
            .in1(N__76291),
            .in2(N__77975),
            .in3(N__78795),
            .lcout(\PROM.ROMDATA.i4_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m338_bm_LC_22_24_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m338_bm_LC_22_24_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m338_bm_LC_22_24_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m338_bm_LC_22_24_1  (
            .in0(N__55238),
            .in1(N__75828),
            .in2(_gnd_net_),
            .in3(N__55226),
            .lcout(\PROM.ROMDATA.m338_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m92_am_1_LC_22_24_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m92_am_1_LC_22_24_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m92_am_1_LC_22_24_2 .LUT_INIT=16'b0011011101110010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m92_am_1_LC_22_24_2  (
            .in0(N__77147),
            .in1(N__76292),
            .in2(N__77976),
            .in3(N__75688),
            .lcout(\PROM.ROMDATA.m92_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m158_LC_22_24_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m158_LC_22_24_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m158_LC_22_24_3 .LUT_INIT=16'b0000000010000100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m158_LC_22_24_3  (
            .in0(N__78797),
            .in1(N__77816),
            .in2(N__75902),
            .in3(N__77148),
            .lcout(\PROM.ROMDATA.m158 ),
            .ltout(\PROM.ROMDATA.m158_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m162_LC_22_24_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m162_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m162_LC_22_24_4 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m162_LC_22_24_4  (
            .in0(N__79838),
            .in1(N__76293),
            .in2(N__55484),
            .in3(N__64925),
            .lcout(\PROM.ROMDATA.m162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m135_LC_22_24_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m135_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m135_LC_22_24_5 .LUT_INIT=16'b0101010010010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m135_LC_22_24_5  (
            .in0(N__78796),
            .in1(N__77812),
            .in2(N__75901),
            .in3(N__77146),
            .lcout(\PROM.ROMDATA.m135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m202_LC_22_24_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m202_LC_22_24_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m202_LC_22_24_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m202_LC_22_24_6  (
            .in0(N__74065),
            .in1(N__72731),
            .in2(N__64142),
            .in3(N__55481),
            .lcout(PROM_ROMDATA_dintern_6ro),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m317_am_LC_22_24_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m317_am_LC_22_24_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m317_am_LC_22_24_7 .LUT_INIT=16'b1101100101100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m317_am_LC_22_24_7  (
            .in0(N__78798),
            .in1(N__75829),
            .in2(N__73891),
            .in3(N__78989),
            .lcout(\PROM.ROMDATA.m317_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_19_4_LC_22_25_0 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_19_4_LC_22_25_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_19_4_LC_22_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_19_4_LC_22_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55333),
            .lcout(\CONTROL.dout_reto_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73279),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_0_c_inv_LC_23_7_0 .C_ON=1'b1;
    defparam \ALU.status_19_cry_0_c_inv_LC_23_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_0_c_inv_LC_23_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_0_c_inv_LC_23_7_0  (
            .in0(_gnd_net_),
            .in1(N__66772),
            .in2(N__55283),
            .in3(N__60579),
            .lcout(\ALU.aluOut_i_0 ),
            .ltout(),
            .carryin(bfn_23_7_0_),
            .carryout(\ALU.status_19_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_1_c_inv_LC_23_7_1 .C_ON=1'b1;
    defparam \ALU.status_19_cry_1_c_inv_LC_23_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_1_c_inv_LC_23_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_1_c_inv_LC_23_7_1  (
            .in0(_gnd_net_),
            .in1(N__66084),
            .in2(N__55274),
            .in3(N__65537),
            .lcout(\ALU.aluOut_i_1 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_0 ),
            .carryout(\ALU.status_19_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_2_c_inv_LC_23_7_2 .C_ON=1'b1;
    defparam \ALU.status_19_cry_2_c_inv_LC_23_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_2_c_inv_LC_23_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_2_c_inv_LC_23_7_2  (
            .in0(_gnd_net_),
            .in1(N__68945),
            .in2(N__55265),
            .in3(N__66320),
            .lcout(\ALU.aluOut_i_2 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_1 ),
            .carryout(\ALU.status_19_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_3_c_inv_LC_23_7_3 .C_ON=1'b1;
    defparam \ALU.status_19_cry_3_c_inv_LC_23_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_3_c_inv_LC_23_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_3_c_inv_LC_23_7_3  (
            .in0(_gnd_net_),
            .in1(N__68525),
            .in2(N__56426),
            .in3(N__60266),
            .lcout(\ALU.aluOut_i_3 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_2 ),
            .carryout(\ALU.status_19_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_4_c_inv_LC_23_7_4 .C_ON=1'b1;
    defparam \ALU.status_19_cry_4_c_inv_LC_23_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_4_c_inv_LC_23_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_4_c_inv_LC_23_7_4  (
            .in0(_gnd_net_),
            .in1(N__56417),
            .in2(N__56285),
            .in3(N__59883),
            .lcout(\ALU.aluOut_i_4 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_3 ),
            .carryout(\ALU.status_19_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_5_c_inv_LC_23_7_5 .C_ON=1'b1;
    defparam \ALU.status_19_cry_5_c_inv_LC_23_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_5_c_inv_LC_23_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_5_c_inv_LC_23_7_5  (
            .in0(_gnd_net_),
            .in1(N__56276),
            .in2(N__56150),
            .in3(N__59644),
            .lcout(\ALU.aluOut_i_5 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_4 ),
            .carryout(\ALU.status_19_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_6_c_inv_LC_23_7_6 .C_ON=1'b1;
    defparam \ALU.status_19_cry_6_c_inv_LC_23_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_6_c_inv_LC_23_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_6_c_inv_LC_23_7_6  (
            .in0(_gnd_net_),
            .in1(N__56131),
            .in2(N__56003),
            .in3(N__62550),
            .lcout(\ALU.aluOut_i_6 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_5 ),
            .carryout(\ALU.status_19_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_7_c_inv_LC_23_7_7 .C_ON=1'b1;
    defparam \ALU.status_19_cry_7_c_inv_LC_23_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_7_c_inv_LC_23_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_7_c_inv_LC_23_7_7  (
            .in0(_gnd_net_),
            .in1(N__55991),
            .in2(N__55835),
            .in3(N__62298),
            .lcout(\ALU.aluOut_i_7 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_6 ),
            .carryout(\ALU.status_19_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_8_c_inv_LC_23_8_0 .C_ON=1'b1;
    defparam \ALU.status_19_cry_8_c_inv_LC_23_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_8_c_inv_LC_23_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_8_c_inv_LC_23_8_0  (
            .in0(_gnd_net_),
            .in1(N__55822),
            .in2(N__55697),
            .in3(N__62024),
            .lcout(\ALU.aluOut_i_8 ),
            .ltout(),
            .carryin(bfn_23_8_0_),
            .carryout(\ALU.status_19_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_9_c_inv_LC_23_8_1 .C_ON=1'b1;
    defparam \ALU.status_19_cry_9_c_inv_LC_23_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_9_c_inv_LC_23_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_9_c_inv_LC_23_8_1  (
            .in0(_gnd_net_),
            .in1(N__55687),
            .in2(N__55598),
            .in3(N__62889),
            .lcout(\ALU.aluOut_i_9 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_8 ),
            .carryout(\ALU.status_19_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_10_c_inv_LC_23_8_2 .C_ON=1'b1;
    defparam \ALU.status_19_cry_10_c_inv_LC_23_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_10_c_inv_LC_23_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_10_c_inv_LC_23_8_2  (
            .in0(_gnd_net_),
            .in1(N__55589),
            .in2(N__55517),
            .in3(N__61701),
            .lcout(\ALU.aluOut_i_10 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_9 ),
            .carryout(\ALU.status_19_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_11_c_inv_LC_23_8_3 .C_ON=1'b1;
    defparam \ALU.status_19_cry_11_c_inv_LC_23_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_11_c_inv_LC_23_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.status_19_cry_11_c_inv_LC_23_8_3  (
            .in0(N__61475),
            .in1(N__57053),
            .in2(N__56942),
            .in3(_gnd_net_),
            .lcout(\ALU.aluOut_i_11 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_10 ),
            .carryout(\ALU.status_19_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_12_c_inv_LC_23_8_4 .C_ON=1'b1;
    defparam \ALU.status_19_cry_12_c_inv_LC_23_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_12_c_inv_LC_23_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_12_c_inv_LC_23_8_4  (
            .in0(_gnd_net_),
            .in1(N__56933),
            .in2(N__56852),
            .in3(N__61226),
            .lcout(\ALU.aluOut_i_12 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_11 ),
            .carryout(\ALU.status_19_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_13_c_inv_LC_23_8_5 .C_ON=1'b1;
    defparam \ALU.status_19_cry_13_c_inv_LC_23_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_13_c_inv_LC_23_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_13_c_inv_LC_23_8_5  (
            .in0(_gnd_net_),
            .in1(N__56759),
            .in2(N__56843),
            .in3(N__61011),
            .lcout(\ALU.aluOut_i_13 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_12 ),
            .carryout(\ALU.status_19_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_14_c_inv_LC_23_8_6 .C_ON=1'b1;
    defparam \ALU.status_19_cry_14_c_inv_LC_23_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_14_c_inv_LC_23_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.status_19_cry_14_c_inv_LC_23_8_6  (
            .in0(_gnd_net_),
            .in1(N__56749),
            .in2(N__56678),
            .in3(N__63852),
            .lcout(\ALU.aluOut_i_14 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_13 ),
            .carryout(\ALU.status_19_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_19_cry_15_c_inv_LC_23_8_7 .C_ON=1'b1;
    defparam \ALU.status_19_cry_15_c_inv_LC_23_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.status_19_cry_15_c_inv_LC_23_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ALU.status_19_cry_15_c_inv_LC_23_8_7  (
            .in0(N__63640),
            .in1(N__74603),
            .in2(N__56669),
            .in3(_gnd_net_),
            .lcout(\ALU.aluOut_i_15 ),
            .ltout(),
            .carryin(\ALU.status_19_cry_14 ),
            .carryout(\ALU.status_19Z0Z_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_5_LC_23_9_0 .C_ON=1'b0;
    defparam \ALU.status_5_LC_23_9_0 .SEQ_MODE=4'b1000;
    defparam \ALU.status_5_LC_23_9_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ALU.status_5_LC_23_9_0  (
            .in0(N__69513),
            .in1(N__56622),
            .in2(N__56647),
            .in3(N__56660),
            .lcout(aluStatus_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73159),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_1_LC_23_9_1 .C_ON=1'b0;
    defparam \ALU.status_1_LC_23_9_1 .SEQ_MODE=4'b1000;
    defparam \ALU.status_1_LC_23_9_1 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \ALU.status_1_LC_23_9_1  (
            .in0(N__56621),
            .in1(N__63414),
            .in2(N__56542),
            .in3(N__63389),
            .lcout(aluStatus_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73159),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI12L8C5_2_LC_23_9_3 .C_ON=1'b0;
    defparam \ALU.d_RNI12L8C5_2_LC_23_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI12L8C5_2_LC_23_9_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ALU.d_RNI12L8C5_2_LC_23_9_3  (
            .in0(N__56492),
            .in1(N__68524),
            .in2(N__56472),
            .in3(N__68944),
            .lcout(\ALU.d_RNI12L8C5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_18_0_LC_23_9_5 .C_ON=1'b0;
    defparam \ALU.status_RNO_18_0_LC_23_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_18_0_LC_23_9_5 .LUT_INIT=16'b0001111011101000;
    LogicCell40 \ALU.status_RNO_18_0_LC_23_9_5  (
            .in0(N__63113),
            .in1(N__60265),
            .in2(N__74902),
            .in3(N__68523),
            .lcout(\ALU.log_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_12_c_RNIP50IR3_LC_23_10_1 .C_ON=1'b0;
    defparam \ALU.addsub_cry_12_c_RNIP50IR3_LC_23_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_12_c_RNIP50IR3_LC_23_10_1 .LUT_INIT=16'b0000011111110111;
    LogicCell40 \ALU.addsub_cry_12_c_RNIP50IR3_LC_23_10_1  (
            .in0(N__57242),
            .in1(N__68565),
            .in2(N__67243),
            .in3(N__60835),
            .lcout(),
            .ltout(\ALU.a_15_d_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_558_c_RNIB75F9G_LC_23_10_2 .C_ON=1'b0;
    defparam \ALU.mult_558_c_RNIB75F9G_LC_23_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_558_c_RNIB75F9G_LC_23_10_2 .LUT_INIT=16'b0000111100101110;
    LogicCell40 \ALU.mult_558_c_RNIB75F9G_LC_23_10_2  (
            .in0(N__57185),
            .in1(N__57121),
            .in2(N__57176),
            .in3(N__67183),
            .lcout(\ALU.mult_558_c_RNIB75F9GZ0 ),
            .ltout(\ALU.mult_558_c_RNIB75F9GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_13_LC_23_10_3 .C_ON=1'b0;
    defparam \ALU.a_13_LC_23_10_3 .SEQ_MODE=4'b1000;
    defparam \ALU.a_13_LC_23_10_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ALU.a_13_LC_23_10_3  (
            .in0(N__67493),
            .in1(_gnd_net_),
            .in2(N__57173),
            .in3(N__67450),
            .lcout(\ALU.aZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73165),
            .ce(N__71214),
            .sr(_gnd_net_));
    defparam \ALU.a_15_d_s_10_LC_23_10_4 .C_ON=1'b0;
    defparam \ALU.a_15_d_s_10_LC_23_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_d_s_10_LC_23_10_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.a_15_d_s_10_LC_23_10_4  (
            .in0(N__59136),
            .in1(N__67179),
            .in2(_gnd_net_),
            .in3(N__69908),
            .lcout(\ALU.a_15_d_sZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJ7J1M5_0_2_LC_23_10_5 .C_ON=1'b0;
    defparam \ALU.d_RNIJ7J1M5_0_2_LC_23_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJ7J1M5_0_2_LC_23_10_5 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \ALU.d_RNIJ7J1M5_0_2_LC_23_10_5  (
            .in0(N__59159),
            .in1(N__57109),
            .in2(N__57122),
            .in3(N__57073),
            .lcout(\ALU.d_RNIJ7J1M5_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m3_d_s_8_LC_23_10_6 .C_ON=1'b0;
    defparam \ALU.a_15_m3_d_s_8_LC_23_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m3_d_s_8_LC_23_10_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \ALU.a_15_m3_d_s_8_LC_23_10_6  (
            .in0(N__59137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__69907),
            .lcout(\ALU.a_15_m3_d_sZ0Z_8 ),
            .ltout(\ALU.a_15_m3_d_sZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJ7J1M5_2_LC_23_10_7 .C_ON=1'b0;
    defparam \ALU.d_RNIJ7J1M5_2_LC_23_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJ7J1M5_2_LC_23_10_7 .LUT_INIT=16'b1111101100001011;
    LogicCell40 \ALU.d_RNIJ7J1M5_2_LC_23_10_7  (
            .in0(N__59158),
            .in1(N__57110),
            .in2(N__57077),
            .in3(N__57074),
            .lcout(\ALU.d_RNIJ7J1M5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_12_LC_23_11_0 .C_ON=1'b0;
    defparam \ALU.f_12_LC_23_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.f_12_LC_23_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.f_12_LC_23_11_0  (
            .in0(N__67754),
            .in1(N__67672),
            .in2(_gnd_net_),
            .in3(N__67603),
            .lcout(f_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73176),
            .ce(N__67864),
            .sr(_gnd_net_));
    defparam \ALU.f_13_LC_23_11_1 .C_ON=1'b0;
    defparam \ALU.f_13_LC_23_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.f_13_LC_23_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.f_13_LC_23_11_1  (
            .in0(N__67449),
            .in1(N__67504),
            .in2(_gnd_net_),
            .in3(N__67390),
            .lcout(f_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73176),
            .ce(N__67864),
            .sr(_gnd_net_));
    defparam \ALU.f_14_LC_23_11_2 .C_ON=1'b0;
    defparam \ALU.f_14_LC_23_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.f_14_LC_23_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.f_14_LC_23_11_2  (
            .in0(N__68058),
            .in1(N__68123),
            .in2(_gnd_net_),
            .in3(N__68000),
            .lcout(f_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73176),
            .ce(N__67864),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_13_c_RNIBVHEA1_LC_23_12_0 .C_ON=1'b0;
    defparam \ALU.addsub_cry_13_c_RNIBVHEA1_LC_23_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_13_c_RNIBVHEA1_LC_23_12_0 .LUT_INIT=16'b1010111110100011;
    LogicCell40 \ALU.addsub_cry_13_c_RNIBVHEA1_LC_23_12_0  (
            .in0(N__63701),
            .in1(N__59287),
            .in2(N__67270),
            .in3(N__57523),
            .lcout(\ALU.addsub_cry_13_c_RNIBVHEAZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_13_c_RNIBVHEA1_0_LC_23_12_1 .C_ON=1'b0;
    defparam \ALU.addsub_cry_13_c_RNIBVHEA1_0_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_13_c_RNIBVHEA1_0_LC_23_12_1 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \ALU.addsub_cry_13_c_RNIBVHEA1_0_LC_23_12_1  (
            .in0(N__59288),
            .in1(N__67248),
            .in2(N__57527),
            .in3(N__63700),
            .lcout(),
            .ltout(\ALU.addsub_cry_13_c_RNIBVHEA1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_13_c_RNIJMTGA5_LC_23_12_2 .C_ON=1'b0;
    defparam \ALU.addsub_cry_13_c_RNIJMTGA5_LC_23_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_13_c_RNIJMTGA5_LC_23_12_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.addsub_cry_13_c_RNIJMTGA5_LC_23_12_2  (
            .in0(_gnd_net_),
            .in1(N__57503),
            .in2(N__57488),
            .in3(N__57485),
            .lcout(),
            .ltout(\ALU.addsub_cry_13_c_RNIJMTGAZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_561_c_RNI1EB5TL_LC_23_12_3 .C_ON=1'b0;
    defparam \ALU.mult_561_c_RNI1EB5TL_LC_23_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_561_c_RNI1EB5TL_LC_23_12_3 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \ALU.mult_561_c_RNI1EB5TL_LC_23_12_3  (
            .in0(N__59107),
            .in1(N__67251),
            .in2(N__57479),
            .in3(N__57476),
            .lcout(\ALU.a_15_ns_rn_0_14 ),
            .ltout(\ALU.a_15_ns_rn_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_14_LC_23_12_4 .C_ON=1'b0;
    defparam \ALU.a_14_LC_23_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.a_14_LC_23_12_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.a_14_LC_23_12_4  (
            .in0(_gnd_net_),
            .in1(N__68122),
            .in2(N__57461),
            .in3(N__68087),
            .lcout(\ALU.aZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73187),
            .ce(N__71200),
            .sr(_gnd_net_));
    defparam \ALU.a_15_s_3_LC_23_12_5 .C_ON=1'b0;
    defparam \ALU.a_15_s_3_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_s_3_LC_23_12_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ALU.a_15_s_3_LC_23_12_5  (
            .in0(N__59286),
            .in1(N__59102),
            .in2(_gnd_net_),
            .in3(N__67244),
            .lcout(\ALU.a_15_sZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_ns_sn_14_LC_23_12_6 .C_ON=1'b0;
    defparam \ALU.a_15_ns_sn_14_LC_23_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_ns_sn_14_LC_23_12_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.a_15_ns_sn_14_LC_23_12_6  (
            .in0(N__67249),
            .in1(N__59106),
            .in2(_gnd_net_),
            .in3(N__59339),
            .lcout(\ALU.a_15_ns_snZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_6_c_RNIJ7U2L_LC_23_12_7 .C_ON=1'b0;
    defparam \ALU.addsub_cry_6_c_RNIJ7U2L_LC_23_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_6_c_RNIJ7U2L_LC_23_12_7 .LUT_INIT=16'b0000000111001101;
    LogicCell40 \ALU.addsub_cry_6_c_RNIJ7U2L_LC_23_12_7  (
            .in0(N__59289),
            .in1(N__67250),
            .in2(N__59138),
            .in3(N__62048),
            .lcout(\ALU.a_15_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_3_LC_23_13_0 .C_ON=1'b0;
    defparam \ALU.h_3_LC_23_13_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_3_LC_23_13_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \ALU.h_3_LC_23_13_0  (
            .in0(_gnd_net_),
            .in1(N__58817),
            .in2(N__58756),
            .in3(N__58677),
            .lcout(h_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73193),
            .ce(N__69451),
            .sr(_gnd_net_));
    defparam \ALU.h_10_LC_23_13_1 .C_ON=1'b0;
    defparam \ALU.h_10_LC_23_13_1 .SEQ_MODE=4'b1000;
    defparam \ALU.h_10_LC_23_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.h_10_LC_23_13_1  (
            .in0(N__58562),
            .in1(N__58372),
            .in2(_gnd_net_),
            .in3(N__58301),
            .lcout(h_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73193),
            .ce(N__69451),
            .sr(_gnd_net_));
    defparam \ALU.h_11_LC_23_13_2 .C_ON=1'b0;
    defparam \ALU.h_11_LC_23_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.h_11_LC_23_13_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.h_11_LC_23_13_2  (
            .in0(_gnd_net_),
            .in1(N__58195),
            .in2(N__58127),
            .in3(N__58056),
            .lcout(h_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73193),
            .ce(N__69451),
            .sr(_gnd_net_));
    defparam \ALU.h_12_LC_23_13_3 .C_ON=1'b0;
    defparam \ALU.h_12_LC_23_13_3 .SEQ_MODE=4'b1000;
    defparam \ALU.h_12_LC_23_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.h_12_LC_23_13_3  (
            .in0(N__67755),
            .in1(N__67687),
            .in2(_gnd_net_),
            .in3(N__67617),
            .lcout(h_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73193),
            .ce(N__69451),
            .sr(_gnd_net_));
    defparam \ALU.h_13_LC_23_13_4 .C_ON=1'b0;
    defparam \ALU.h_13_LC_23_13_4 .SEQ_MODE=4'b1000;
    defparam \ALU.h_13_LC_23_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.h_13_LC_23_13_4  (
            .in0(N__67460),
            .in1(N__67517),
            .in2(_gnd_net_),
            .in3(N__67399),
            .lcout(h_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73193),
            .ce(N__69451),
            .sr(_gnd_net_));
    defparam \ALU.h_14_LC_23_13_5 .C_ON=1'b0;
    defparam \ALU.h_14_LC_23_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.h_14_LC_23_13_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.h_14_LC_23_13_5  (
            .in0(N__68078),
            .in1(N__68139),
            .in2(_gnd_net_),
            .in3(N__68002),
            .lcout(h_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73193),
            .ce(N__69451),
            .sr(_gnd_net_));
    defparam \CONTROL.addrstackptr_RNI0D361_4_LC_23_13_6 .C_ON=1'b0;
    defparam \CONTROL.addrstackptr_RNI0D361_4_LC_23_13_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.addrstackptr_RNI0D361_4_LC_23_13_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \CONTROL.addrstackptr_RNI0D361_4_LC_23_13_6  (
            .in0(N__57801),
            .in1(_gnd_net_),
            .in2(N__60818),
            .in3(N__60736),
            .lcout(\CONTROL.g1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_0_c_THRU_CRY_0_LC_23_14_0 .C_ON=1'b1;
    defparam \ALU.addsub_cry_0_c_THRU_CRY_0_LC_23_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_0_c_THRU_CRY_0_LC_23_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.addsub_cry_0_c_THRU_CRY_0_LC_23_14_0  (
            .in0(_gnd_net_),
            .in1(N__63276),
            .in2(N__63297),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_23_14_0_),
            .carryout(\ALU.addsub_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4KF5H_0_LC_23_14_1 .C_ON=1'b1;
    defparam \ALU.d_RNI4KF5H_0_LC_23_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4KF5H_0_LC_23_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.d_RNI4KF5H_0_LC_23_14_1  (
            .in0(_gnd_net_),
            .in1(N__60625),
            .in2(N__60386),
            .in3(N__60347),
            .lcout(\ALU.addsub_0 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_0_c_THRU_CO ),
            .carryout(\ALU.addsub_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_0_c_RNISBATS_LC_23_14_2 .C_ON=1'b1;
    defparam \ALU.addsub_cry_0_c_RNISBATS_LC_23_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_0_c_RNISBATS_LC_23_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_0_c_RNISBATS_LC_23_14_2  (
            .in0(_gnd_net_),
            .in1(N__65536),
            .in2(N__60344),
            .in3(N__60308),
            .lcout(\ALU.addsub_1 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_0 ),
            .carryout(\ALU.addsub_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_1_c_RNIRBVRO_LC_23_14_3 .C_ON=1'b1;
    defparam \ALU.addsub_cry_1_c_RNIRBVRO_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_1_c_RNIRBVRO_LC_23_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_1_c_RNIRBVRO_LC_23_14_3  (
            .in0(_gnd_net_),
            .in1(N__66303),
            .in2(N__60305),
            .in3(N__60269),
            .lcout(\ALU.addsub_2 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_1 ),
            .carryout(\ALU.addsub_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_2_c_RNIDOASJ_LC_23_14_4 .C_ON=1'b1;
    defparam \ALU.addsub_cry_2_c_RNIDOASJ_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_2_c_RNIDOASJ_LC_23_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_2_c_RNIDOASJ_LC_23_14_4  (
            .in0(_gnd_net_),
            .in1(N__60236),
            .in2(N__59957),
            .in3(N__59915),
            .lcout(\ALU.addsub_3 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_2 ),
            .carryout(\ALU.addsub_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_3_c_RNI67KIM_LC_23_14_5 .C_ON=1'b1;
    defparam \ALU.addsub_cry_3_c_RNI67KIM_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_3_c_RNI67KIM_LC_23_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_3_c_RNI67KIM_LC_23_14_5  (
            .in0(_gnd_net_),
            .in1(N__59882),
            .in2(N__59693),
            .in3(N__59648),
            .lcout(\ALU.addsub_4 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_3 ),
            .carryout(\ALU.addsub_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_4_c_RNIDE0RM_LC_23_14_6 .C_ON=1'b1;
    defparam \ALU.addsub_cry_4_c_RNIDE0RM_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_4_c_RNIDE0RM_LC_23_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_4_c_RNIDE0RM_LC_23_14_6  (
            .in0(_gnd_net_),
            .in1(N__59639),
            .in2(N__59384),
            .in3(N__59342),
            .lcout(\ALU.addsub_5 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_4 ),
            .carryout(\ALU.addsub_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_5_c_RNIR5MEM_LC_23_14_7 .C_ON=1'b1;
    defparam \ALU.addsub_cry_5_c_RNIR5MEM_LC_23_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_5_c_RNIR5MEM_LC_23_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_5_c_RNIR5MEM_LC_23_14_7  (
            .in0(_gnd_net_),
            .in1(N__62586),
            .in2(N__62366),
            .in3(N__62327),
            .lcout(\ALU.addsub_6 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_5 ),
            .carryout(\ALU.addsub_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_6_c_RNI112DK_LC_23_15_0 .C_ON=1'b1;
    defparam \ALU.addsub_cry_6_c_RNI112DK_LC_23_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_6_c_RNI112DK_LC_23_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_6_c_RNI112DK_LC_23_15_0  (
            .in0(_gnd_net_),
            .in1(N__62219),
            .in2(N__62060),
            .in3(N__62030),
            .lcout(\ALU.addsub_7 ),
            .ltout(),
            .carryin(bfn_23_15_0_),
            .carryout(\ALU.addsub_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_7_c_RNI7LOOL_LC_23_15_1 .C_ON=1'b1;
    defparam \ALU.addsub_cry_7_c_RNI7LOOL_LC_23_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_7_c_RNI7LOOL_LC_23_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_7_c_RNI7LOOL_LC_23_15_1  (
            .in0(_gnd_net_),
            .in1(N__62027),
            .in2(N__61781),
            .in3(N__61742),
            .lcout(\ALU.addsub_8 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_7 ),
            .carryout(\ALU.addsub_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_8_c_RNINRS3M_LC_23_15_2 .C_ON=1'b1;
    defparam \ALU.addsub_cry_8_c_RNINRS3M_LC_23_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_8_c_RNINRS3M_LC_23_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_8_c_RNINRS3M_LC_23_15_2  (
            .in0(_gnd_net_),
            .in1(N__62801),
            .in2(N__62672),
            .in3(N__61739),
            .lcout(\ALU.addsub_9 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_8 ),
            .carryout(\ALU.addsub_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_9_c_RNI8MSRO_LC_23_15_3 .C_ON=1'b1;
    defparam \ALU.addsub_cry_9_c_RNI8MSRO_LC_23_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_9_c_RNI8MSRO_LC_23_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_9_c_RNI8MSRO_LC_23_15_3  (
            .in0(_gnd_net_),
            .in1(N__61736),
            .in2(N__61710),
            .in3(N__61478),
            .lcout(\ALU.addsub_10 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_9 ),
            .carryout(\ALU.addsub_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_10_c_RNIS0BKM_LC_23_15_4 .C_ON=1'b1;
    defparam \ALU.addsub_cry_10_c_RNIS0BKM_LC_23_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_10_c_RNIS0BKM_LC_23_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_10_c_RNIS0BKM_LC_23_15_4  (
            .in0(_gnd_net_),
            .in1(N__61364),
            .in2(N__61298),
            .in3(N__61247),
            .lcout(\ALU.addsub_11 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_10 ),
            .carryout(\ALU.addsub_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_11_c_RNI0C50P_LC_23_15_5 .C_ON=1'b1;
    defparam \ALU.addsub_cry_11_c_RNI0C50P_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_11_c_RNI0C50P_LC_23_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_11_c_RNI0C50P_LC_23_15_5  (
            .in0(_gnd_net_),
            .in1(N__61244),
            .in2(N__61224),
            .in3(N__61028),
            .lcout(\ALU.addsub_12 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_11 ),
            .carryout(\ALU.addsub_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_12_c_RNIEV1GP_LC_23_15_6 .C_ON=1'b1;
    defparam \ALU.addsub_cry_12_c_RNIEV1GP_LC_23_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_12_c_RNIEV1GP_LC_23_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_12_c_RNIEV1GP_LC_23_15_6  (
            .in0(_gnd_net_),
            .in1(N__61025),
            .in2(N__61019),
            .in3(N__63863),
            .lcout(\ALU.addsub_13 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_12 ),
            .carryout(\ALU.addsub_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_13_c_RNI9HJ8N_LC_23_15_7 .C_ON=1'b1;
    defparam \ALU.addsub_cry_13_c_RNI9HJ8N_LC_23_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_13_c_RNI9HJ8N_LC_23_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_13_c_RNI9HJ8N_LC_23_15_7  (
            .in0(_gnd_net_),
            .in1(N__63860),
            .in2(N__63819),
            .in3(N__63683),
            .lcout(\ALU.addsub_14 ),
            .ltout(),
            .carryin(\ALU.addsub_cry_13 ),
            .carryout(\ALU.addsub_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_14_c_RNIORHUL_LC_23_16_0 .C_ON=1'b1;
    defparam \ALU.addsub_cry_14_c_RNIORHUL_LC_23_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_14_c_RNIORHUL_LC_23_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.addsub_cry_14_c_RNIORHUL_LC_23_16_0  (
            .in0(_gnd_net_),
            .in1(N__63680),
            .in2(N__63612),
            .in3(N__63488),
            .lcout(\ALU.addsub_15 ),
            .ltout(),
            .carryin(bfn_23_16_0_),
            .carryout(\ALU.addsub_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.status_RNO_0_1_LC_23_16_1 .C_ON=1'b0;
    defparam \ALU.status_RNO_0_1_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.status_RNO_0_1_LC_23_16_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \ALU.status_RNO_0_1_LC_23_16_1  (
            .in0(N__63442),
            .in1(N__63239),
            .in2(N__69496),
            .in3(N__63392),
            .lcout(\ALU.N_545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIPBAG72_14_LC_23_16_4 .C_ON=1'b0;
    defparam \ALU.c_RNIPBAG72_14_LC_23_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIPBAG72_14_LC_23_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNIPBAG72_14_LC_23_16_4  (
            .in0(N__69988),
            .in1(N__63360),
            .in2(_gnd_net_),
            .in3(N__62627),
            .lcout(\ALU.c_RNIPBAG72Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI70I1I_9_LC_23_16_6 .C_ON=1'b0;
    defparam \ALU.d_RNI70I1I_9_LC_23_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI70I1I_9_LC_23_16_6 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \ALU.d_RNI70I1I_9_LC_23_16_6  (
            .in0(N__63238),
            .in1(N__62927),
            .in2(_gnd_net_),
            .in3(N__62881),
            .lcout(\ALU.d_RNI70I1IZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNISS7FV1_14_LC_23_16_7 .C_ON=1'b0;
    defparam \ALU.c_RNISS7FV1_14_LC_23_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNISS7FV1_14_LC_23_16_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ALU.c_RNISS7FV1_14_LC_23_16_7  (
            .in0(N__62663),
            .in1(N__68933),
            .in2(_gnd_net_),
            .in3(N__66075),
            .lcout(\ALU.N_1029 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m500_ns_LC_23_17_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m500_ns_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m500_ns_LC_23_17_0 .LUT_INIT=16'b0110010011101100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m500_ns_LC_23_17_0  (
            .in0(N__79497),
            .in1(N__62621),
            .in2(N__63935),
            .in3(N__63869),
            .lcout(\PROM.ROMDATA.m500_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m498_am_LC_23_17_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m498_am_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m498_am_LC_23_17_1 .LUT_INIT=16'b1111111100100111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m498_am_LC_23_17_1  (
            .in0(N__75995),
            .in1(N__78997),
            .in2(N__73919),
            .in3(N__78744),
            .lcout(),
            .ltout(\PROM.ROMDATA.m498_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m498_ns_LC_23_17_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m498_ns_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m498_ns_LC_23_17_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m498_ns_LC_23_17_2  (
            .in0(_gnd_net_),
            .in1(N__63950),
            .in2(N__63938),
            .in3(N__76572),
            .lcout(\PROM.ROMDATA.m498_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m317_bm_LC_23_17_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m317_bm_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m317_bm_LC_23_17_3 .LUT_INIT=16'b0010010010101100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m317_bm_LC_23_17_3  (
            .in0(N__75996),
            .in1(N__78745),
            .in2(N__73918),
            .in3(N__78041),
            .lcout(),
            .ltout(\PROM.ROMDATA.m317_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m317_ns_LC_23_17_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m317_ns_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m317_ns_LC_23_17_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m317_ns_LC_23_17_4  (
            .in0(N__63926),
            .in1(_gnd_net_),
            .in2(N__63914),
            .in3(N__76573),
            .lcout(),
            .ltout(\PROM.ROMDATA.m317_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m325_ns_1_LC_23_17_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m325_ns_1_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m325_ns_1_LC_23_17_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m325_ns_1_LC_23_17_5  (
            .in0(N__63911),
            .in1(N__79498),
            .in2(N__63899),
            .in3(N__79895),
            .lcout(),
            .ltout(\PROM.ROMDATA.m325_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m325_ns_LC_23_17_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m325_ns_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m325_ns_LC_23_17_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m325_ns_LC_23_17_6  (
            .in0(N__79499),
            .in1(N__74912),
            .in2(N__63896),
            .in3(N__63893),
            .lcout(\PROM.ROMDATA.m325_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m329_LC_23_18_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m329_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m329_LC_23_18_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m329_LC_23_18_0  (
            .in0(N__74070),
            .in1(N__72770),
            .in2(N__63884),
            .in3(N__64124),
            .lcout(),
            .ltout(PROM_ROMDATA_dintern_14ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.results_1_LC_23_18_1 .C_ON=1'b0;
    defparam \CONTROL.results_1_LC_23_18_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.results_1_LC_23_18_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \CONTROL.results_1_LC_23_18_1  (
            .in0(N__70882),
            .in1(N__64084),
            .in2(N__63872),
            .in3(N__72299),
            .lcout(aluResults_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.results_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m494_ns_LC_23_18_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m494_ns_LC_23_18_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m494_ns_LC_23_18_2 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m494_ns_LC_23_18_2  (
            .in0(N__73829),
            .in1(N__65192),
            .in2(N__73469),
            .in3(N__76575),
            .lcout(\PROM.ROMDATA.m494_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m414_ns_LC_23_18_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m414_ns_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m414_ns_LC_23_18_3 .LUT_INIT=16'b1011100100110001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m414_ns_LC_23_18_3  (
            .in0(N__76574),
            .in1(N__64187),
            .in2(N__64181),
            .in3(N__64346),
            .lcout(\PROM.ROMDATA.m414_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m308_LC_23_18_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m308_LC_23_18_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m308_LC_23_18_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m308_LC_23_18_4  (
            .in0(N__74069),
            .in1(N__74258),
            .in2(N__64157),
            .in3(N__72771),
            .lcout(),
            .ltout(PROM_ROMDATA_dintern_13ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.results_0_LC_23_18_5 .C_ON=1'b0;
    defparam \CONTROL.results_0_LC_23_18_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.results_0_LC_23_18_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \CONTROL.results_0_LC_23_18_5  (
            .in0(N__69270),
            .in1(N__64083),
            .in2(N__64145),
            .in3(N__72298),
            .lcout(aluResults_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.results_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m198_LC_23_19_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m198_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m198_LC_23_19_0 .LUT_INIT=16'b0000001010010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m198_LC_23_19_0  (
            .in0(N__78404),
            .in1(N__77896),
            .in2(N__75954),
            .in3(N__77252),
            .lcout(\PROM.ROMDATA.m198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m344_LC_23_19_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m344_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m344_LC_23_19_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m344_LC_23_19_1  (
            .in0(N__72697),
            .in1(N__74067),
            .in2(N__79064),
            .in3(N__64123),
            .lcout(),
            .ltout(PROM_ROMDATA_dintern_15ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.results_2_LC_23_19_2 .C_ON=1'b0;
    defparam \CONTROL.results_2_LC_23_19_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.results_2_LC_23_19_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \CONTROL.results_2_LC_23_19_2  (
            .in0(N__70913),
            .in1(N__64085),
            .in2(N__64070),
            .in3(N__72304),
            .lcout(aluResults_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.results_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m367_LC_23_19_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m367_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m367_LC_23_19_3 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m367_LC_23_19_3  (
            .in0(N__65013),
            .in1(N__74066),
            .in2(N__64067),
            .in3(N__75800),
            .lcout(\PROM.ROMDATA.N_564_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m298_bm_LC_23_19_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m298_bm_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m298_bm_LC_23_19_4 .LUT_INIT=16'b0110001100101100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m298_bm_LC_23_19_4  (
            .in0(N__78406),
            .in1(N__77898),
            .in2(N__75955),
            .in3(N__77255),
            .lcout(\PROM.ROMDATA.m298_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m386_LC_23_19_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m386_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m386_LC_23_19_5 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m386_LC_23_19_5  (
            .in0(N__74068),
            .in1(N__64261),
            .in2(N__64018),
            .in3(N__75804),
            .lcout(\PROM.ROMDATA.N_565_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m287_LC_23_19_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m287_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m287_LC_23_19_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m287_LC_23_19_6  (
            .in0(N__78405),
            .in1(N__77897),
            .in2(_gnd_net_),
            .in3(N__77253),
            .lcout(\PROM.ROMDATA.m287 ),
            .ltout(\PROM.ROMDATA.m287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m410_bm_LC_23_19_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m410_bm_LC_23_19_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m410_bm_LC_23_19_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m410_bm_LC_23_19_7  (
            .in0(N__77254),
            .in1(N__77940),
            .in2(N__64349),
            .in3(N__75799),
            .lcout(\PROM.ROMDATA.m410_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m66_LC_23_20_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m66_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m66_LC_23_20_0 .LUT_INIT=16'b0011000011111010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m66_LC_23_20_0  (
            .in0(N__77250),
            .in1(N__75668),
            .in2(N__78021),
            .in3(N__78359),
            .lcout(\PROM.ROMDATA.m66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m490_LC_23_20_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m490_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m490_LC_23_20_1 .LUT_INIT=16'b1000100001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m490_LC_23_20_1  (
            .in0(N__75669),
            .in1(N__74963),
            .in2(N__64328),
            .in3(N__76404),
            .lcout(\PROM.ROMDATA.m490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m446_am_LC_23_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m446_am_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m446_am_LC_23_20_2 .LUT_INIT=16'b1000000001000001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m446_am_LC_23_20_2  (
            .in0(N__77251),
            .in1(N__75672),
            .in2(N__78022),
            .in3(N__78361),
            .lcout(\PROM.ROMDATA.m446_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m149_LC_23_20_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m149_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m149_LC_23_20_3 .LUT_INIT=16'b0101010111101110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m149_LC_23_20_3  (
            .in0(N__78358),
            .in1(N__77899),
            .in2(_gnd_net_),
            .in3(N__77249),
            .lcout(\PROM.ROMDATA.m149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m120_bm_LC_23_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m120_bm_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m120_bm_LC_23_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m120_bm_LC_23_20_4  (
            .in0(N__76403),
            .in1(N__64277),
            .in2(_gnd_net_),
            .in3(N__64271),
            .lcout(\PROM.ROMDATA.m120_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m456_ns_1_LC_23_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m456_ns_1_LC_23_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m456_ns_1_LC_23_20_5 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m456_ns_1_LC_23_20_5  (
            .in0(N__75670),
            .in1(N__64793),
            .in2(N__79891),
            .in3(N__64966),
            .lcout(),
            .ltout(\PROM.ROMDATA.m456_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m456_ns_LC_23_20_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m456_ns_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m456_ns_LC_23_20_6 .LUT_INIT=16'b0100100000001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m456_ns_LC_23_20_6  (
            .in0(N__76405),
            .in1(N__64250),
            .in2(N__64202),
            .in3(N__75671),
            .lcout(\PROM.ROMDATA.m456_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m166_e_LC_23_20_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m166_e_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m166_e_LC_23_20_7 .LUT_INIT=16'b0000000101010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m166_e_LC_23_20_7  (
            .in0(N__78360),
            .in1(N__64524),
            .in2(N__73740),
            .in3(N__64486),
            .lcout(\PROM.ROMDATA.m166_e ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m107_LC_23_21_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m107_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m107_LC_23_21_0 .LUT_INIT=16'b0110100010111010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m107_LC_23_21_0  (
            .in0(N__78482),
            .in1(N__77966),
            .in2(N__75795),
            .in3(N__77244),
            .lcout(\PROM.ROMDATA.m107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m361_am_LC_23_21_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m361_am_LC_23_21_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m361_am_LC_23_21_1 .LUT_INIT=16'b1111101100111000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m361_am_LC_23_21_1  (
            .in0(N__77245),
            .in1(N__75500),
            .in2(N__78573),
            .in3(N__79033),
            .lcout(\PROM.ROMDATA.m361_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m104_ns_LC_23_21_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m104_ns_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m104_ns_LC_23_21_2 .LUT_INIT=16'b0101010111100100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m104_ns_LC_23_21_2  (
            .in0(N__75499),
            .in1(N__78988),
            .in2(N__79043),
            .in3(N__64433),
            .lcout(),
            .ltout(\PROM.ROMDATA.m104_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m109_bm_LC_23_21_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m109_bm_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m109_bm_LC_23_21_3 .LUT_INIT=16'b0011001111110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m109_bm_LC_23_21_3  (
            .in0(_gnd_net_),
            .in1(N__64424),
            .in2(N__64418),
            .in3(N__76272),
            .lcout(),
            .ltout(\PROM.ROMDATA.m109_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m121_ns_LC_23_21_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m121_ns_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m121_ns_LC_23_21_4 .LUT_INIT=16'b0101010111011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m121_ns_LC_23_21_4  (
            .in0(N__64355),
            .in1(N__64415),
            .in2(N__64400),
            .in3(N__79322),
            .lcout(\PROM.ROMDATA.m121_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m357_bm_LC_23_21_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m357_bm_LC_23_21_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m357_bm_LC_23_21_5 .LUT_INIT=16'b0001100111100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m357_bm_LC_23_21_5  (
            .in0(N__77246),
            .in1(N__75501),
            .in2(N__78043),
            .in3(N__78483),
            .lcout(\PROM.ROMDATA.m357_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m120_am_LC_23_21_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m120_am_LC_23_21_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m120_am_LC_23_21_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m120_am_LC_23_21_6  (
            .in0(N__76271),
            .in1(N__64376),
            .in2(_gnd_net_),
            .in3(N__64370),
            .lcout(),
            .ltout(\PROM.ROMDATA.m120_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m121_ns_1_LC_23_21_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m121_ns_1_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m121_ns_1_LC_23_21_7 .LUT_INIT=16'b0001001110011011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m121_ns_1_LC_23_21_7  (
            .in0(N__79321),
            .in1(N__79834),
            .in2(N__64364),
            .in3(N__64361),
            .lcout(\PROM.ROMDATA.m121_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m138_LC_23_22_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m138_LC_23_22_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m138_LC_23_22_0 .LUT_INIT=16'b0111010011110001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m138_LC_23_22_0  (
            .in0(N__78334),
            .in1(N__77692),
            .in2(N__75909),
            .in3(N__77067),
            .lcout(),
            .ltout(\PROM.ROMDATA.m138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m147_am_LC_23_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m147_am_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m147_am_LC_23_22_1 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m147_am_LC_23_22_1  (
            .in0(_gnd_net_),
            .in1(N__64769),
            .in2(N__64763),
            .in3(N__76350),
            .lcout(\PROM.ROMDATA.m147_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m80_bm_1_LC_23_22_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m80_bm_1_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m80_bm_1_LC_23_22_2 .LUT_INIT=16'b0100010001100111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m80_bm_1_LC_23_22_2  (
            .in0(N__78333),
            .in1(N__77690),
            .in2(N__76498),
            .in3(N__77065),
            .lcout(),
            .ltout(\PROM.ROMDATA.m80_bm_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m80_bm_LC_23_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m80_bm_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m80_bm_LC_23_22_3 .LUT_INIT=16'b0011110010100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m80_bm_LC_23_22_3  (
            .in0(N__77691),
            .in1(N__76349),
            .in2(N__64760),
            .in3(N__75711),
            .lcout(\PROM.ROMDATA.m80_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m4_LC_23_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m4_LC_23_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m4_LC_23_22_4 .LUT_INIT=16'b0011010111001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m4_LC_23_22_4  (
            .in0(N__64740),
            .in1(N__64710),
            .in2(N__64662),
            .in3(N__77066),
            .lcout(\PROM.ROMDATA.m4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m347_LC_23_22_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m347_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m347_LC_23_22_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m347_LC_23_22_5  (
            .in0(N__77069),
            .in1(N__78336),
            .in2(_gnd_net_),
            .in3(N__77744),
            .lcout(\PROM.ROMDATA.m347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m292_LC_23_22_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m292_LC_23_22_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m292_LC_23_22_6 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m292_LC_23_22_6  (
            .in0(N__73552),
            .in1(N__73809),
            .in2(N__73730),
            .in3(N__77070),
            .lcout(\PROM.ROMDATA.m292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m112_LC_23_22_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m112_LC_23_22_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m112_LC_23_22_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m112_LC_23_22_7  (
            .in0(N__77068),
            .in1(N__78335),
            .in2(_gnd_net_),
            .in3(N__77743),
            .lcout(\PROM.ROMDATA.m112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m137_bm_LC_23_23_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m137_bm_LC_23_23_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m137_bm_LC_23_23_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m137_bm_LC_23_23_0  (
            .in0(N__76263),
            .in1(N__64544),
            .in2(_gnd_net_),
            .in3(N__64538),
            .lcout(\PROM.ROMDATA.m137_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m83_LC_23_23_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m83_LC_23_23_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m83_LC_23_23_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m83_LC_23_23_1  (
            .in0(N__78793),
            .in1(N__77888),
            .in2(_gnd_net_),
            .in3(N__77238),
            .lcout(\PROM.ROMDATA.m83 ),
            .ltout(\PROM.ROMDATA.m83_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m161_LC_23_23_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m161_LC_23_23_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m161_LC_23_23_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m161_LC_23_23_2  (
            .in0(N__76261),
            .in1(N__75636),
            .in2(N__64976),
            .in3(N__64940),
            .lcout(\PROM.ROMDATA.m161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m15_LC_23_23_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m15_LC_23_23_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m15_LC_23_23_3 .LUT_INIT=16'b0110011000010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m15_LC_23_23_3  (
            .in0(N__78792),
            .in1(N__77887),
            .in2(_gnd_net_),
            .in3(N__77237),
            .lcout(\PROM.ROMDATA.m15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m128_LC_23_23_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m128_LC_23_23_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m128_LC_23_23_4 .LUT_INIT=16'b0000101010101101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m128_LC_23_23_4  (
            .in0(N__77239),
            .in1(N__75637),
            .in2(N__78020),
            .in3(N__78794),
            .lcout(\PROM.ROMDATA.m128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m171_ns_LC_23_23_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m171_ns_LC_23_23_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m171_ns_LC_23_23_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m171_ns_LC_23_23_5  (
            .in0(N__64778),
            .in1(_gnd_net_),
            .in2(N__79890),
            .in3(N__65102),
            .lcout(),
            .ltout(\PROM.ROMDATA.m171_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m172_LC_23_23_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m172_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m172_LC_23_23_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m172_LC_23_23_6  (
            .in0(N__79454),
            .in1(_gnd_net_),
            .in2(N__64913),
            .in3(N__64910),
            .lcout(\PROM.ROMDATA.m172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m171_bm_LC_23_23_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m171_bm_LC_23_23_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m171_bm_LC_23_23_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m171_bm_LC_23_23_7  (
            .in0(N__75638),
            .in1(N__76262),
            .in2(N__64876),
            .in3(N__64789),
            .lcout(\PROM.ROMDATA.m171_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m383_LC_23_24_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m383_LC_23_24_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m383_LC_23_24_0 .LUT_INIT=16'b0010100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m383_LC_23_24_0  (
            .in0(N__77886),
            .in1(N__77236),
            .in2(N__75900),
            .in3(N__78506),
            .lcout(),
            .ltout(\PROM.ROMDATA.m383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m427_am_LC_23_24_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m427_am_LC_23_24_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m427_am_LC_23_24_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m427_am_LC_23_24_1  (
            .in0(N__76448),
            .in1(N__74406),
            .in2(N__64772),
            .in3(N__75684),
            .lcout(),
            .ltout(\PROM.ROMDATA.m427_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m427_ns_LC_23_24_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m427_ns_LC_23_24_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m427_ns_LC_23_24_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m427_ns_LC_23_24_2  (
            .in0(_gnd_net_),
            .in1(N__65249),
            .in2(N__65240),
            .in3(N__79857),
            .lcout(\PROM.ROMDATA.m427_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m494_ns_1_LC_23_24_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m494_ns_1_LC_23_24_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m494_ns_1_LC_23_24_3 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m494_ns_1_LC_23_24_3  (
            .in0(N__76447),
            .in1(N__65213),
            .in2(N__65201),
            .in3(N__75680),
            .lcout(\PROM.ROMDATA.m494_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m88_LC_23_24_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m88_LC_23_24_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m88_LC_23_24_4 .LUT_INIT=16'b0001001100111001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m88_LC_23_24_4  (
            .in0(N__77884),
            .in1(N__77234),
            .in2(N__75899),
            .in3(N__78505),
            .lcout(\PROM.ROMDATA.m88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m181_LC_23_24_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m181_LC_23_24_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m181_LC_23_24_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m181_LC_23_24_5  (
            .in0(N__77235),
            .in1(N__78542),
            .in2(_gnd_net_),
            .in3(N__77885),
            .lcout(\PROM.ROMDATA.m181 ),
            .ltout(\PROM.ROMDATA.m181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m514_ns_LC_23_24_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m514_ns_LC_23_24_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m514_ns_LC_23_24_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m514_ns_LC_23_24_6  (
            .in0(N__74489),
            .in1(N__65171),
            .in2(N__65153),
            .in3(N__79487),
            .lcout(\PROM.ROMDATA.m514_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m171_am_LC_23_24_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m171_am_LC_23_24_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m171_am_LC_23_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m171_am_LC_23_24_7  (
            .in0(N__76446),
            .in1(N__65114),
            .in2(_gnd_net_),
            .in3(N__65108),
            .lcout(\PROM.ROMDATA.m171_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_12_LC_24_10_0 .C_ON=1'b0;
    defparam \ALU.d_12_LC_24_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.d_12_LC_24_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_12_LC_24_10_0  (
            .in0(N__67756),
            .in1(N__67686),
            .in2(_gnd_net_),
            .in3(N__67621),
            .lcout(\ALU.dZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73177),
            .ce(N__70239),
            .sr(_gnd_net_));
    defparam \ALU.d_13_LC_24_10_1 .C_ON=1'b0;
    defparam \ALU.d_13_LC_24_10_1 .SEQ_MODE=4'b1000;
    defparam \ALU.d_13_LC_24_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_13_LC_24_10_1  (
            .in0(N__67451),
            .in1(N__67508),
            .in2(_gnd_net_),
            .in3(N__67389),
            .lcout(\ALU.dZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73177),
            .ce(N__70239),
            .sr(_gnd_net_));
    defparam \ALU.d_14_LC_24_10_2 .C_ON=1'b0;
    defparam \ALU.d_14_LC_24_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.d_14_LC_24_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_14_LC_24_10_2  (
            .in0(N__68144),
            .in1(N__68077),
            .in2(_gnd_net_),
            .in3(N__68012),
            .lcout(\ALU.dZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73177),
            .ce(N__70239),
            .sr(_gnd_net_));
    defparam \ALU.c_12_LC_24_11_0 .C_ON=1'b0;
    defparam \ALU.c_12_LC_24_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.c_12_LC_24_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_12_LC_24_11_0  (
            .in0(N__67753),
            .in1(N__67685),
            .in2(_gnd_net_),
            .in3(N__67610),
            .lcout(\ALU.cZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73188),
            .ce(N__71553),
            .sr(_gnd_net_));
    defparam \ALU.c_13_LC_24_11_1 .C_ON=1'b0;
    defparam \ALU.c_13_LC_24_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.c_13_LC_24_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.c_13_LC_24_11_1  (
            .in0(N__67516),
            .in1(N__67459),
            .in2(_gnd_net_),
            .in3(N__67391),
            .lcout(\ALU.cZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73188),
            .ce(N__71553),
            .sr(_gnd_net_));
    defparam \ALU.c_14_LC_24_11_2 .C_ON=1'b0;
    defparam \ALU.c_14_LC_24_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.c_14_LC_24_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_14_LC_24_11_2  (
            .in0(N__68136),
            .in1(N__68076),
            .in2(_gnd_net_),
            .in3(N__68003),
            .lcout(\ALU.cZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73188),
            .ce(N__71553),
            .sr(_gnd_net_));
    defparam \ALU.addsub_cry_8_c_RNI6UUIV5_LC_24_13_0 .C_ON=1'b0;
    defparam \ALU.addsub_cry_8_c_RNI6UUIV5_LC_24_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.addsub_cry_8_c_RNI6UUIV5_LC_24_13_0 .LUT_INIT=16'b0011000000111010;
    LogicCell40 \ALU.addsub_cry_8_c_RNI6UUIV5_LC_24_13_0  (
            .in0(N__67164),
            .in1(N__68150),
            .in2(N__66897),
            .in3(N__66860),
            .lcout(\ALU.a_15_d_ns_sx_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMGKJC1_0_2_LC_24_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIMGKJC1_0_2_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMGKJC1_0_2_LC_24_13_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \ALU.d_RNIMGKJC1_0_2_LC_24_13_1  (
            .in0(N__66315),
            .in1(N__66085),
            .in2(N__65585),
            .in3(N__66761),
            .lcout(\ALU.d_RNIMGKJC1_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMGKJC1_2_LC_24_13_2 .C_ON=1'b0;
    defparam \ALU.d_RNIMGKJC1_2_LC_24_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMGKJC1_2_LC_24_13_2 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \ALU.d_RNIMGKJC1_2_LC_24_13_2  (
            .in0(N__66762),
            .in1(N__66316),
            .in2(N__66089),
            .in3(N__65584),
            .lcout(),
            .ltout(\ALU.d_RNIMGKJC1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0TK6H3_2_LC_24_13_3 .C_ON=1'b0;
    defparam \ALU.d_RNI0TK6H3_2_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0TK6H3_2_LC_24_13_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.d_RNI0TK6H3_2_LC_24_13_3  (
            .in0(_gnd_net_),
            .in1(N__65285),
            .in2(N__65279),
            .in3(N__65272),
            .lcout(),
            .ltout(\ALU.N_859_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISGV438_2_LC_24_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNISGV438_2_LC_24_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISGV438_2_LC_24_13_4 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.d_RNISGV438_2_LC_24_13_4  (
            .in0(N__69188),
            .in1(N__68521),
            .in2(N__69176),
            .in3(N__68897),
            .lcout(),
            .ltout(\ALU.rshift_15_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI0UFMPC_15_LC_24_13_5 .C_ON=1'b0;
    defparam \ALU.c_RNI0UFMPC_15_LC_24_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI0UFMPC_15_LC_24_13_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNI0UFMPC_15_LC_24_13_5  (
            .in0(N__68522),
            .in1(N__68567),
            .in2(N__69173),
            .in3(N__68167),
            .lcout(),
            .ltout(\ALU.rshift_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI98D92D_15_LC_24_13_6 .C_ON=1'b0;
    defparam \ALU.c_RNI98D92D_15_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI98D92D_15_LC_24_13_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.c_RNI98D92D_15_LC_24_13_6  (
            .in0(N__69150),
            .in1(_gnd_net_),
            .in2(N__69077),
            .in3(N__69057),
            .lcout(\ALU.c_RNI98D92DZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNICBIG85_15_LC_24_13_7 .C_ON=1'b0;
    defparam \ALU.c_RNICBIG85_15_LC_24_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNICBIG85_15_LC_24_13_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.c_RNICBIG85_15_LC_24_13_7  (
            .in0(N__68896),
            .in1(N__68566),
            .in2(N__68531),
            .in3(N__68166),
            .lcout(\ALU.c_RNICBIG85Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_14_LC_24_14_0 .C_ON=1'b0;
    defparam \ALU.b_14_LC_24_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.b_14_LC_24_14_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_14_LC_24_14_0  (
            .in0(N__68140),
            .in1(N__68079),
            .in2(_gnd_net_),
            .in3(N__68011),
            .lcout(\ALU.bZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73209),
            .ce(N__67921),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_8_LC_24_15_0 .C_ON=1'b0;
    defparam \ALU.un1_a41_8_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_8_LC_24_15_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ALU.un1_a41_8_LC_24_15_0  (
            .in0(N__70268),
            .in1(N__70891),
            .in2(N__69338),
            .in3(N__69284),
            .lcout(\ALU.un1_a41_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_4_LC_24_15_1 .C_ON=1'b0;
    defparam \ALU.un1_a41_4_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_4_LC_24_15_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ALU.un1_a41_4_LC_24_15_1  (
            .in0(N__70889),
            .in1(N__69333),
            .in2(N__70942),
            .in3(N__70259),
            .lcout(\ALU.un1_a41_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_operation_10_LC_24_15_2 .C_ON=1'b0;
    defparam \ALU.un1_operation_10_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_operation_10_LC_24_15_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \ALU.un1_operation_10_LC_24_15_2  (
            .in0(N__67820),
            .in1(N__69966),
            .in2(N__67808),
            .in3(N__69799),
            .lcout(\ALU.un1_operation_10_0 ),
            .ltout(\ALU.un1_operation_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_7_2_LC_24_15_3 .C_ON=1'b0;
    defparam \ALU.un1_a41_7_2_LC_24_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_7_2_LC_24_15_3 .LUT_INIT=16'b0101000100010001;
    LogicCell40 \ALU.un1_a41_7_2_LC_24_15_3  (
            .in0(N__70931),
            .in1(N__71515),
            .in2(N__67787),
            .in3(N__71469),
            .lcout(\ALU.un1_a41_7_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_operation_13_2_LC_24_15_4 .C_ON=1'b0;
    defparam \ALU.un1_operation_13_2_LC_24_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_operation_13_2_LC_24_15_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ALU.un1_operation_13_2_LC_24_15_4  (
            .in0(N__69967),
            .in1(N__69798),
            .in2(N__69716),
            .in3(N__70157),
            .lcout(\ALU.un1_operation_13Z0Z_2 ),
            .ltout(\ALU.un1_operation_13Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_4_2_LC_24_15_5 .C_ON=1'b0;
    defparam \ALU.un1_a41_4_2_LC_24_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_4_2_LC_24_15_5 .LUT_INIT=16'b1000101000001010;
    LogicCell40 \ALU.un1_a41_4_2_LC_24_15_5  (
            .in0(N__69283),
            .in1(N__71491),
            .in2(N__70262),
            .in3(N__71468),
            .lcout(\ALU.un1_a41_4_0_2 ),
            .ltout(\ALU.un1_a41_4_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_6_LC_24_15_6 .C_ON=1'b0;
    defparam \ALU.un1_a41_6_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_6_LC_24_15_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ALU.un1_a41_6_LC_24_15_6  (
            .in0(N__69337),
            .in1(N__70935),
            .in2(N__70253),
            .in3(N__70890),
            .lcout(\ALU.un1_a41_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_operation_7_LC_24_15_7 .C_ON=1'b0;
    defparam \ALU.un1_operation_7_LC_24_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_operation_7_LC_24_15_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ALU.un1_operation_7_LC_24_15_7  (
            .in0(N__70158),
            .in1(N__69968),
            .in2(N__69803),
            .in3(N__69697),
            .lcout(\ALU.un1_operationZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_2_LC_24_16_0 .C_ON=1'b0;
    defparam \ALU.un1_a41_2_LC_24_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_2_LC_24_16_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ALU.un1_a41_2_LC_24_16_0  (
            .in0(N__71007),
            .in1(N__69332),
            .in2(N__70844),
            .in3(N__69282),
            .lcout(\ALU.un1_a41_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m160_LC_24_16_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m160_LC_24_16_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m160_LC_24_16_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m160_LC_24_16_1  (
            .in0(N__78842),
            .in1(N__78066),
            .in2(N__76003),
            .in3(N__77317),
            .lcout(\PROM.ROMDATA.m160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_3_1_LC_24_16_2 .C_ON=1'b0;
    defparam \ALU.un1_a41_3_1_LC_24_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_3_1_LC_24_16_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ALU.un1_a41_3_1_LC_24_16_2  (
            .in0(_gnd_net_),
            .in1(N__69331),
            .in2(_gnd_net_),
            .in3(N__69281),
            .lcout(\ALU.un1_a41_3_0_1 ),
            .ltout(\ALU.un1_a41_3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_5_LC_24_16_3 .C_ON=1'b0;
    defparam \ALU.un1_a41_5_LC_24_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_5_LC_24_16_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.un1_a41_5_LC_24_16_3  (
            .in0(N__70940),
            .in1(N__70883),
            .in2(N__69248),
            .in3(N__71008),
            .lcout(\ALU.un1_a41_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_7_LC_24_16_4 .C_ON=1'b0;
    defparam \ALU.un1_a41_7_LC_24_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_7_LC_24_16_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ALU.un1_a41_7_LC_24_16_4  (
            .in0(N__71009),
            .in1(N__70941),
            .in2(N__70892),
            .in3(N__71019),
            .lcout(\ALU.un1_a41_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_operation_13_LC_24_16_5 .C_ON=1'b0;
    defparam \ALU.un1_operation_13_LC_24_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_operation_13_LC_24_16_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \ALU.un1_operation_13_LC_24_16_5  (
            .in0(N__71519),
            .in1(N__71490),
            .in2(_gnd_net_),
            .in3(N__71470),
            .lcout(\ALU.un1_operation_13_0 ),
            .ltout(\ALU.un1_operation_13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_9_LC_24_16_6 .C_ON=1'b0;
    defparam \ALU.un1_a41_9_LC_24_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_9_LC_24_16_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ALU.un1_a41_9_LC_24_16_6  (
            .in0(N__70887),
            .in1(N__70936),
            .in2(N__71219),
            .in3(N__71020),
            .lcout(\ALU.un1_a41_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_3_LC_24_16_7 .C_ON=1'b0;
    defparam \ALU.un1_a41_3_LC_24_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_3_LC_24_16_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ALU.un1_a41_3_LC_24_16_7  (
            .in0(N__71021),
            .in1(N__70888),
            .in2(N__70943),
            .in3(N__71006),
            .lcout(\ALU.un1_a41_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un1_a41_2_1_LC_24_17_0 .C_ON=1'b0;
    defparam \ALU.un1_a41_2_1_LC_24_17_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un1_a41_2_1_LC_24_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.un1_a41_2_1_LC_24_17_0  (
            .in0(_gnd_net_),
            .in1(N__70914),
            .in2(_gnd_net_),
            .in3(N__70865),
            .lcout(\ALU.un1_a41_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.ramAddReg_6_LC_24_18_3 .C_ON=1'b0;
    defparam \CONTROL.ramAddReg_6_LC_24_18_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.ramAddReg_6_LC_24_18_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \CONTROL.ramAddReg_6_LC_24_18_3  (
            .in0(N__70835),
            .in1(N__70799),
            .in2(N__70613),
            .in3(N__70556),
            .lcout(A6_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVCONTROL.ramAddReg_6C_net ),
            .ce(N__70329),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m281_LC_24_19_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m281_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m281_LC_24_19_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m281_LC_24_19_0  (
            .in0(N__78714),
            .in1(N__77907),
            .in2(_gnd_net_),
            .in3(N__77257),
            .lcout(),
            .ltout(\PROM.ROMDATA.m281_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m480_bm_LC_24_19_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m480_bm_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m480_bm_LC_24_19_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m480_bm_LC_24_19_1  (
            .in0(_gnd_net_),
            .in1(N__76559),
            .in2(N__70271),
            .in3(N__75808),
            .lcout(\PROM.ROMDATA.m480_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m60_LC_24_19_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m60_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m60_LC_24_19_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m60_LC_24_19_2  (
            .in0(N__78713),
            .in1(N__77906),
            .in2(_gnd_net_),
            .in3(N__77256),
            .lcout(\PROM.ROMDATA.m60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.programCounter_ret_1_7_LC_24_19_3 .C_ON=1'b0;
    defparam \CONTROL.programCounter_ret_1_7_LC_24_19_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.programCounter_ret_1_7_LC_24_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.programCounter_ret_1_7_LC_24_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__73355),
            .lcout(\CONTROL.programCounter_1_reto_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__73258),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m480_am_LC_24_19_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m480_am_LC_24_19_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m480_am_LC_24_19_4 .LUT_INIT=16'b0101100000001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m480_am_LC_24_19_4  (
            .in0(N__75809),
            .in1(N__72827),
            .in2(N__76616),
            .in3(N__74488),
            .lcout(),
            .ltout(\PROM.ROMDATA.m480_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m480_ns_LC_24_19_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m480_ns_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m480_ns_LC_24_19_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m480_ns_LC_24_19_5  (
            .in0(_gnd_net_),
            .in1(N__72815),
            .in2(N__72809),
            .in3(N__79898),
            .lcout(),
            .ltout(\PROM.ROMDATA.m480_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m485_LC_24_19_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m485_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m485_LC_24_19_6 .LUT_INIT=16'b0010001010111000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m485_LC_24_19_6  (
            .in0(N__72806),
            .in1(N__72696),
            .in2(N__72383),
            .in3(N__79502),
            .lcout(PROM_ROMDATA_dintern_25ro),
            .ltout(PROM_ROMDATA_dintern_25ro_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.romAddReg_7_9_LC_24_19_7 .C_ON=1'b0;
    defparam \CONTROL.romAddReg_7_9_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \CONTROL.romAddReg_7_9_LC_24_19_7 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \CONTROL.romAddReg_7_9_LC_24_19_7  (
            .in0(N__72352),
            .in1(N__72318),
            .in2(N__71879),
            .in3(N__71875),
            .lcout(CONTROL_romAddReg_7_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m262_LC_24_20_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m262_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m262_LC_24_20_1 .LUT_INIT=16'b0000100000000100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m262_LC_24_20_1  (
            .in0(N__77247),
            .in1(N__75891),
            .in2(N__78839),
            .in3(N__77908),
            .lcout(\PROM.ROMDATA.m262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m447_ns_LC_24_20_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m447_ns_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m447_ns_LC_24_20_2 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m447_ns_LC_24_20_2  (
            .in0(N__71615),
            .in1(N__71603),
            .in2(N__71588),
            .in3(N__79866),
            .lcout(\PROM.ROMDATA.m447_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m488_ns_1_LC_24_20_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m488_ns_1_LC_24_20_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m488_ns_1_LC_24_20_4 .LUT_INIT=16'b0001000101010010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m488_ns_1_LC_24_20_4  (
            .in0(N__75892),
            .in1(N__78718),
            .in2(N__76601),
            .in3(N__77248),
            .lcout(\PROM.ROMDATA.m488_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m503_LC_24_20_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m503_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m503_LC_24_20_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m503_LC_24_20_5  (
            .in0(N__78719),
            .in1(N__74071),
            .in2(N__75986),
            .in3(N__73505),
            .lcout(\PROM.ROMDATA.N_570_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m493_am_LC_24_20_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m493_am_LC_24_20_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m493_am_LC_24_20_6 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m493_am_LC_24_20_6  (
            .in0(N__73728),
            .in1(N__73565),
            .in2(N__73911),
            .in3(N__73812),
            .lcout(\PROM.ROMDATA.m493_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m493_bm_LC_24_20_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m493_bm_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m493_bm_LC_24_20_7 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m493_bm_LC_24_20_7  (
            .in0(N__73813),
            .in1(N__73729),
            .in2(N__73573),
            .in3(N__73504),
            .lcout(\PROM.ROMDATA.m493_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m361_ns_LC_24_21_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m361_ns_LC_24_21_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m361_ns_LC_24_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m361_ns_LC_24_21_0  (
            .in0(N__74192),
            .in1(N__73454),
            .in2(_gnd_net_),
            .in3(N__76522),
            .lcout(\PROM.ROMDATA.m361_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m211_ns_LC_24_21_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m211_ns_LC_24_21_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m211_ns_LC_24_21_1 .LUT_INIT=16'b0000011010110100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m211_ns_LC_24_21_1  (
            .in0(N__78473),
            .in1(N__77961),
            .in2(N__73448),
            .in3(N__77241),
            .lcout(\PROM.ROMDATA.m211_ns ),
            .ltout(\PROM.ROMDATA.m211_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m221cf0_1_LC_24_21_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf0_1_LC_24_21_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf0_1_LC_24_21_2 .LUT_INIT=16'b0011001111000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m221cf0_1_LC_24_21_2  (
            .in0(_gnd_net_),
            .in1(N__79323),
            .in2(N__73436),
            .in3(N__79831),
            .lcout(\PROM.ROMDATA.m221cf0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m221cf1_1_LC_24_21_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf1_1_LC_24_21_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m221cf1_1_LC_24_21_3 .LUT_INIT=16'b0000111101011111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m221cf1_1_LC_24_21_3  (
            .in0(N__79832),
            .in1(_gnd_net_),
            .in2(N__79414),
            .in3(N__73418),
            .lcout(\PROM.ROMDATA.m221cf1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m369_LC_24_21_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m369_LC_24_21_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m369_LC_24_21_4 .LUT_INIT=16'b0101011111100011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m369_LC_24_21_4  (
            .in0(N__77242),
            .in1(N__75810),
            .in2(N__78042),
            .in3(N__78474),
            .lcout(\PROM.ROMDATA.m369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m373_LC_24_21_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m373_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m373_LC_24_21_5 .LUT_INIT=16'b0100001001000101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m373_LC_24_21_5  (
            .in0(N__78475),
            .in1(N__77965),
            .in2(N__75959),
            .in3(N__77243),
            .lcout(\PROM.ROMDATA.m373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m303_ns_LC_24_21_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m303_ns_LC_24_21_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m303_ns_LC_24_21_6 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m303_ns_LC_24_21_6  (
            .in0(N__74270),
            .in1(N__79327),
            .in2(N__74360),
            .in3(N__74093),
            .lcout(\PROM.ROMDATA.m303_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m424_LC_24_21_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m424_LC_24_21_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m424_LC_24_21_7 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m424_LC_24_21_7  (
            .in0(N__79833),
            .in1(N__74239),
            .in2(_gnd_net_),
            .in3(N__74225),
            .lcout(\PROM.ROMDATA.m424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m361_bm_LC_24_22_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m361_bm_LC_24_22_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m361_bm_LC_24_22_0 .LUT_INIT=16'b0011010110111111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m361_bm_LC_24_22_0  (
            .in0(N__77172),
            .in1(N__75718),
            .in2(N__78035),
            .in3(N__78858),
            .lcout(\PROM.ROMDATA.m361_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m137_am_LC_24_22_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m137_am_LC_24_22_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m137_am_LC_24_22_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m137_am_LC_24_22_1  (
            .in0(N__74186),
            .in1(N__76372),
            .in2(_gnd_net_),
            .in3(N__74171),
            .lcout(),
            .ltout(\PROM.ROMDATA.m137_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m148_ns_1_LC_24_22_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m148_ns_1_LC_24_22_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m148_ns_1_LC_24_22_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m148_ns_1_LC_24_22_2  (
            .in0(N__79452),
            .in1(N__79858),
            .in2(N__74165),
            .in3(N__74162),
            .lcout(),
            .ltout(\PROM.ROMDATA.m148_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m148_ns_LC_24_22_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m148_ns_LC_24_22_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m148_ns_LC_24_22_3 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m148_ns_LC_24_22_3  (
            .in0(N__74156),
            .in1(N__74150),
            .in2(N__74141),
            .in3(N__79453),
            .lcout(\PROM.ROMDATA.m148_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m301_LC_24_22_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m301_LC_24_22_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m301_LC_24_22_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m301_LC_24_22_4  (
            .in0(N__76374),
            .in1(N__74125),
            .in2(N__74108),
            .in3(N__75720),
            .lcout(\PROM.ROMDATA.m301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m349_am_LC_24_22_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m349_am_LC_24_22_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m349_am_LC_24_22_5 .LUT_INIT=16'b1001111101110101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m349_am_LC_24_22_5  (
            .in0(N__78857),
            .in1(N__77933),
            .in2(N__75910),
            .in3(N__77171),
            .lcout(\PROM.ROMDATA.m349_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m357_am_LC_24_22_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m357_am_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m357_am_LC_24_22_6 .LUT_INIT=16'b1000111111011011;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m357_am_LC_24_22_6  (
            .in0(N__77173),
            .in1(N__75719),
            .in2(N__78036),
            .in3(N__78859),
            .lcout(),
            .ltout(\PROM.ROMDATA.m357_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m357_ns_LC_24_22_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m357_ns_LC_24_22_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m357_ns_LC_24_22_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m357_ns_LC_24_22_7  (
            .in0(_gnd_net_),
            .in1(N__74501),
            .in2(N__74495),
            .in3(N__76373),
            .lcout(\PROM.ROMDATA.m357_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m290_LC_24_23_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m290_LC_24_23_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m290_LC_24_23_0 .LUT_INIT=16'b0101000010001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m290_LC_24_23_0  (
            .in0(N__76533),
            .in1(N__74490),
            .in2(N__74411),
            .in3(N__75725),
            .lcout(),
            .ltout(\PROM.ROMDATA.m290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m303_ns_1_LC_24_23_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m303_ns_1_LC_24_23_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m303_ns_1_LC_24_23_1 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m303_ns_1_LC_24_23_1  (
            .in0(N__74378),
            .in1(N__79457),
            .in2(N__74363),
            .in3(N__79860),
            .lcout(\PROM.ROMDATA.m303_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m363_ns_LC_24_23_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m363_ns_LC_24_23_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m363_ns_LC_24_23_2 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m363_ns_LC_24_23_2  (
            .in0(N__79456),
            .in1(N__74348),
            .in2(N__74339),
            .in3(N__74291),
            .lcout(\PROM.ROMDATA.m363_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m353_am_LC_24_23_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m353_am_LC_24_23_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m353_am_LC_24_23_3 .LUT_INIT=16'b1000111111011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m353_am_LC_24_23_3  (
            .in0(N__78720),
            .in1(N__77892),
            .in2(N__75911),
            .in3(N__77240),
            .lcout(),
            .ltout(\PROM.ROMDATA.m353_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m353_ns_LC_24_23_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m353_ns_LC_24_23_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m353_ns_LC_24_23_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m353_ns_LC_24_23_4  (
            .in0(N__76532),
            .in1(_gnd_net_),
            .in2(N__74312),
            .in3(N__74309),
            .lcout(),
            .ltout(\PROM.ROMDATA.m353_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m363_ns_1_LC_24_23_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m363_ns_1_LC_24_23_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m363_ns_1_LC_24_23_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m363_ns_1_LC_24_23_5  (
            .in0(N__74936),
            .in1(N__79455),
            .in2(N__74294),
            .in3(N__79859),
            .lcout(\PROM.ROMDATA.m363_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m349_bm_LC_24_23_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m349_bm_LC_24_23_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m349_bm_LC_24_23_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m349_bm_LC_24_23_6  (
            .in0(N__74972),
            .in1(N__74962),
            .in2(_gnd_net_),
            .in3(N__75721),
            .lcout(),
            .ltout(\PROM.ROMDATA.m349_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m349_ns_LC_24_23_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m349_ns_LC_24_23_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m349_ns_LC_24_23_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m349_ns_LC_24_23_7  (
            .in0(_gnd_net_),
            .in1(N__74945),
            .in2(N__74939),
            .in3(N__76531),
            .lcout(\PROM.ROMDATA.m349_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m331_bm_LC_26_16_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m331_bm_LC_26_16_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m331_bm_LC_26_16_6 .LUT_INIT=16'b0000100100001000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m331_bm_LC_26_16_6  (
            .in0(N__78843),
            .in1(N__78011),
            .in2(N__76010),
            .in3(N__77309),
            .lcout(),
            .ltout(\PROM.ROMDATA.m331_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m331_ns_LC_26_16_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m331_ns_LC_26_16_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m331_ns_LC_26_16_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m331_ns_LC_26_16_7  (
            .in0(_gnd_net_),
            .in1(N__74507),
            .in2(N__74930),
            .in3(N__76617),
            .lcout(\PROM.ROMDATA.m331_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m323_am_LC_26_17_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m323_am_LC_26_17_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m323_am_LC_26_17_2 .LUT_INIT=16'b0010110000111000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m323_am_LC_26_17_2  (
            .in0(N__78841),
            .in1(N__78069),
            .in2(N__76016),
            .in3(N__77310),
            .lcout(),
            .ltout(\PROM.ROMDATA.m323_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m323_ns_LC_26_17_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m323_ns_LC_26_17_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m323_ns_LC_26_17_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m323_ns_LC_26_17_3  (
            .in0(_gnd_net_),
            .in1(N__74927),
            .in2(N__74915),
            .in3(N__76618),
            .lcout(\PROM.ROMDATA.m323_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFS1RP_15_LC_26_17_5 .C_ON=1'b0;
    defparam \ALU.c_RNIFS1RP_15_LC_26_17_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFS1RP_15_LC_26_17_5 .LUT_INIT=16'b0101010110111011;
    LogicCell40 \ALU.c_RNIFS1RP_15_LC_26_17_5  (
            .in0(N__74855),
            .in1(N__74618),
            .in2(_gnd_net_),
            .in3(N__74596),
            .lcout(\ALU.N_586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m331_am_LC_26_17_6 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m331_am_LC_26_17_6 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m331_am_LC_26_17_6 .LUT_INIT=16'b0010000010101000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m331_am_LC_26_17_6  (
            .in0(N__76011),
            .in1(N__78840),
            .in2(N__79049),
            .in3(N__78068),
            .lcout(\PROM.ROMDATA.m331_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m341_ns_1_LC_26_18_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m341_ns_1_LC_26_18_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m341_ns_1_LC_26_18_3 .LUT_INIT=16'b0000011100111110;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m341_ns_1_LC_26_18_3  (
            .in0(N__78637),
            .in1(N__78067),
            .in2(N__76008),
            .in3(N__77318),
            .lcout(\PROM.ROMDATA.m341_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m343_ns_1_LC_26_19_0 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m343_ns_1_LC_26_19_0 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m343_ns_1_LC_26_19_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m343_ns_1_LC_26_19_0  (
            .in0(N__79907),
            .in1(N__79415),
            .in2(N__78872),
            .in3(N__79883),
            .lcout(),
            .ltout(\PROM.ROMDATA.m343_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m343_ns_LC_26_19_1 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m343_ns_LC_26_19_1 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m343_ns_LC_26_19_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m343_ns_LC_26_19_1  (
            .in0(N__79416),
            .in1(N__74978),
            .in2(N__79067),
            .in3(N__76661),
            .lcout(\PROM.ROMDATA.m343_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m334_ns_1_LC_26_19_2 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m334_ns_1_LC_26_19_2 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m334_ns_1_LC_26_19_2 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m334_ns_1_LC_26_19_2  (
            .in0(N__76569),
            .in1(N__79044),
            .in2(_gnd_net_),
            .in3(N__78998),
            .lcout(),
            .ltout(\PROM.ROMDATA.m334_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m334_ns_LC_26_19_3 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m334_ns_LC_26_19_3 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m334_ns_LC_26_19_3 .LUT_INIT=16'b1101000100000000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m334_ns_LC_26_19_3  (
            .in0(N__78061),
            .in1(N__78887),
            .in2(N__78875),
            .in3(N__78778),
            .lcout(\PROM.ROMDATA.i3_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m338_am_LC_26_19_4 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m338_am_LC_26_19_4 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m338_am_LC_26_19_4 .LUT_INIT=16'b0100011110001100;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m338_am_LC_26_19_4  (
            .in0(N__78777),
            .in1(N__78062),
            .in2(N__76009),
            .in3(N__77311),
            .lcout(),
            .ltout(\PROM.ROMDATA.m338_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m338_ns_LC_26_19_5 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m338_ns_LC_26_19_5 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m338_ns_LC_26_19_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m338_ns_LC_26_19_5  (
            .in0(_gnd_net_),
            .in1(N__76679),
            .in2(N__76664),
            .in3(N__76571),
            .lcout(\PROM.ROMDATA.m338_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PROM.ROMDATA.dintern_31_0__m341_ns_LC_26_19_7 .C_ON=1'b0;
    defparam \PROM.ROMDATA.dintern_31_0__m341_ns_LC_26_19_7 .SEQ_MODE=4'b0000;
    defparam \PROM.ROMDATA.dintern_31_0__m341_ns_LC_26_19_7 .LUT_INIT=16'b0011000011010001;
    LogicCell40 \PROM.ROMDATA.dintern_31_0__m341_ns_LC_26_19_7  (
            .in0(N__76655),
            .in1(N__76570),
            .in2(N__76028),
            .in3(N__75983),
            .lcout(\PROM.ROMDATA.m341_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
