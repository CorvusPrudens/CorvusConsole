-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 27 2020 03:05:38

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    BUFFER_DATA_OUT : out std_logic_vector(15 downto 0);
    BUFFER_DATA_IN : in std_logic_vector(15 downto 0);
    BUFFER_ADDRESS : out std_logic_vector(15 downto 0);
    A13 : out std_logic;
    D6_in : in std_logic;
    A9 : out std_logic;
    D3 : out std_logic;
    CLK : in std_logic;
    A6 : out std_logic;
    RX : in std_logic;
    D8_in : in std_logic;
    D7 : out std_logic;
    D12 : out std_logic;
    CE : out std_logic;
    D9_in : in std_logic;
    D5_in : in std_logic;
    D0_in : in std_logic;
    B_OE : out std_logic;
    A10 : out std_logic;
    D10_in : in std_logic;
    A8 : out std_logic;
    D11_in : in std_logic;
    D0 : out std_logic;
    A1 : out std_logic;
    GPIO11 : out std_logic;
    D4_in : in std_logic;
    GPIO9 : out std_logic;
    A14 : out std_logic;
    LB : out std_logic;
    D4 : out std_logic;
    D13_in : in std_logic;
    D11 : out std_logic;
    B_CE : out std_logic;
    A5 : out std_logic;
    D14_in : in std_logic;
    B_WR : out std_logic;
    A2 : out std_logic;
    A11 : out std_logic;
    D6 : out std_logic;
    D13 : out std_logic;
    B_LB : out std_logic;
    D1 : out std_logic;
    A0 : out std_logic;
    OE : out std_logic;
    D8 : out std_logic;
    D15 : out std_logic;
    D15_in : in std_logic;
    A15 : out std_logic;
    UB : out std_logic;
    D5 : out std_logic;
    D10 : out std_logic;
    A4 : out std_logic;
    GPIO3 : out std_logic;
    D1_in : in std_logic;
    TX : out std_logic;
    D7_in : in std_logic;
    A3 : out std_logic;
    D9 : out std_logic;
    D14 : out std_logic;
    WR : out std_logic;
    D3_in : in std_logic;
    A12 : out std_logic;
    D2_in : in std_logic;
    D12_in : in std_logic;
    D2 : out std_logic;
    B_UB : out std_logic;
    A7 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__80918\ : std_logic;
signal \N__80917\ : std_logic;
signal \N__80916\ : std_logic;
signal \N__80907\ : std_logic;
signal \N__80906\ : std_logic;
signal \N__80905\ : std_logic;
signal \N__80898\ : std_logic;
signal \N__80897\ : std_logic;
signal \N__80896\ : std_logic;
signal \N__80889\ : std_logic;
signal \N__80888\ : std_logic;
signal \N__80887\ : std_logic;
signal \N__80880\ : std_logic;
signal \N__80879\ : std_logic;
signal \N__80878\ : std_logic;
signal \N__80871\ : std_logic;
signal \N__80870\ : std_logic;
signal \N__80869\ : std_logic;
signal \N__80862\ : std_logic;
signal \N__80861\ : std_logic;
signal \N__80860\ : std_logic;
signal \N__80853\ : std_logic;
signal \N__80852\ : std_logic;
signal \N__80851\ : std_logic;
signal \N__80844\ : std_logic;
signal \N__80843\ : std_logic;
signal \N__80842\ : std_logic;
signal \N__80835\ : std_logic;
signal \N__80834\ : std_logic;
signal \N__80833\ : std_logic;
signal \N__80826\ : std_logic;
signal \N__80825\ : std_logic;
signal \N__80824\ : std_logic;
signal \N__80817\ : std_logic;
signal \N__80816\ : std_logic;
signal \N__80815\ : std_logic;
signal \N__80808\ : std_logic;
signal \N__80807\ : std_logic;
signal \N__80806\ : std_logic;
signal \N__80799\ : std_logic;
signal \N__80798\ : std_logic;
signal \N__80797\ : std_logic;
signal \N__80790\ : std_logic;
signal \N__80789\ : std_logic;
signal \N__80788\ : std_logic;
signal \N__80781\ : std_logic;
signal \N__80780\ : std_logic;
signal \N__80779\ : std_logic;
signal \N__80772\ : std_logic;
signal \N__80771\ : std_logic;
signal \N__80770\ : std_logic;
signal \N__80763\ : std_logic;
signal \N__80762\ : std_logic;
signal \N__80761\ : std_logic;
signal \N__80754\ : std_logic;
signal \N__80753\ : std_logic;
signal \N__80752\ : std_logic;
signal \N__80745\ : std_logic;
signal \N__80744\ : std_logic;
signal \N__80743\ : std_logic;
signal \N__80736\ : std_logic;
signal \N__80735\ : std_logic;
signal \N__80734\ : std_logic;
signal \N__80727\ : std_logic;
signal \N__80726\ : std_logic;
signal \N__80725\ : std_logic;
signal \N__80718\ : std_logic;
signal \N__80717\ : std_logic;
signal \N__80716\ : std_logic;
signal \N__80709\ : std_logic;
signal \N__80708\ : std_logic;
signal \N__80707\ : std_logic;
signal \N__80700\ : std_logic;
signal \N__80699\ : std_logic;
signal \N__80698\ : std_logic;
signal \N__80691\ : std_logic;
signal \N__80690\ : std_logic;
signal \N__80689\ : std_logic;
signal \N__80682\ : std_logic;
signal \N__80681\ : std_logic;
signal \N__80680\ : std_logic;
signal \N__80673\ : std_logic;
signal \N__80672\ : std_logic;
signal \N__80671\ : std_logic;
signal \N__80664\ : std_logic;
signal \N__80663\ : std_logic;
signal \N__80662\ : std_logic;
signal \N__80655\ : std_logic;
signal \N__80654\ : std_logic;
signal \N__80653\ : std_logic;
signal \N__80646\ : std_logic;
signal \N__80645\ : std_logic;
signal \N__80644\ : std_logic;
signal \N__80637\ : std_logic;
signal \N__80636\ : std_logic;
signal \N__80635\ : std_logic;
signal \N__80628\ : std_logic;
signal \N__80627\ : std_logic;
signal \N__80626\ : std_logic;
signal \N__80619\ : std_logic;
signal \N__80618\ : std_logic;
signal \N__80617\ : std_logic;
signal \N__80610\ : std_logic;
signal \N__80609\ : std_logic;
signal \N__80608\ : std_logic;
signal \N__80601\ : std_logic;
signal \N__80600\ : std_logic;
signal \N__80599\ : std_logic;
signal \N__80592\ : std_logic;
signal \N__80591\ : std_logic;
signal \N__80590\ : std_logic;
signal \N__80583\ : std_logic;
signal \N__80582\ : std_logic;
signal \N__80581\ : std_logic;
signal \N__80574\ : std_logic;
signal \N__80573\ : std_logic;
signal \N__80572\ : std_logic;
signal \N__80565\ : std_logic;
signal \N__80564\ : std_logic;
signal \N__80563\ : std_logic;
signal \N__80556\ : std_logic;
signal \N__80555\ : std_logic;
signal \N__80554\ : std_logic;
signal \N__80547\ : std_logic;
signal \N__80546\ : std_logic;
signal \N__80545\ : std_logic;
signal \N__80538\ : std_logic;
signal \N__80537\ : std_logic;
signal \N__80536\ : std_logic;
signal \N__80529\ : std_logic;
signal \N__80528\ : std_logic;
signal \N__80527\ : std_logic;
signal \N__80520\ : std_logic;
signal \N__80519\ : std_logic;
signal \N__80518\ : std_logic;
signal \N__80511\ : std_logic;
signal \N__80510\ : std_logic;
signal \N__80509\ : std_logic;
signal \N__80502\ : std_logic;
signal \N__80501\ : std_logic;
signal \N__80500\ : std_logic;
signal \N__80493\ : std_logic;
signal \N__80492\ : std_logic;
signal \N__80491\ : std_logic;
signal \N__80484\ : std_logic;
signal \N__80483\ : std_logic;
signal \N__80482\ : std_logic;
signal \N__80475\ : std_logic;
signal \N__80474\ : std_logic;
signal \N__80473\ : std_logic;
signal \N__80466\ : std_logic;
signal \N__80465\ : std_logic;
signal \N__80464\ : std_logic;
signal \N__80457\ : std_logic;
signal \N__80456\ : std_logic;
signal \N__80455\ : std_logic;
signal \N__80448\ : std_logic;
signal \N__80447\ : std_logic;
signal \N__80446\ : std_logic;
signal \N__80439\ : std_logic;
signal \N__80438\ : std_logic;
signal \N__80437\ : std_logic;
signal \N__80430\ : std_logic;
signal \N__80429\ : std_logic;
signal \N__80428\ : std_logic;
signal \N__80421\ : std_logic;
signal \N__80420\ : std_logic;
signal \N__80419\ : std_logic;
signal \N__80412\ : std_logic;
signal \N__80411\ : std_logic;
signal \N__80410\ : std_logic;
signal \N__80403\ : std_logic;
signal \N__80402\ : std_logic;
signal \N__80401\ : std_logic;
signal \N__80394\ : std_logic;
signal \N__80393\ : std_logic;
signal \N__80392\ : std_logic;
signal \N__80385\ : std_logic;
signal \N__80384\ : std_logic;
signal \N__80383\ : std_logic;
signal \N__80376\ : std_logic;
signal \N__80375\ : std_logic;
signal \N__80374\ : std_logic;
signal \N__80367\ : std_logic;
signal \N__80366\ : std_logic;
signal \N__80365\ : std_logic;
signal \N__80358\ : std_logic;
signal \N__80357\ : std_logic;
signal \N__80356\ : std_logic;
signal \N__80349\ : std_logic;
signal \N__80348\ : std_logic;
signal \N__80347\ : std_logic;
signal \N__80340\ : std_logic;
signal \N__80339\ : std_logic;
signal \N__80338\ : std_logic;
signal \N__80331\ : std_logic;
signal \N__80330\ : std_logic;
signal \N__80329\ : std_logic;
signal \N__80322\ : std_logic;
signal \N__80321\ : std_logic;
signal \N__80320\ : std_logic;
signal \N__80313\ : std_logic;
signal \N__80312\ : std_logic;
signal \N__80311\ : std_logic;
signal \N__80304\ : std_logic;
signal \N__80303\ : std_logic;
signal \N__80302\ : std_logic;
signal \N__80295\ : std_logic;
signal \N__80294\ : std_logic;
signal \N__80293\ : std_logic;
signal \N__80286\ : std_logic;
signal \N__80285\ : std_logic;
signal \N__80284\ : std_logic;
signal \N__80277\ : std_logic;
signal \N__80276\ : std_logic;
signal \N__80275\ : std_logic;
signal \N__80268\ : std_logic;
signal \N__80267\ : std_logic;
signal \N__80266\ : std_logic;
signal \N__80259\ : std_logic;
signal \N__80258\ : std_logic;
signal \N__80257\ : std_logic;
signal \N__80250\ : std_logic;
signal \N__80249\ : std_logic;
signal \N__80248\ : std_logic;
signal \N__80241\ : std_logic;
signal \N__80240\ : std_logic;
signal \N__80239\ : std_logic;
signal \N__80232\ : std_logic;
signal \N__80231\ : std_logic;
signal \N__80230\ : std_logic;
signal \N__80223\ : std_logic;
signal \N__80222\ : std_logic;
signal \N__80221\ : std_logic;
signal \N__80214\ : std_logic;
signal \N__80213\ : std_logic;
signal \N__80212\ : std_logic;
signal \N__80205\ : std_logic;
signal \N__80204\ : std_logic;
signal \N__80203\ : std_logic;
signal \N__80196\ : std_logic;
signal \N__80195\ : std_logic;
signal \N__80194\ : std_logic;
signal \N__80187\ : std_logic;
signal \N__80186\ : std_logic;
signal \N__80185\ : std_logic;
signal \N__80178\ : std_logic;
signal \N__80177\ : std_logic;
signal \N__80176\ : std_logic;
signal \N__80169\ : std_logic;
signal \N__80168\ : std_logic;
signal \N__80167\ : std_logic;
signal \N__80160\ : std_logic;
signal \N__80159\ : std_logic;
signal \N__80158\ : std_logic;
signal \N__80151\ : std_logic;
signal \N__80150\ : std_logic;
signal \N__80149\ : std_logic;
signal \N__80142\ : std_logic;
signal \N__80141\ : std_logic;
signal \N__80140\ : std_logic;
signal \N__80133\ : std_logic;
signal \N__80132\ : std_logic;
signal \N__80131\ : std_logic;
signal \N__80124\ : std_logic;
signal \N__80123\ : std_logic;
signal \N__80122\ : std_logic;
signal \N__80115\ : std_logic;
signal \N__80114\ : std_logic;
signal \N__80113\ : std_logic;
signal \N__80106\ : std_logic;
signal \N__80105\ : std_logic;
signal \N__80104\ : std_logic;
signal \N__80097\ : std_logic;
signal \N__80096\ : std_logic;
signal \N__80095\ : std_logic;
signal \N__80088\ : std_logic;
signal \N__80087\ : std_logic;
signal \N__80086\ : std_logic;
signal \N__80079\ : std_logic;
signal \N__80078\ : std_logic;
signal \N__80077\ : std_logic;
signal \N__80070\ : std_logic;
signal \N__80069\ : std_logic;
signal \N__80068\ : std_logic;
signal \N__80061\ : std_logic;
signal \N__80060\ : std_logic;
signal \N__80059\ : std_logic;
signal \N__80052\ : std_logic;
signal \N__80051\ : std_logic;
signal \N__80050\ : std_logic;
signal \N__80043\ : std_logic;
signal \N__80042\ : std_logic;
signal \N__80041\ : std_logic;
signal \N__80034\ : std_logic;
signal \N__80033\ : std_logic;
signal \N__80032\ : std_logic;
signal \N__80025\ : std_logic;
signal \N__80024\ : std_logic;
signal \N__80023\ : std_logic;
signal \N__80016\ : std_logic;
signal \N__80015\ : std_logic;
signal \N__80014\ : std_logic;
signal \N__80007\ : std_logic;
signal \N__80006\ : std_logic;
signal \N__80005\ : std_logic;
signal \N__79998\ : std_logic;
signal \N__79997\ : std_logic;
signal \N__79996\ : std_logic;
signal \N__79989\ : std_logic;
signal \N__79988\ : std_logic;
signal \N__79987\ : std_logic;
signal \N__79980\ : std_logic;
signal \N__79979\ : std_logic;
signal \N__79978\ : std_logic;
signal \N__79971\ : std_logic;
signal \N__79970\ : std_logic;
signal \N__79969\ : std_logic;
signal \N__79962\ : std_logic;
signal \N__79961\ : std_logic;
signal \N__79960\ : std_logic;
signal \N__79953\ : std_logic;
signal \N__79952\ : std_logic;
signal \N__79951\ : std_logic;
signal \N__79944\ : std_logic;
signal \N__79943\ : std_logic;
signal \N__79942\ : std_logic;
signal \N__79935\ : std_logic;
signal \N__79934\ : std_logic;
signal \N__79933\ : std_logic;
signal \N__79926\ : std_logic;
signal \N__79925\ : std_logic;
signal \N__79924\ : std_logic;
signal \N__79907\ : std_logic;
signal \N__79904\ : std_logic;
signal \N__79901\ : std_logic;
signal \N__79898\ : std_logic;
signal \N__79897\ : std_logic;
signal \N__79896\ : std_logic;
signal \N__79895\ : std_logic;
signal \N__79892\ : std_logic;
signal \N__79891\ : std_logic;
signal \N__79890\ : std_logic;
signal \N__79887\ : std_logic;
signal \N__79884\ : std_logic;
signal \N__79883\ : std_logic;
signal \N__79882\ : std_logic;
signal \N__79881\ : std_logic;
signal \N__79880\ : std_logic;
signal \N__79879\ : std_logic;
signal \N__79878\ : std_logic;
signal \N__79875\ : std_logic;
signal \N__79874\ : std_logic;
signal \N__79873\ : std_logic;
signal \N__79872\ : std_logic;
signal \N__79871\ : std_logic;
signal \N__79870\ : std_logic;
signal \N__79867\ : std_logic;
signal \N__79866\ : std_logic;
signal \N__79863\ : std_logic;
signal \N__79862\ : std_logic;
signal \N__79861\ : std_logic;
signal \N__79860\ : std_logic;
signal \N__79859\ : std_logic;
signal \N__79858\ : std_logic;
signal \N__79857\ : std_logic;
signal \N__79854\ : std_logic;
signal \N__79851\ : std_logic;
signal \N__79850\ : std_logic;
signal \N__79847\ : std_logic;
signal \N__79846\ : std_logic;
signal \N__79845\ : std_logic;
signal \N__79844\ : std_logic;
signal \N__79843\ : std_logic;
signal \N__79842\ : std_logic;
signal \N__79841\ : std_logic;
signal \N__79840\ : std_logic;
signal \N__79839\ : std_logic;
signal \N__79838\ : std_logic;
signal \N__79835\ : std_logic;
signal \N__79834\ : std_logic;
signal \N__79833\ : std_logic;
signal \N__79832\ : std_logic;
signal \N__79831\ : std_logic;
signal \N__79830\ : std_logic;
signal \N__79819\ : std_logic;
signal \N__79818\ : std_logic;
signal \N__79815\ : std_logic;
signal \N__79812\ : std_logic;
signal \N__79809\ : std_logic;
signal \N__79808\ : std_logic;
signal \N__79801\ : std_logic;
signal \N__79798\ : std_logic;
signal \N__79795\ : std_logic;
signal \N__79792\ : std_logic;
signal \N__79789\ : std_logic;
signal \N__79788\ : std_logic;
signal \N__79787\ : std_logic;
signal \N__79784\ : std_logic;
signal \N__79783\ : std_logic;
signal \N__79778\ : std_logic;
signal \N__79775\ : std_logic;
signal \N__79772\ : std_logic;
signal \N__79769\ : std_logic;
signal \N__79766\ : std_logic;
signal \N__79763\ : std_logic;
signal \N__79762\ : std_logic;
signal \N__79761\ : std_logic;
signal \N__79758\ : std_logic;
signal \N__79755\ : std_logic;
signal \N__79752\ : std_logic;
signal \N__79751\ : std_logic;
signal \N__79748\ : std_logic;
signal \N__79747\ : std_logic;
signal \N__79744\ : std_logic;
signal \N__79741\ : std_logic;
signal \N__79738\ : std_logic;
signal \N__79735\ : std_logic;
signal \N__79732\ : std_logic;
signal \N__79729\ : std_logic;
signal \N__79726\ : std_logic;
signal \N__79723\ : std_logic;
signal \N__79716\ : std_logic;
signal \N__79715\ : std_logic;
signal \N__79714\ : std_logic;
signal \N__79711\ : std_logic;
signal \N__79708\ : std_logic;
signal \N__79705\ : std_logic;
signal \N__79698\ : std_logic;
signal \N__79695\ : std_logic;
signal \N__79692\ : std_logic;
signal \N__79683\ : std_logic;
signal \N__79678\ : std_logic;
signal \N__79675\ : std_logic;
signal \N__79672\ : std_logic;
signal \N__79667\ : std_logic;
signal \N__79662\ : std_logic;
signal \N__79657\ : std_logic;
signal \N__79652\ : std_logic;
signal \N__79649\ : std_logic;
signal \N__79644\ : std_logic;
signal \N__79641\ : std_logic;
signal \N__79638\ : std_logic;
signal \N__79635\ : std_logic;
signal \N__79628\ : std_logic;
signal \N__79621\ : std_logic;
signal \N__79614\ : std_logic;
signal \N__79613\ : std_logic;
signal \N__79610\ : std_logic;
signal \N__79605\ : std_logic;
signal \N__79598\ : std_logic;
signal \N__79591\ : std_logic;
signal \N__79584\ : std_logic;
signal \N__79581\ : std_logic;
signal \N__79578\ : std_logic;
signal \N__79573\ : std_logic;
signal \N__79556\ : std_logic;
signal \N__79553\ : std_logic;
signal \N__79532\ : std_logic;
signal \N__79531\ : std_logic;
signal \N__79530\ : std_logic;
signal \N__79529\ : std_logic;
signal \N__79528\ : std_logic;
signal \N__79527\ : std_logic;
signal \N__79524\ : std_logic;
signal \N__79523\ : std_logic;
signal \N__79522\ : std_logic;
signal \N__79519\ : std_logic;
signal \N__79516\ : std_logic;
signal \N__79515\ : std_logic;
signal \N__79514\ : std_logic;
signal \N__79511\ : std_logic;
signal \N__79508\ : std_logic;
signal \N__79507\ : std_logic;
signal \N__79504\ : std_logic;
signal \N__79503\ : std_logic;
signal \N__79502\ : std_logic;
signal \N__79501\ : std_logic;
signal \N__79500\ : std_logic;
signal \N__79499\ : std_logic;
signal \N__79498\ : std_logic;
signal \N__79497\ : std_logic;
signal \N__79496\ : std_logic;
signal \N__79495\ : std_logic;
signal \N__79490\ : std_logic;
signal \N__79489\ : std_logic;
signal \N__79488\ : std_logic;
signal \N__79487\ : std_logic;
signal \N__79486\ : std_logic;
signal \N__79483\ : std_logic;
signal \N__79474\ : std_logic;
signal \N__79469\ : std_logic;
signal \N__79464\ : std_logic;
signal \N__79461\ : std_logic;
signal \N__79458\ : std_logic;
signal \N__79457\ : std_logic;
signal \N__79456\ : std_logic;
signal \N__79455\ : std_logic;
signal \N__79454\ : std_logic;
signal \N__79453\ : std_logic;
signal \N__79452\ : std_logic;
signal \N__79447\ : std_logic;
signal \N__79440\ : std_logic;
signal \N__79437\ : std_logic;
signal \N__79434\ : std_logic;
signal \N__79433\ : std_logic;
signal \N__79432\ : std_logic;
signal \N__79431\ : std_logic;
signal \N__79428\ : std_logic;
signal \N__79425\ : std_logic;
signal \N__79422\ : std_logic;
signal \N__79421\ : std_logic;
signal \N__79420\ : std_logic;
signal \N__79419\ : std_logic;
signal \N__79418\ : std_logic;
signal \N__79417\ : std_logic;
signal \N__79416\ : std_logic;
signal \N__79415\ : std_logic;
signal \N__79414\ : std_logic;
signal \N__79413\ : std_logic;
signal \N__79412\ : std_logic;
signal \N__79411\ : std_logic;
signal \N__79408\ : std_logic;
signal \N__79405\ : std_logic;
signal \N__79398\ : std_logic;
signal \N__79395\ : std_logic;
signal \N__79392\ : std_logic;
signal \N__79391\ : std_logic;
signal \N__79388\ : std_logic;
signal \N__79381\ : std_logic;
signal \N__79378\ : std_logic;
signal \N__79373\ : std_logic;
signal \N__79370\ : std_logic;
signal \N__79367\ : std_logic;
signal \N__79358\ : std_logic;
signal \N__79355\ : std_logic;
signal \N__79352\ : std_logic;
signal \N__79343\ : std_logic;
signal \N__79342\ : std_logic;
signal \N__79341\ : std_logic;
signal \N__79336\ : std_logic;
signal \N__79333\ : std_logic;
signal \N__79328\ : std_logic;
signal \N__79327\ : std_logic;
signal \N__79324\ : std_logic;
signal \N__79323\ : std_logic;
signal \N__79322\ : std_logic;
signal \N__79321\ : std_logic;
signal \N__79320\ : std_logic;
signal \N__79319\ : std_logic;
signal \N__79318\ : std_logic;
signal \N__79315\ : std_logic;
signal \N__79314\ : std_logic;
signal \N__79309\ : std_logic;
signal \N__79306\ : std_logic;
signal \N__79301\ : std_logic;
signal \N__79300\ : std_logic;
signal \N__79299\ : std_logic;
signal \N__79298\ : std_logic;
signal \N__79297\ : std_logic;
signal \N__79294\ : std_logic;
signal \N__79293\ : std_logic;
signal \N__79290\ : std_logic;
signal \N__79287\ : std_logic;
signal \N__79286\ : std_logic;
signal \N__79277\ : std_logic;
signal \N__79274\ : std_logic;
signal \N__79269\ : std_logic;
signal \N__79262\ : std_logic;
signal \N__79259\ : std_logic;
signal \N__79256\ : std_logic;
signal \N__79253\ : std_logic;
signal \N__79250\ : std_logic;
signal \N__79249\ : std_logic;
signal \N__79248\ : std_logic;
signal \N__79245\ : std_logic;
signal \N__79238\ : std_logic;
signal \N__79233\ : std_logic;
signal \N__79228\ : std_logic;
signal \N__79223\ : std_logic;
signal \N__79220\ : std_logic;
signal \N__79217\ : std_logic;
signal \N__79214\ : std_logic;
signal \N__79211\ : std_logic;
signal \N__79210\ : std_logic;
signal \N__79209\ : std_logic;
signal \N__79208\ : std_logic;
signal \N__79207\ : std_logic;
signal \N__79204\ : std_logic;
signal \N__79201\ : std_logic;
signal \N__79196\ : std_logic;
signal \N__79193\ : std_logic;
signal \N__79190\ : std_logic;
signal \N__79185\ : std_logic;
signal \N__79182\ : std_logic;
signal \N__79179\ : std_logic;
signal \N__79176\ : std_logic;
signal \N__79171\ : std_logic;
signal \N__79162\ : std_logic;
signal \N__79157\ : std_logic;
signal \N__79150\ : std_logic;
signal \N__79143\ : std_logic;
signal \N__79142\ : std_logic;
signal \N__79139\ : std_logic;
signal \N__79134\ : std_logic;
signal \N__79131\ : std_logic;
signal \N__79126\ : std_logic;
signal \N__79123\ : std_logic;
signal \N__79116\ : std_logic;
signal \N__79111\ : std_logic;
signal \N__79104\ : std_logic;
signal \N__79091\ : std_logic;
signal \N__79088\ : std_logic;
signal \N__79067\ : std_logic;
signal \N__79064\ : std_logic;
signal \N__79061\ : std_logic;
signal \N__79058\ : std_logic;
signal \N__79055\ : std_logic;
signal \N__79052\ : std_logic;
signal \N__79049\ : std_logic;
signal \N__79048\ : std_logic;
signal \N__79045\ : std_logic;
signal \N__79044\ : std_logic;
signal \N__79043\ : std_logic;
signal \N__79040\ : std_logic;
signal \N__79037\ : std_logic;
signal \N__79034\ : std_logic;
signal \N__79033\ : std_logic;
signal \N__79030\ : std_logic;
signal \N__79027\ : std_logic;
signal \N__79024\ : std_logic;
signal \N__79021\ : std_logic;
signal \N__79016\ : std_logic;
signal \N__79011\ : std_logic;
signal \N__79006\ : std_logic;
signal \N__79001\ : std_logic;
signal \N__78998\ : std_logic;
signal \N__78997\ : std_logic;
signal \N__78996\ : std_logic;
signal \N__78995\ : std_logic;
signal \N__78994\ : std_logic;
signal \N__78993\ : std_logic;
signal \N__78990\ : std_logic;
signal \N__78989\ : std_logic;
signal \N__78988\ : std_logic;
signal \N__78985\ : std_logic;
signal \N__78984\ : std_logic;
signal \N__78981\ : std_logic;
signal \N__78980\ : std_logic;
signal \N__78977\ : std_logic;
signal \N__78972\ : std_logic;
signal \N__78969\ : std_logic;
signal \N__78966\ : std_logic;
signal \N__78963\ : std_logic;
signal \N__78960\ : std_logic;
signal \N__78957\ : std_logic;
signal \N__78956\ : std_logic;
signal \N__78955\ : std_logic;
signal \N__78952\ : std_logic;
signal \N__78949\ : std_logic;
signal \N__78944\ : std_logic;
signal \N__78943\ : std_logic;
signal \N__78940\ : std_logic;
signal \N__78937\ : std_logic;
signal \N__78934\ : std_logic;
signal \N__78929\ : std_logic;
signal \N__78924\ : std_logic;
signal \N__78921\ : std_logic;
signal \N__78918\ : std_logic;
signal \N__78915\ : std_logic;
signal \N__78912\ : std_logic;
signal \N__78905\ : std_logic;
signal \N__78900\ : std_logic;
signal \N__78887\ : std_logic;
signal \N__78884\ : std_logic;
signal \N__78881\ : std_logic;
signal \N__78878\ : std_logic;
signal \N__78875\ : std_logic;
signal \N__78872\ : std_logic;
signal \N__78869\ : std_logic;
signal \N__78866\ : std_logic;
signal \N__78863\ : std_logic;
signal \N__78862\ : std_logic;
signal \N__78861\ : std_logic;
signal \N__78860\ : std_logic;
signal \N__78859\ : std_logic;
signal \N__78858\ : std_logic;
signal \N__78857\ : std_logic;
signal \N__78856\ : std_logic;
signal \N__78855\ : std_logic;
signal \N__78854\ : std_logic;
signal \N__78853\ : std_logic;
signal \N__78852\ : std_logic;
signal \N__78851\ : std_logic;
signal \N__78850\ : std_logic;
signal \N__78849\ : std_logic;
signal \N__78846\ : std_logic;
signal \N__78845\ : std_logic;
signal \N__78844\ : std_logic;
signal \N__78843\ : std_logic;
signal \N__78842\ : std_logic;
signal \N__78841\ : std_logic;
signal \N__78840\ : std_logic;
signal \N__78839\ : std_logic;
signal \N__78838\ : std_logic;
signal \N__78837\ : std_logic;
signal \N__78836\ : std_logic;
signal \N__78835\ : std_logic;
signal \N__78834\ : std_logic;
signal \N__78833\ : std_logic;
signal \N__78832\ : std_logic;
signal \N__78831\ : std_logic;
signal \N__78830\ : std_logic;
signal \N__78829\ : std_logic;
signal \N__78828\ : std_logic;
signal \N__78827\ : std_logic;
signal \N__78824\ : std_logic;
signal \N__78823\ : std_logic;
signal \N__78820\ : std_logic;
signal \N__78819\ : std_logic;
signal \N__78818\ : std_logic;
signal \N__78815\ : std_logic;
signal \N__78814\ : std_logic;
signal \N__78813\ : std_logic;
signal \N__78812\ : std_logic;
signal \N__78811\ : std_logic;
signal \N__78810\ : std_logic;
signal \N__78809\ : std_logic;
signal \N__78808\ : std_logic;
signal \N__78807\ : std_logic;
signal \N__78806\ : std_logic;
signal \N__78799\ : std_logic;
signal \N__78798\ : std_logic;
signal \N__78797\ : std_logic;
signal \N__78796\ : std_logic;
signal \N__78795\ : std_logic;
signal \N__78794\ : std_logic;
signal \N__78793\ : std_logic;
signal \N__78792\ : std_logic;
signal \N__78791\ : std_logic;
signal \N__78790\ : std_logic;
signal \N__78789\ : std_logic;
signal \N__78788\ : std_logic;
signal \N__78787\ : std_logic;
signal \N__78780\ : std_logic;
signal \N__78779\ : std_logic;
signal \N__78778\ : std_logic;
signal \N__78777\ : std_logic;
signal \N__78776\ : std_logic;
signal \N__78775\ : std_logic;
signal \N__78774\ : std_logic;
signal \N__78773\ : std_logic;
signal \N__78770\ : std_logic;
signal \N__78769\ : std_logic;
signal \N__78768\ : std_logic;
signal \N__78767\ : std_logic;
signal \N__78766\ : std_logic;
signal \N__78761\ : std_logic;
signal \N__78754\ : std_logic;
signal \N__78753\ : std_logic;
signal \N__78750\ : std_logic;
signal \N__78747\ : std_logic;
signal \N__78746\ : std_logic;
signal \N__78745\ : std_logic;
signal \N__78744\ : std_logic;
signal \N__78741\ : std_logic;
signal \N__78738\ : std_logic;
signal \N__78737\ : std_logic;
signal \N__78736\ : std_logic;
signal \N__78735\ : std_logic;
signal \N__78734\ : std_logic;
signal \N__78733\ : std_logic;
signal \N__78732\ : std_logic;
signal \N__78731\ : std_logic;
signal \N__78730\ : std_logic;
signal \N__78729\ : std_logic;
signal \N__78728\ : std_logic;
signal \N__78727\ : std_logic;
signal \N__78724\ : std_logic;
signal \N__78721\ : std_logic;
signal \N__78720\ : std_logic;
signal \N__78719\ : std_logic;
signal \N__78718\ : std_logic;
signal \N__78715\ : std_logic;
signal \N__78714\ : std_logic;
signal \N__78713\ : std_logic;
signal \N__78712\ : std_logic;
signal \N__78705\ : std_logic;
signal \N__78704\ : std_logic;
signal \N__78701\ : std_logic;
signal \N__78700\ : std_logic;
signal \N__78697\ : std_logic;
signal \N__78696\ : std_logic;
signal \N__78695\ : std_logic;
signal \N__78694\ : std_logic;
signal \N__78693\ : std_logic;
signal \N__78692\ : std_logic;
signal \N__78689\ : std_logic;
signal \N__78688\ : std_logic;
signal \N__78687\ : std_logic;
signal \N__78686\ : std_logic;
signal \N__78685\ : std_logic;
signal \N__78680\ : std_logic;
signal \N__78679\ : std_logic;
signal \N__78678\ : std_logic;
signal \N__78677\ : std_logic;
signal \N__78672\ : std_logic;
signal \N__78663\ : std_logic;
signal \N__78652\ : std_logic;
signal \N__78641\ : std_logic;
signal \N__78640\ : std_logic;
signal \N__78639\ : std_logic;
signal \N__78638\ : std_logic;
signal \N__78637\ : std_logic;
signal \N__78636\ : std_logic;
signal \N__78635\ : std_logic;
signal \N__78634\ : std_logic;
signal \N__78631\ : std_logic;
signal \N__78626\ : std_logic;
signal \N__78625\ : std_logic;
signal \N__78622\ : std_logic;
signal \N__78613\ : std_logic;
signal \N__78606\ : std_logic;
signal \N__78597\ : std_logic;
signal \N__78594\ : std_logic;
signal \N__78591\ : std_logic;
signal \N__78588\ : std_logic;
signal \N__78583\ : std_logic;
signal \N__78574\ : std_logic;
signal \N__78573\ : std_logic;
signal \N__78570\ : std_logic;
signal \N__78569\ : std_logic;
signal \N__78560\ : std_logic;
signal \N__78555\ : std_logic;
signal \N__78552\ : std_logic;
signal \N__78547\ : std_logic;
signal \N__78544\ : std_logic;
signal \N__78543\ : std_logic;
signal \N__78542\ : std_logic;
signal \N__78537\ : std_logic;
signal \N__78532\ : std_logic;
signal \N__78523\ : std_logic;
signal \N__78516\ : std_logic;
signal \N__78507\ : std_logic;
signal \N__78506\ : std_logic;
signal \N__78505\ : std_logic;
signal \N__78502\ : std_logic;
signal \N__78499\ : std_logic;
signal \N__78496\ : std_logic;
signal \N__78489\ : std_logic;
signal \N__78484\ : std_logic;
signal \N__78483\ : std_logic;
signal \N__78482\ : std_logic;
signal \N__78479\ : std_logic;
signal \N__78476\ : std_logic;
signal \N__78475\ : std_logic;
signal \N__78474\ : std_logic;
signal \N__78473\ : std_logic;
signal \N__78472\ : std_logic;
signal \N__78469\ : std_logic;
signal \N__78468\ : std_logic;
signal \N__78457\ : std_logic;
signal \N__78454\ : std_logic;
signal \N__78447\ : std_logic;
signal \N__78442\ : std_logic;
signal \N__78437\ : std_logic;
signal \N__78434\ : std_logic;
signal \N__78431\ : std_logic;
signal \N__78426\ : std_logic;
signal \N__78417\ : std_logic;
signal \N__78410\ : std_logic;
signal \N__78407\ : std_logic;
signal \N__78406\ : std_logic;
signal \N__78405\ : std_logic;
signal \N__78404\ : std_logic;
signal \N__78399\ : std_logic;
signal \N__78396\ : std_logic;
signal \N__78391\ : std_logic;
signal \N__78388\ : std_logic;
signal \N__78379\ : std_logic;
signal \N__78372\ : std_logic;
signal \N__78369\ : std_logic;
signal \N__78366\ : std_logic;
signal \N__78363\ : std_logic;
signal \N__78362\ : std_logic;
signal \N__78361\ : std_logic;
signal \N__78360\ : std_logic;
signal \N__78359\ : std_logic;
signal \N__78358\ : std_logic;
signal \N__78355\ : std_logic;
signal \N__78352\ : std_logic;
signal \N__78345\ : std_logic;
signal \N__78340\ : std_logic;
signal \N__78339\ : std_logic;
signal \N__78338\ : std_logic;
signal \N__78337\ : std_logic;
signal \N__78336\ : std_logic;
signal \N__78335\ : std_logic;
signal \N__78334\ : std_logic;
signal \N__78333\ : std_logic;
signal \N__78332\ : std_logic;
signal \N__78331\ : std_logic;
signal \N__78330\ : std_logic;
signal \N__78329\ : std_logic;
signal \N__78328\ : std_logic;
signal \N__78327\ : std_logic;
signal \N__78326\ : std_logic;
signal \N__78325\ : std_logic;
signal \N__78324\ : std_logic;
signal \N__78323\ : std_logic;
signal \N__78322\ : std_logic;
signal \N__78321\ : std_logic;
signal \N__78320\ : std_logic;
signal \N__78319\ : std_logic;
signal \N__78316\ : std_logic;
signal \N__78315\ : std_logic;
signal \N__78312\ : std_logic;
signal \N__78305\ : std_logic;
signal \N__78300\ : std_logic;
signal \N__78295\ : std_logic;
signal \N__78290\ : std_logic;
signal \N__78287\ : std_logic;
signal \N__78282\ : std_logic;
signal \N__78277\ : std_logic;
signal \N__78272\ : std_logic;
signal \N__78265\ : std_logic;
signal \N__78258\ : std_logic;
signal \N__78237\ : std_logic;
signal \N__78234\ : std_logic;
signal \N__78227\ : std_logic;
signal \N__78214\ : std_logic;
signal \N__78209\ : std_logic;
signal \N__78206\ : std_logic;
signal \N__78203\ : std_logic;
signal \N__78194\ : std_logic;
signal \N__78185\ : std_logic;
signal \N__78178\ : std_logic;
signal \N__78169\ : std_logic;
signal \N__78160\ : std_logic;
signal \N__78151\ : std_logic;
signal \N__78142\ : std_logic;
signal \N__78133\ : std_logic;
signal \N__78124\ : std_logic;
signal \N__78107\ : std_logic;
signal \N__78100\ : std_logic;
signal \N__78071\ : std_logic;
signal \N__78070\ : std_logic;
signal \N__78069\ : std_logic;
signal \N__78068\ : std_logic;
signal \N__78067\ : std_logic;
signal \N__78066\ : std_logic;
signal \N__78065\ : std_logic;
signal \N__78064\ : std_logic;
signal \N__78063\ : std_logic;
signal \N__78062\ : std_logic;
signal \N__78061\ : std_logic;
signal \N__78060\ : std_logic;
signal \N__78059\ : std_logic;
signal \N__78056\ : std_logic;
signal \N__78055\ : std_logic;
signal \N__78054\ : std_logic;
signal \N__78051\ : std_logic;
signal \N__78050\ : std_logic;
signal \N__78049\ : std_logic;
signal \N__78044\ : std_logic;
signal \N__78043\ : std_logic;
signal \N__78042\ : std_logic;
signal \N__78041\ : std_logic;
signal \N__78040\ : std_logic;
signal \N__78039\ : std_logic;
signal \N__78038\ : std_logic;
signal \N__78037\ : std_logic;
signal \N__78036\ : std_logic;
signal \N__78035\ : std_logic;
signal \N__78032\ : std_logic;
signal \N__78029\ : std_logic;
signal \N__78028\ : std_logic;
signal \N__78027\ : std_logic;
signal \N__78026\ : std_logic;
signal \N__78025\ : std_logic;
signal \N__78024\ : std_logic;
signal \N__78023\ : std_logic;
signal \N__78022\ : std_logic;
signal \N__78021\ : std_logic;
signal \N__78020\ : std_logic;
signal \N__78017\ : std_logic;
signal \N__78012\ : std_logic;
signal \N__78011\ : std_logic;
signal \N__78006\ : std_logic;
signal \N__78003\ : std_logic;
signal \N__77996\ : std_logic;
signal \N__77995\ : std_logic;
signal \N__77994\ : std_logic;
signal \N__77993\ : std_logic;
signal \N__77990\ : std_logic;
signal \N__77989\ : std_logic;
signal \N__77988\ : std_logic;
signal \N__77983\ : std_logic;
signal \N__77982\ : std_logic;
signal \N__77981\ : std_logic;
signal \N__77978\ : std_logic;
signal \N__77977\ : std_logic;
signal \N__77976\ : std_logic;
signal \N__77975\ : std_logic;
signal \N__77974\ : std_logic;
signal \N__77973\ : std_logic;
signal \N__77970\ : std_logic;
signal \N__77967\ : std_logic;
signal \N__77966\ : std_logic;
signal \N__77965\ : std_logic;
signal \N__77962\ : std_logic;
signal \N__77961\ : std_logic;
signal \N__77958\ : std_logic;
signal \N__77957\ : std_logic;
signal \N__77956\ : std_logic;
signal \N__77955\ : std_logic;
signal \N__77954\ : std_logic;
signal \N__77953\ : std_logic;
signal \N__77950\ : std_logic;
signal \N__77947\ : std_logic;
signal \N__77944\ : std_logic;
signal \N__77941\ : std_logic;
signal \N__77940\ : std_logic;
signal \N__77937\ : std_logic;
signal \N__77934\ : std_logic;
signal \N__77933\ : std_logic;
signal \N__77932\ : std_logic;
signal \N__77929\ : std_logic;
signal \N__77926\ : std_logic;
signal \N__77921\ : std_logic;
signal \N__77912\ : std_logic;
signal \N__77911\ : std_logic;
signal \N__77910\ : std_logic;
signal \N__77909\ : std_logic;
signal \N__77908\ : std_logic;
signal \N__77907\ : std_logic;
signal \N__77906\ : std_logic;
signal \N__77903\ : std_logic;
signal \N__77900\ : std_logic;
signal \N__77899\ : std_logic;
signal \N__77898\ : std_logic;
signal \N__77897\ : std_logic;
signal \N__77896\ : std_logic;
signal \N__77895\ : std_logic;
signal \N__77894\ : std_logic;
signal \N__77893\ : std_logic;
signal \N__77892\ : std_logic;
signal \N__77889\ : std_logic;
signal \N__77888\ : std_logic;
signal \N__77887\ : std_logic;
signal \N__77886\ : std_logic;
signal \N__77885\ : std_logic;
signal \N__77884\ : std_logic;
signal \N__77883\ : std_logic;
signal \N__77882\ : std_logic;
signal \N__77881\ : std_logic;
signal \N__77880\ : std_logic;
signal \N__77879\ : std_logic;
signal \N__77878\ : std_logic;
signal \N__77877\ : std_logic;
signal \N__77876\ : std_logic;
signal \N__77875\ : std_logic;
signal \N__77874\ : std_logic;
signal \N__77873\ : std_logic;
signal \N__77870\ : std_logic;
signal \N__77867\ : std_logic;
signal \N__77866\ : std_logic;
signal \N__77865\ : std_logic;
signal \N__77864\ : std_logic;
signal \N__77863\ : std_logic;
signal \N__77862\ : std_logic;
signal \N__77859\ : std_logic;
signal \N__77856\ : std_logic;
signal \N__77853\ : std_logic;
signal \N__77850\ : std_logic;
signal \N__77847\ : std_logic;
signal \N__77844\ : std_logic;
signal \N__77843\ : std_logic;
signal \N__77842\ : std_logic;
signal \N__77841\ : std_logic;
signal \N__77840\ : std_logic;
signal \N__77839\ : std_logic;
signal \N__77838\ : std_logic;
signal \N__77829\ : std_logic;
signal \N__77826\ : std_logic;
signal \N__77817\ : std_logic;
signal \N__77816\ : std_logic;
signal \N__77813\ : std_logic;
signal \N__77812\ : std_logic;
signal \N__77809\ : std_logic;
signal \N__77808\ : std_logic;
signal \N__77807\ : std_logic;
signal \N__77806\ : std_logic;
signal \N__77805\ : std_logic;
signal \N__77804\ : std_logic;
signal \N__77803\ : std_logic;
signal \N__77800\ : std_logic;
signal \N__77797\ : std_logic;
signal \N__77796\ : std_logic;
signal \N__77795\ : std_logic;
signal \N__77794\ : std_logic;
signal \N__77793\ : std_logic;
signal \N__77790\ : std_logic;
signal \N__77785\ : std_logic;
signal \N__77778\ : std_logic;
signal \N__77775\ : std_logic;
signal \N__77766\ : std_logic;
signal \N__77755\ : std_logic;
signal \N__77752\ : std_logic;
signal \N__77745\ : std_logic;
signal \N__77744\ : std_logic;
signal \N__77743\ : std_logic;
signal \N__77740\ : std_logic;
signal \N__77733\ : std_logic;
signal \N__77730\ : std_logic;
signal \N__77723\ : std_logic;
signal \N__77720\ : std_logic;
signal \N__77715\ : std_logic;
signal \N__77708\ : std_logic;
signal \N__77701\ : std_logic;
signal \N__77700\ : std_logic;
signal \N__77697\ : std_logic;
signal \N__77694\ : std_logic;
signal \N__77693\ : std_logic;
signal \N__77692\ : std_logic;
signal \N__77691\ : std_logic;
signal \N__77690\ : std_logic;
signal \N__77689\ : std_logic;
signal \N__77688\ : std_logic;
signal \N__77685\ : std_logic;
signal \N__77682\ : std_logic;
signal \N__77675\ : std_logic;
signal \N__77668\ : std_logic;
signal \N__77659\ : std_logic;
signal \N__77654\ : std_logic;
signal \N__77647\ : std_logic;
signal \N__77642\ : std_logic;
signal \N__77639\ : std_logic;
signal \N__77636\ : std_logic;
signal \N__77627\ : std_logic;
signal \N__77624\ : std_logic;
signal \N__77621\ : std_logic;
signal \N__77620\ : std_logic;
signal \N__77619\ : std_logic;
signal \N__77618\ : std_logic;
signal \N__77617\ : std_logic;
signal \N__77616\ : std_logic;
signal \N__77615\ : std_logic;
signal \N__77614\ : std_logic;
signal \N__77613\ : std_logic;
signal \N__77612\ : std_logic;
signal \N__77611\ : std_logic;
signal \N__77610\ : std_logic;
signal \N__77609\ : std_logic;
signal \N__77608\ : std_logic;
signal \N__77605\ : std_logic;
signal \N__77598\ : std_logic;
signal \N__77591\ : std_logic;
signal \N__77590\ : std_logic;
signal \N__77587\ : std_logic;
signal \N__77584\ : std_logic;
signal \N__77583\ : std_logic;
signal \N__77580\ : std_logic;
signal \N__77577\ : std_logic;
signal \N__77576\ : std_logic;
signal \N__77575\ : std_logic;
signal \N__77568\ : std_logic;
signal \N__77559\ : std_logic;
signal \N__77548\ : std_logic;
signal \N__77539\ : std_logic;
signal \N__77532\ : std_logic;
signal \N__77525\ : std_logic;
signal \N__77518\ : std_logic;
signal \N__77515\ : std_logic;
signal \N__77512\ : std_logic;
signal \N__77507\ : std_logic;
signal \N__77498\ : std_logic;
signal \N__77489\ : std_logic;
signal \N__77480\ : std_logic;
signal \N__77473\ : std_logic;
signal \N__77466\ : std_logic;
signal \N__77459\ : std_logic;
signal \N__77450\ : std_logic;
signal \N__77441\ : std_logic;
signal \N__77438\ : std_logic;
signal \N__77427\ : std_logic;
signal \N__77420\ : std_logic;
signal \N__77415\ : std_logic;
signal \N__77408\ : std_logic;
signal \N__77401\ : std_logic;
signal \N__77392\ : std_logic;
signal \N__77383\ : std_logic;
signal \N__77378\ : std_logic;
signal \N__77373\ : std_logic;
signal \N__77366\ : std_logic;
signal \N__77343\ : std_logic;
signal \N__77318\ : std_logic;
signal \N__77317\ : std_logic;
signal \N__77316\ : std_logic;
signal \N__77315\ : std_logic;
signal \N__77314\ : std_logic;
signal \N__77313\ : std_logic;
signal \N__77312\ : std_logic;
signal \N__77311\ : std_logic;
signal \N__77310\ : std_logic;
signal \N__77309\ : std_logic;
signal \N__77308\ : std_logic;
signal \N__77305\ : std_logic;
signal \N__77304\ : std_logic;
signal \N__77303\ : std_logic;
signal \N__77302\ : std_logic;
signal \N__77301\ : std_logic;
signal \N__77298\ : std_logic;
signal \N__77297\ : std_logic;
signal \N__77296\ : std_logic;
signal \N__77295\ : std_logic;
signal \N__77294\ : std_logic;
signal \N__77293\ : std_logic;
signal \N__77292\ : std_logic;
signal \N__77287\ : std_logic;
signal \N__77284\ : std_logic;
signal \N__77283\ : std_logic;
signal \N__77282\ : std_logic;
signal \N__77281\ : std_logic;
signal \N__77280\ : std_logic;
signal \N__77275\ : std_logic;
signal \N__77274\ : std_logic;
signal \N__77273\ : std_logic;
signal \N__77272\ : std_logic;
signal \N__77271\ : std_logic;
signal \N__77268\ : std_logic;
signal \N__77265\ : std_logic;
signal \N__77262\ : std_logic;
signal \N__77259\ : std_logic;
signal \N__77258\ : std_logic;
signal \N__77257\ : std_logic;
signal \N__77256\ : std_logic;
signal \N__77255\ : std_logic;
signal \N__77254\ : std_logic;
signal \N__77253\ : std_logic;
signal \N__77252\ : std_logic;
signal \N__77251\ : std_logic;
signal \N__77250\ : std_logic;
signal \N__77249\ : std_logic;
signal \N__77248\ : std_logic;
signal \N__77247\ : std_logic;
signal \N__77246\ : std_logic;
signal \N__77245\ : std_logic;
signal \N__77244\ : std_logic;
signal \N__77243\ : std_logic;
signal \N__77242\ : std_logic;
signal \N__77241\ : std_logic;
signal \N__77240\ : std_logic;
signal \N__77239\ : std_logic;
signal \N__77238\ : std_logic;
signal \N__77237\ : std_logic;
signal \N__77236\ : std_logic;
signal \N__77235\ : std_logic;
signal \N__77234\ : std_logic;
signal \N__77231\ : std_logic;
signal \N__77222\ : std_logic;
signal \N__77219\ : std_logic;
signal \N__77214\ : std_logic;
signal \N__77205\ : std_logic;
signal \N__77202\ : std_logic;
signal \N__77201\ : std_logic;
signal \N__77200\ : std_logic;
signal \N__77199\ : std_logic;
signal \N__77198\ : std_logic;
signal \N__77197\ : std_logic;
signal \N__77196\ : std_logic;
signal \N__77193\ : std_logic;
signal \N__77192\ : std_logic;
signal \N__77191\ : std_logic;
signal \N__77190\ : std_logic;
signal \N__77189\ : std_logic;
signal \N__77188\ : std_logic;
signal \N__77187\ : std_logic;
signal \N__77186\ : std_logic;
signal \N__77185\ : std_logic;
signal \N__77184\ : std_logic;
signal \N__77183\ : std_logic;
signal \N__77182\ : std_logic;
signal \N__77181\ : std_logic;
signal \N__77176\ : std_logic;
signal \N__77175\ : std_logic;
signal \N__77174\ : std_logic;
signal \N__77173\ : std_logic;
signal \N__77172\ : std_logic;
signal \N__77171\ : std_logic;
signal \N__77166\ : std_logic;
signal \N__77165\ : std_logic;
signal \N__77164\ : std_logic;
signal \N__77161\ : std_logic;
signal \N__77152\ : std_logic;
signal \N__77151\ : std_logic;
signal \N__77150\ : std_logic;
signal \N__77149\ : std_logic;
signal \N__77148\ : std_logic;
signal \N__77147\ : std_logic;
signal \N__77146\ : std_logic;
signal \N__77145\ : std_logic;
signal \N__77144\ : std_logic;
signal \N__77143\ : std_logic;
signal \N__77142\ : std_logic;
signal \N__77141\ : std_logic;
signal \N__77140\ : std_logic;
signal \N__77137\ : std_logic;
signal \N__77132\ : std_logic;
signal \N__77129\ : std_logic;
signal \N__77126\ : std_logic;
signal \N__77125\ : std_logic;
signal \N__77124\ : std_logic;
signal \N__77123\ : std_logic;
signal \N__77122\ : std_logic;
signal \N__77121\ : std_logic;
signal \N__77120\ : std_logic;
signal \N__77119\ : std_logic;
signal \N__77118\ : std_logic;
signal \N__77117\ : std_logic;
signal \N__77116\ : std_logic;
signal \N__77115\ : std_logic;
signal \N__77114\ : std_logic;
signal \N__77109\ : std_logic;
signal \N__77100\ : std_logic;
signal \N__77093\ : std_logic;
signal \N__77088\ : std_logic;
signal \N__77081\ : std_logic;
signal \N__77074\ : std_logic;
signal \N__77073\ : std_logic;
signal \N__77072\ : std_logic;
signal \N__77071\ : std_logic;
signal \N__77070\ : std_logic;
signal \N__77069\ : std_logic;
signal \N__77068\ : std_logic;
signal \N__77067\ : std_logic;
signal \N__77066\ : std_logic;
signal \N__77065\ : std_logic;
signal \N__77062\ : std_logic;
signal \N__77055\ : std_logic;
signal \N__77048\ : std_logic;
signal \N__77039\ : std_logic;
signal \N__77034\ : std_logic;
signal \N__77027\ : std_logic;
signal \N__77020\ : std_logic;
signal \N__77017\ : std_logic;
signal \N__77010\ : std_logic;
signal \N__77003\ : std_logic;
signal \N__76998\ : std_logic;
signal \N__76995\ : std_logic;
signal \N__76988\ : std_logic;
signal \N__76985\ : std_logic;
signal \N__76982\ : std_logic;
signal \N__76979\ : std_logic;
signal \N__76978\ : std_logic;
signal \N__76977\ : std_logic;
signal \N__76970\ : std_logic;
signal \N__76967\ : std_logic;
signal \N__76966\ : std_logic;
signal \N__76965\ : std_logic;
signal \N__76960\ : std_logic;
signal \N__76957\ : std_logic;
signal \N__76954\ : std_logic;
signal \N__76947\ : std_logic;
signal \N__76938\ : std_logic;
signal \N__76937\ : std_logic;
signal \N__76936\ : std_logic;
signal \N__76935\ : std_logic;
signal \N__76934\ : std_logic;
signal \N__76933\ : std_logic;
signal \N__76932\ : std_logic;
signal \N__76931\ : std_logic;
signal \N__76930\ : std_logic;
signal \N__76929\ : std_logic;
signal \N__76928\ : std_logic;
signal \N__76927\ : std_logic;
signal \N__76926\ : std_logic;
signal \N__76925\ : std_logic;
signal \N__76914\ : std_logic;
signal \N__76913\ : std_logic;
signal \N__76912\ : std_logic;
signal \N__76911\ : std_logic;
signal \N__76910\ : std_logic;
signal \N__76909\ : std_logic;
signal \N__76904\ : std_logic;
signal \N__76899\ : std_logic;
signal \N__76890\ : std_logic;
signal \N__76879\ : std_logic;
signal \N__76872\ : std_logic;
signal \N__76865\ : std_logic;
signal \N__76858\ : std_logic;
signal \N__76851\ : std_logic;
signal \N__76838\ : std_logic;
signal \N__76831\ : std_logic;
signal \N__76822\ : std_logic;
signal \N__76811\ : std_logic;
signal \N__76802\ : std_logic;
signal \N__76797\ : std_logic;
signal \N__76792\ : std_logic;
signal \N__76787\ : std_logic;
signal \N__76784\ : std_logic;
signal \N__76775\ : std_logic;
signal \N__76762\ : std_logic;
signal \N__76753\ : std_logic;
signal \N__76746\ : std_logic;
signal \N__76743\ : std_logic;
signal \N__76732\ : std_logic;
signal \N__76723\ : std_logic;
signal \N__76704\ : std_logic;
signal \N__76679\ : std_logic;
signal \N__76676\ : std_logic;
signal \N__76673\ : std_logic;
signal \N__76670\ : std_logic;
signal \N__76667\ : std_logic;
signal \N__76664\ : std_logic;
signal \N__76661\ : std_logic;
signal \N__76658\ : std_logic;
signal \N__76655\ : std_logic;
signal \N__76652\ : std_logic;
signal \N__76649\ : std_logic;
signal \N__76648\ : std_logic;
signal \N__76645\ : std_logic;
signal \N__76642\ : std_logic;
signal \N__76637\ : std_logic;
signal \N__76636\ : std_logic;
signal \N__76635\ : std_logic;
signal \N__76634\ : std_logic;
signal \N__76633\ : std_logic;
signal \N__76626\ : std_logic;
signal \N__76625\ : std_logic;
signal \N__76624\ : std_logic;
signal \N__76623\ : std_logic;
signal \N__76620\ : std_logic;
signal \N__76619\ : std_logic;
signal \N__76618\ : std_logic;
signal \N__76617\ : std_logic;
signal \N__76616\ : std_logic;
signal \N__76613\ : std_logic;
signal \N__76610\ : std_logic;
signal \N__76609\ : std_logic;
signal \N__76608\ : std_logic;
signal \N__76607\ : std_logic;
signal \N__76606\ : std_logic;
signal \N__76605\ : std_logic;
signal \N__76604\ : std_logic;
signal \N__76603\ : std_logic;
signal \N__76602\ : std_logic;
signal \N__76601\ : std_logic;
signal \N__76600\ : std_logic;
signal \N__76597\ : std_logic;
signal \N__76594\ : std_logic;
signal \N__76593\ : std_logic;
signal \N__76592\ : std_logic;
signal \N__76591\ : std_logic;
signal \N__76588\ : std_logic;
signal \N__76587\ : std_logic;
signal \N__76586\ : std_logic;
signal \N__76585\ : std_logic;
signal \N__76584\ : std_logic;
signal \N__76583\ : std_logic;
signal \N__76580\ : std_logic;
signal \N__76579\ : std_logic;
signal \N__76576\ : std_logic;
signal \N__76575\ : std_logic;
signal \N__76574\ : std_logic;
signal \N__76573\ : std_logic;
signal \N__76572\ : std_logic;
signal \N__76571\ : std_logic;
signal \N__76570\ : std_logic;
signal \N__76569\ : std_logic;
signal \N__76566\ : std_logic;
signal \N__76563\ : std_logic;
signal \N__76560\ : std_logic;
signal \N__76559\ : std_logic;
signal \N__76554\ : std_logic;
signal \N__76551\ : std_logic;
signal \N__76546\ : std_logic;
signal \N__76541\ : std_logic;
signal \N__76536\ : std_logic;
signal \N__76535\ : std_logic;
signal \N__76534\ : std_logic;
signal \N__76533\ : std_logic;
signal \N__76532\ : std_logic;
signal \N__76531\ : std_logic;
signal \N__76530\ : std_logic;
signal \N__76529\ : std_logic;
signal \N__76528\ : std_logic;
signal \N__76527\ : std_logic;
signal \N__76526\ : std_logic;
signal \N__76523\ : std_logic;
signal \N__76522\ : std_logic;
signal \N__76519\ : std_logic;
signal \N__76516\ : std_logic;
signal \N__76513\ : std_logic;
signal \N__76510\ : std_logic;
signal \N__76507\ : std_logic;
signal \N__76504\ : std_logic;
signal \N__76501\ : std_logic;
signal \N__76500\ : std_logic;
signal \N__76499\ : std_logic;
signal \N__76498\ : std_logic;
signal \N__76493\ : std_logic;
signal \N__76486\ : std_logic;
signal \N__76485\ : std_logic;
signal \N__76484\ : std_logic;
signal \N__76483\ : std_logic;
signal \N__76482\ : std_logic;
signal \N__76481\ : std_logic;
signal \N__76480\ : std_logic;
signal \N__76479\ : std_logic;
signal \N__76476\ : std_logic;
signal \N__76475\ : std_logic;
signal \N__76474\ : std_logic;
signal \N__76473\ : std_logic;
signal \N__76472\ : std_logic;
signal \N__76471\ : std_logic;
signal \N__76470\ : std_logic;
signal \N__76467\ : std_logic;
signal \N__76464\ : std_logic;
signal \N__76463\ : std_logic;
signal \N__76462\ : std_logic;
signal \N__76461\ : std_logic;
signal \N__76460\ : std_logic;
signal \N__76459\ : std_logic;
signal \N__76458\ : std_logic;
signal \N__76455\ : std_logic;
signal \N__76454\ : std_logic;
signal \N__76449\ : std_logic;
signal \N__76448\ : std_logic;
signal \N__76447\ : std_logic;
signal \N__76446\ : std_logic;
signal \N__76441\ : std_logic;
signal \N__76434\ : std_logic;
signal \N__76429\ : std_logic;
signal \N__76424\ : std_logic;
signal \N__76421\ : std_logic;
signal \N__76414\ : std_logic;
signal \N__76411\ : std_logic;
signal \N__76406\ : std_logic;
signal \N__76405\ : std_logic;
signal \N__76404\ : std_logic;
signal \N__76403\ : std_logic;
signal \N__76396\ : std_logic;
signal \N__76391\ : std_logic;
signal \N__76388\ : std_logic;
signal \N__76381\ : std_logic;
signal \N__76378\ : std_logic;
signal \N__76375\ : std_logic;
signal \N__76374\ : std_logic;
signal \N__76373\ : std_logic;
signal \N__76372\ : std_logic;
signal \N__76369\ : std_logic;
signal \N__76362\ : std_logic;
signal \N__76357\ : std_logic;
signal \N__76354\ : std_logic;
signal \N__76351\ : std_logic;
signal \N__76350\ : std_logic;
signal \N__76349\ : std_logic;
signal \N__76346\ : std_logic;
signal \N__76341\ : std_logic;
signal \N__76336\ : std_logic;
signal \N__76331\ : std_logic;
signal \N__76326\ : std_logic;
signal \N__76323\ : std_logic;
signal \N__76322\ : std_logic;
signal \N__76321\ : std_logic;
signal \N__76318\ : std_logic;
signal \N__76313\ : std_logic;
signal \N__76310\ : std_logic;
signal \N__76305\ : std_logic;
signal \N__76302\ : std_logic;
signal \N__76299\ : std_logic;
signal \N__76294\ : std_logic;
signal \N__76293\ : std_logic;
signal \N__76292\ : std_logic;
signal \N__76291\ : std_logic;
signal \N__76288\ : std_logic;
signal \N__76287\ : std_logic;
signal \N__76286\ : std_logic;
signal \N__76277\ : std_logic;
signal \N__76274\ : std_logic;
signal \N__76273\ : std_logic;
signal \N__76272\ : std_logic;
signal \N__76271\ : std_logic;
signal \N__76270\ : std_logic;
signal \N__76269\ : std_logic;
signal \N__76268\ : std_logic;
signal \N__76265\ : std_logic;
signal \N__76264\ : std_logic;
signal \N__76263\ : std_logic;
signal \N__76262\ : std_logic;
signal \N__76261\ : std_logic;
signal \N__76258\ : std_logic;
signal \N__76251\ : std_logic;
signal \N__76248\ : std_logic;
signal \N__76241\ : std_logic;
signal \N__76232\ : std_logic;
signal \N__76225\ : std_logic;
signal \N__76222\ : std_logic;
signal \N__76215\ : std_logic;
signal \N__76210\ : std_logic;
signal \N__76203\ : std_logic;
signal \N__76192\ : std_logic;
signal \N__76185\ : std_logic;
signal \N__76174\ : std_logic;
signal \N__76173\ : std_logic;
signal \N__76168\ : std_logic;
signal \N__76159\ : std_logic;
signal \N__76152\ : std_logic;
signal \N__76145\ : std_logic;
signal \N__76142\ : std_logic;
signal \N__76139\ : std_logic;
signal \N__76136\ : std_logic;
signal \N__76131\ : std_logic;
signal \N__76128\ : std_logic;
signal \N__76123\ : std_logic;
signal \N__76118\ : std_logic;
signal \N__76113\ : std_logic;
signal \N__76110\ : std_logic;
signal \N__76103\ : std_logic;
signal \N__76098\ : std_logic;
signal \N__76089\ : std_logic;
signal \N__76074\ : std_logic;
signal \N__76071\ : std_logic;
signal \N__76062\ : std_logic;
signal \N__76059\ : std_logic;
signal \N__76028\ : std_logic;
signal \N__76025\ : std_logic;
signal \N__76022\ : std_logic;
signal \N__76019\ : std_logic;
signal \N__76016\ : std_logic;
signal \N__76015\ : std_logic;
signal \N__76012\ : std_logic;
signal \N__76011\ : std_logic;
signal \N__76010\ : std_logic;
signal \N__76009\ : std_logic;
signal \N__76008\ : std_logic;
signal \N__76005\ : std_logic;
signal \N__76004\ : std_logic;
signal \N__76003\ : std_logic;
signal \N__76002\ : std_logic;
signal \N__75997\ : std_logic;
signal \N__75996\ : std_logic;
signal \N__75995\ : std_logic;
signal \N__75994\ : std_logic;
signal \N__75993\ : std_logic;
signal \N__75992\ : std_logic;
signal \N__75991\ : std_logic;
signal \N__75990\ : std_logic;
signal \N__75987\ : std_logic;
signal \N__75986\ : std_logic;
signal \N__75985\ : std_logic;
signal \N__75984\ : std_logic;
signal \N__75983\ : std_logic;
signal \N__75980\ : std_logic;
signal \N__75977\ : std_logic;
signal \N__75974\ : std_logic;
signal \N__75973\ : std_logic;
signal \N__75970\ : std_logic;
signal \N__75969\ : std_logic;
signal \N__75968\ : std_logic;
signal \N__75967\ : std_logic;
signal \N__75966\ : std_logic;
signal \N__75965\ : std_logic;
signal \N__75964\ : std_logic;
signal \N__75963\ : std_logic;
signal \N__75962\ : std_logic;
signal \N__75961\ : std_logic;
signal \N__75960\ : std_logic;
signal \N__75959\ : std_logic;
signal \N__75956\ : std_logic;
signal \N__75955\ : std_logic;
signal \N__75954\ : std_logic;
signal \N__75951\ : std_logic;
signal \N__75950\ : std_logic;
signal \N__75947\ : std_logic;
signal \N__75942\ : std_logic;
signal \N__75941\ : std_logic;
signal \N__75940\ : std_logic;
signal \N__75939\ : std_logic;
signal \N__75938\ : std_logic;
signal \N__75935\ : std_logic;
signal \N__75934\ : std_logic;
signal \N__75933\ : std_logic;
signal \N__75932\ : std_logic;
signal \N__75929\ : std_logic;
signal \N__75926\ : std_logic;
signal \N__75923\ : std_logic;
signal \N__75920\ : std_logic;
signal \N__75919\ : std_logic;
signal \N__75918\ : std_logic;
signal \N__75917\ : std_logic;
signal \N__75916\ : std_logic;
signal \N__75915\ : std_logic;
signal \N__75914\ : std_logic;
signal \N__75913\ : std_logic;
signal \N__75912\ : std_logic;
signal \N__75911\ : std_logic;
signal \N__75910\ : std_logic;
signal \N__75909\ : std_logic;
signal \N__75908\ : std_logic;
signal \N__75907\ : std_logic;
signal \N__75906\ : std_logic;
signal \N__75905\ : std_logic;
signal \N__75904\ : std_logic;
signal \N__75903\ : std_logic;
signal \N__75902\ : std_logic;
signal \N__75901\ : std_logic;
signal \N__75900\ : std_logic;
signal \N__75899\ : std_logic;
signal \N__75896\ : std_logic;
signal \N__75893\ : std_logic;
signal \N__75892\ : std_logic;
signal \N__75891\ : std_logic;
signal \N__75890\ : std_logic;
signal \N__75889\ : std_logic;
signal \N__75888\ : std_logic;
signal \N__75887\ : std_logic;
signal \N__75886\ : std_logic;
signal \N__75885\ : std_logic;
signal \N__75882\ : std_logic;
signal \N__75881\ : std_logic;
signal \N__75880\ : std_logic;
signal \N__75879\ : std_logic;
signal \N__75876\ : std_logic;
signal \N__75871\ : std_logic;
signal \N__75868\ : std_logic;
signal \N__75865\ : std_logic;
signal \N__75860\ : std_logic;
signal \N__75857\ : std_logic;
signal \N__75856\ : std_logic;
signal \N__75853\ : std_logic;
signal \N__75852\ : std_logic;
signal \N__75851\ : std_logic;
signal \N__75848\ : std_logic;
signal \N__75847\ : std_logic;
signal \N__75846\ : std_logic;
signal \N__75843\ : std_logic;
signal \N__75840\ : std_logic;
signal \N__75839\ : std_logic;
signal \N__75836\ : std_logic;
signal \N__75833\ : std_logic;
signal \N__75832\ : std_logic;
signal \N__75831\ : std_logic;
signal \N__75830\ : std_logic;
signal \N__75829\ : std_logic;
signal \N__75828\ : std_logic;
signal \N__75825\ : std_logic;
signal \N__75822\ : std_logic;
signal \N__75821\ : std_logic;
signal \N__75818\ : std_logic;
signal \N__75817\ : std_logic;
signal \N__75816\ : std_logic;
signal \N__75815\ : std_logic;
signal \N__75814\ : std_logic;
signal \N__75811\ : std_logic;
signal \N__75810\ : std_logic;
signal \N__75809\ : std_logic;
signal \N__75808\ : std_logic;
signal \N__75805\ : std_logic;
signal \N__75804\ : std_logic;
signal \N__75801\ : std_logic;
signal \N__75800\ : std_logic;
signal \N__75799\ : std_logic;
signal \N__75796\ : std_logic;
signal \N__75795\ : std_logic;
signal \N__75792\ : std_logic;
signal \N__75791\ : std_logic;
signal \N__75790\ : std_logic;
signal \N__75789\ : std_logic;
signal \N__75786\ : std_logic;
signal \N__75781\ : std_logic;
signal \N__75770\ : std_logic;
signal \N__75763\ : std_logic;
signal \N__75754\ : std_logic;
signal \N__75751\ : std_logic;
signal \N__75750\ : std_logic;
signal \N__75747\ : std_logic;
signal \N__75746\ : std_logic;
signal \N__75743\ : std_logic;
signal \N__75740\ : std_logic;
signal \N__75737\ : std_logic;
signal \N__75736\ : std_logic;
signal \N__75733\ : std_logic;
signal \N__75730\ : std_logic;
signal \N__75727\ : std_logic;
signal \N__75726\ : std_logic;
signal \N__75725\ : std_logic;
signal \N__75722\ : std_logic;
signal \N__75721\ : std_logic;
signal \N__75720\ : std_logic;
signal \N__75719\ : std_logic;
signal \N__75718\ : std_logic;
signal \N__75715\ : std_logic;
signal \N__75712\ : std_logic;
signal \N__75711\ : std_logic;
signal \N__75710\ : std_logic;
signal \N__75709\ : std_logic;
signal \N__75708\ : std_logic;
signal \N__75705\ : std_logic;
signal \N__75702\ : std_logic;
signal \N__75695\ : std_logic;
signal \N__75692\ : std_logic;
signal \N__75689\ : std_logic;
signal \N__75688\ : std_logic;
signal \N__75685\ : std_logic;
signal \N__75684\ : std_logic;
signal \N__75681\ : std_logic;
signal \N__75680\ : std_logic;
signal \N__75677\ : std_logic;
signal \N__75676\ : std_logic;
signal \N__75673\ : std_logic;
signal \N__75672\ : std_logic;
signal \N__75671\ : std_logic;
signal \N__75670\ : std_logic;
signal \N__75669\ : std_logic;
signal \N__75668\ : std_logic;
signal \N__75665\ : std_logic;
signal \N__75660\ : std_logic;
signal \N__75659\ : std_logic;
signal \N__75656\ : std_logic;
signal \N__75655\ : std_logic;
signal \N__75654\ : std_logic;
signal \N__75653\ : std_logic;
signal \N__75650\ : std_logic;
signal \N__75647\ : std_logic;
signal \N__75646\ : std_logic;
signal \N__75645\ : std_logic;
signal \N__75642\ : std_logic;
signal \N__75639\ : std_logic;
signal \N__75638\ : std_logic;
signal \N__75637\ : std_logic;
signal \N__75636\ : std_logic;
signal \N__75635\ : std_logic;
signal \N__75632\ : std_logic;
signal \N__75631\ : std_logic;
signal \N__75630\ : std_logic;
signal \N__75627\ : std_logic;
signal \N__75620\ : std_logic;
signal \N__75619\ : std_logic;
signal \N__75616\ : std_logic;
signal \N__75615\ : std_logic;
signal \N__75614\ : std_logic;
signal \N__75613\ : std_logic;
signal \N__75612\ : std_logic;
signal \N__75611\ : std_logic;
signal \N__75606\ : std_logic;
signal \N__75599\ : std_logic;
signal \N__75598\ : std_logic;
signal \N__75597\ : std_logic;
signal \N__75594\ : std_logic;
signal \N__75587\ : std_logic;
signal \N__75580\ : std_logic;
signal \N__75577\ : std_logic;
signal \N__75570\ : std_logic;
signal \N__75561\ : std_logic;
signal \N__75556\ : std_logic;
signal \N__75551\ : std_logic;
signal \N__75546\ : std_logic;
signal \N__75541\ : std_logic;
signal \N__75540\ : std_logic;
signal \N__75539\ : std_logic;
signal \N__75538\ : std_logic;
signal \N__75535\ : std_logic;
signal \N__75534\ : std_logic;
signal \N__75533\ : std_logic;
signal \N__75530\ : std_logic;
signal \N__75529\ : std_logic;
signal \N__75528\ : std_logic;
signal \N__75527\ : std_logic;
signal \N__75526\ : std_logic;
signal \N__75521\ : std_logic;
signal \N__75516\ : std_logic;
signal \N__75513\ : std_logic;
signal \N__75502\ : std_logic;
signal \N__75501\ : std_logic;
signal \N__75500\ : std_logic;
signal \N__75499\ : std_logic;
signal \N__75496\ : std_logic;
signal \N__75493\ : std_logic;
signal \N__75490\ : std_logic;
signal \N__75483\ : std_logic;
signal \N__75474\ : std_logic;
signal \N__75467\ : std_logic;
signal \N__75460\ : std_logic;
signal \N__75453\ : std_logic;
signal \N__75446\ : std_logic;
signal \N__75439\ : std_logic;
signal \N__75430\ : std_logic;
signal \N__75425\ : std_logic;
signal \N__75424\ : std_logic;
signal \N__75423\ : std_logic;
signal \N__75422\ : std_logic;
signal \N__75419\ : std_logic;
signal \N__75416\ : std_logic;
signal \N__75413\ : std_logic;
signal \N__75410\ : std_logic;
signal \N__75407\ : std_logic;
signal \N__75404\ : std_logic;
signal \N__75401\ : std_logic;
signal \N__75394\ : std_logic;
signal \N__75385\ : std_logic;
signal \N__75384\ : std_logic;
signal \N__75383\ : std_logic;
signal \N__75380\ : std_logic;
signal \N__75377\ : std_logic;
signal \N__75366\ : std_logic;
signal \N__75361\ : std_logic;
signal \N__75348\ : std_logic;
signal \N__75339\ : std_logic;
signal \N__75336\ : std_logic;
signal \N__75329\ : std_logic;
signal \N__75320\ : std_logic;
signal \N__75317\ : std_logic;
signal \N__75314\ : std_logic;
signal \N__75311\ : std_logic;
signal \N__75308\ : std_logic;
signal \N__75307\ : std_logic;
signal \N__75306\ : std_logic;
signal \N__75305\ : std_logic;
signal \N__75304\ : std_logic;
signal \N__75303\ : std_logic;
signal \N__75300\ : std_logic;
signal \N__75299\ : std_logic;
signal \N__75296\ : std_logic;
signal \N__75293\ : std_logic;
signal \N__75292\ : std_logic;
signal \N__75291\ : std_logic;
signal \N__75288\ : std_logic;
signal \N__75287\ : std_logic;
signal \N__75284\ : std_logic;
signal \N__75283\ : std_logic;
signal \N__75280\ : std_logic;
signal \N__75277\ : std_logic;
signal \N__75272\ : std_logic;
signal \N__75263\ : std_logic;
signal \N__75258\ : std_logic;
signal \N__75249\ : std_logic;
signal \N__75248\ : std_logic;
signal \N__75247\ : std_logic;
signal \N__75244\ : std_logic;
signal \N__75243\ : std_logic;
signal \N__75240\ : std_logic;
signal \N__75237\ : std_logic;
signal \N__75236\ : std_logic;
signal \N__75235\ : std_logic;
signal \N__75234\ : std_logic;
signal \N__75231\ : std_logic;
signal \N__75224\ : std_logic;
signal \N__75215\ : std_logic;
signal \N__75212\ : std_logic;
signal \N__75205\ : std_logic;
signal \N__75196\ : std_logic;
signal \N__75179\ : std_logic;
signal \N__75172\ : std_logic;
signal \N__75161\ : std_logic;
signal \N__75158\ : std_logic;
signal \N__75151\ : std_logic;
signal \N__75144\ : std_logic;
signal \N__75137\ : std_logic;
signal \N__75126\ : std_logic;
signal \N__75123\ : std_logic;
signal \N__75118\ : std_logic;
signal \N__75109\ : std_logic;
signal \N__75106\ : std_logic;
signal \N__75101\ : std_logic;
signal \N__75090\ : std_logic;
signal \N__75083\ : std_logic;
signal \N__75074\ : std_logic;
signal \N__75061\ : std_logic;
signal \N__75050\ : std_logic;
signal \N__75041\ : std_logic;
signal \N__75034\ : std_logic;
signal \N__75021\ : std_logic;
signal \N__75010\ : std_logic;
signal \N__75003\ : std_logic;
signal \N__74978\ : std_logic;
signal \N__74975\ : std_logic;
signal \N__74972\ : std_logic;
signal \N__74969\ : std_logic;
signal \N__74966\ : std_logic;
signal \N__74963\ : std_logic;
signal \N__74962\ : std_logic;
signal \N__74959\ : std_logic;
signal \N__74956\ : std_logic;
signal \N__74953\ : std_logic;
signal \N__74950\ : std_logic;
signal \N__74945\ : std_logic;
signal \N__74942\ : std_logic;
signal \N__74939\ : std_logic;
signal \N__74936\ : std_logic;
signal \N__74933\ : std_logic;
signal \N__74930\ : std_logic;
signal \N__74927\ : std_logic;
signal \N__74924\ : std_logic;
signal \N__74921\ : std_logic;
signal \N__74918\ : std_logic;
signal \N__74915\ : std_logic;
signal \N__74912\ : std_logic;
signal \N__74909\ : std_logic;
signal \N__74906\ : std_logic;
signal \N__74903\ : std_logic;
signal \N__74902\ : std_logic;
signal \N__74899\ : std_logic;
signal \N__74896\ : std_logic;
signal \N__74895\ : std_logic;
signal \N__74894\ : std_logic;
signal \N__74891\ : std_logic;
signal \N__74890\ : std_logic;
signal \N__74889\ : std_logic;
signal \N__74888\ : std_logic;
signal \N__74887\ : std_logic;
signal \N__74886\ : std_logic;
signal \N__74883\ : std_logic;
signal \N__74882\ : std_logic;
signal \N__74879\ : std_logic;
signal \N__74876\ : std_logic;
signal \N__74873\ : std_logic;
signal \N__74870\ : std_logic;
signal \N__74867\ : std_logic;
signal \N__74864\ : std_logic;
signal \N__74861\ : std_logic;
signal \N__74860\ : std_logic;
signal \N__74857\ : std_logic;
signal \N__74856\ : std_logic;
signal \N__74855\ : std_logic;
signal \N__74854\ : std_logic;
signal \N__74853\ : std_logic;
signal \N__74850\ : std_logic;
signal \N__74847\ : std_logic;
signal \N__74844\ : std_logic;
signal \N__74841\ : std_logic;
signal \N__74838\ : std_logic;
signal \N__74835\ : std_logic;
signal \N__74834\ : std_logic;
signal \N__74833\ : std_logic;
signal \N__74832\ : std_logic;
signal \N__74827\ : std_logic;
signal \N__74826\ : std_logic;
signal \N__74825\ : std_logic;
signal \N__74824\ : std_logic;
signal \N__74817\ : std_logic;
signal \N__74816\ : std_logic;
signal \N__74815\ : std_logic;
signal \N__74812\ : std_logic;
signal \N__74809\ : std_logic;
signal \N__74804\ : std_logic;
signal \N__74801\ : std_logic;
signal \N__74798\ : std_logic;
signal \N__74793\ : std_logic;
signal \N__74788\ : std_logic;
signal \N__74785\ : std_logic;
signal \N__74782\ : std_logic;
signal \N__74779\ : std_logic;
signal \N__74778\ : std_logic;
signal \N__74775\ : std_logic;
signal \N__74772\ : std_logic;
signal \N__74771\ : std_logic;
signal \N__74768\ : std_logic;
signal \N__74765\ : std_logic;
signal \N__74762\ : std_logic;
signal \N__74759\ : std_logic;
signal \N__74756\ : std_logic;
signal \N__74753\ : std_logic;
signal \N__74750\ : std_logic;
signal \N__74739\ : std_logic;
signal \N__74736\ : std_logic;
signal \N__74733\ : std_logic;
signal \N__74730\ : std_logic;
signal \N__74727\ : std_logic;
signal \N__74724\ : std_logic;
signal \N__74715\ : std_logic;
signal \N__74712\ : std_logic;
signal \N__74709\ : std_logic;
signal \N__74706\ : std_logic;
signal \N__74703\ : std_logic;
signal \N__74700\ : std_logic;
signal \N__74697\ : std_logic;
signal \N__74694\ : std_logic;
signal \N__74691\ : std_logic;
signal \N__74686\ : std_logic;
signal \N__74683\ : std_logic;
signal \N__74682\ : std_logic;
signal \N__74681\ : std_logic;
signal \N__74674\ : std_logic;
signal \N__74671\ : std_logic;
signal \N__74666\ : std_logic;
signal \N__74663\ : std_logic;
signal \N__74658\ : std_logic;
signal \N__74655\ : std_logic;
signal \N__74652\ : std_logic;
signal \N__74649\ : std_logic;
signal \N__74646\ : std_logic;
signal \N__74643\ : std_logic;
signal \N__74636\ : std_logic;
signal \N__74629\ : std_logic;
signal \N__74618\ : std_logic;
signal \N__74615\ : std_logic;
signal \N__74612\ : std_logic;
signal \N__74609\ : std_logic;
signal \N__74608\ : std_logic;
signal \N__74607\ : std_logic;
signal \N__74604\ : std_logic;
signal \N__74603\ : std_logic;
signal \N__74600\ : std_logic;
signal \N__74597\ : std_logic;
signal \N__74596\ : std_logic;
signal \N__74593\ : std_logic;
signal \N__74590\ : std_logic;
signal \N__74587\ : std_logic;
signal \N__74584\ : std_logic;
signal \N__74581\ : std_logic;
signal \N__74578\ : std_logic;
signal \N__74575\ : std_logic;
signal \N__74572\ : std_logic;
signal \N__74571\ : std_logic;
signal \N__74570\ : std_logic;
signal \N__74569\ : std_logic;
signal \N__74566\ : std_logic;
signal \N__74563\ : std_logic;
signal \N__74560\ : std_logic;
signal \N__74555\ : std_logic;
signal \N__74548\ : std_logic;
signal \N__74545\ : std_logic;
signal \N__74542\ : std_logic;
signal \N__74539\ : std_logic;
signal \N__74528\ : std_logic;
signal \N__74525\ : std_logic;
signal \N__74524\ : std_logic;
signal \N__74521\ : std_logic;
signal \N__74518\ : std_logic;
signal \N__74515\ : std_logic;
signal \N__74512\ : std_logic;
signal \N__74507\ : std_logic;
signal \N__74504\ : std_logic;
signal \N__74501\ : std_logic;
signal \N__74498\ : std_logic;
signal \N__74495\ : std_logic;
signal \N__74492\ : std_logic;
signal \N__74491\ : std_logic;
signal \N__74490\ : std_logic;
signal \N__74489\ : std_logic;
signal \N__74488\ : std_logic;
signal \N__74487\ : std_logic;
signal \N__74484\ : std_logic;
signal \N__74481\ : std_logic;
signal \N__74480\ : std_logic;
signal \N__74477\ : std_logic;
signal \N__74474\ : std_logic;
signal \N__74471\ : std_logic;
signal \N__74468\ : std_logic;
signal \N__74465\ : std_logic;
signal \N__74462\ : std_logic;
signal \N__74459\ : std_logic;
signal \N__74454\ : std_logic;
signal \N__74451\ : std_logic;
signal \N__74448\ : std_logic;
signal \N__74447\ : std_logic;
signal \N__74444\ : std_logic;
signal \N__74439\ : std_logic;
signal \N__74434\ : std_logic;
signal \N__74431\ : std_logic;
signal \N__74428\ : std_logic;
signal \N__74423\ : std_logic;
signal \N__74416\ : std_logic;
signal \N__74411\ : std_logic;
signal \N__74410\ : std_logic;
signal \N__74407\ : std_logic;
signal \N__74406\ : std_logic;
signal \N__74403\ : std_logic;
signal \N__74400\ : std_logic;
signal \N__74397\ : std_logic;
signal \N__74394\ : std_logic;
signal \N__74391\ : std_logic;
signal \N__74386\ : std_logic;
signal \N__74383\ : std_logic;
signal \N__74378\ : std_logic;
signal \N__74375\ : std_logic;
signal \N__74372\ : std_logic;
signal \N__74369\ : std_logic;
signal \N__74366\ : std_logic;
signal \N__74363\ : std_logic;
signal \N__74360\ : std_logic;
signal \N__74357\ : std_logic;
signal \N__74354\ : std_logic;
signal \N__74351\ : std_logic;
signal \N__74348\ : std_logic;
signal \N__74345\ : std_logic;
signal \N__74342\ : std_logic;
signal \N__74339\ : std_logic;
signal \N__74336\ : std_logic;
signal \N__74333\ : std_logic;
signal \N__74330\ : std_logic;
signal \N__74329\ : std_logic;
signal \N__74324\ : std_logic;
signal \N__74321\ : std_logic;
signal \N__74318\ : std_logic;
signal \N__74315\ : std_logic;
signal \N__74312\ : std_logic;
signal \N__74309\ : std_logic;
signal \N__74306\ : std_logic;
signal \N__74303\ : std_logic;
signal \N__74300\ : std_logic;
signal \N__74297\ : std_logic;
signal \N__74294\ : std_logic;
signal \N__74291\ : std_logic;
signal \N__74288\ : std_logic;
signal \N__74285\ : std_logic;
signal \N__74282\ : std_logic;
signal \N__74279\ : std_logic;
signal \N__74276\ : std_logic;
signal \N__74273\ : std_logic;
signal \N__74270\ : std_logic;
signal \N__74267\ : std_logic;
signal \N__74264\ : std_logic;
signal \N__74261\ : std_logic;
signal \N__74258\ : std_logic;
signal \N__74255\ : std_logic;
signal \N__74252\ : std_logic;
signal \N__74249\ : std_logic;
signal \N__74246\ : std_logic;
signal \N__74243\ : std_logic;
signal \N__74240\ : std_logic;
signal \N__74239\ : std_logic;
signal \N__74236\ : std_logic;
signal \N__74233\ : std_logic;
signal \N__74230\ : std_logic;
signal \N__74225\ : std_logic;
signal \N__74222\ : std_logic;
signal \N__74219\ : std_logic;
signal \N__74216\ : std_logic;
signal \N__74213\ : std_logic;
signal \N__74212\ : std_logic;
signal \N__74207\ : std_logic;
signal \N__74204\ : std_logic;
signal \N__74201\ : std_logic;
signal \N__74198\ : std_logic;
signal \N__74195\ : std_logic;
signal \N__74192\ : std_logic;
signal \N__74189\ : std_logic;
signal \N__74186\ : std_logic;
signal \N__74185\ : std_logic;
signal \N__74182\ : std_logic;
signal \N__74179\ : std_logic;
signal \N__74176\ : std_logic;
signal \N__74171\ : std_logic;
signal \N__74168\ : std_logic;
signal \N__74165\ : std_logic;
signal \N__74162\ : std_logic;
signal \N__74159\ : std_logic;
signal \N__74156\ : std_logic;
signal \N__74153\ : std_logic;
signal \N__74150\ : std_logic;
signal \N__74147\ : std_logic;
signal \N__74144\ : std_logic;
signal \N__74141\ : std_logic;
signal \N__74138\ : std_logic;
signal \N__74135\ : std_logic;
signal \N__74132\ : std_logic;
signal \N__74129\ : std_logic;
signal \N__74126\ : std_logic;
signal \N__74125\ : std_logic;
signal \N__74122\ : std_logic;
signal \N__74119\ : std_logic;
signal \N__74116\ : std_logic;
signal \N__74111\ : std_logic;
signal \N__74108\ : std_logic;
signal \N__74105\ : std_logic;
signal \N__74102\ : std_logic;
signal \N__74099\ : std_logic;
signal \N__74096\ : std_logic;
signal \N__74093\ : std_logic;
signal \N__74090\ : std_logic;
signal \N__74087\ : std_logic;
signal \N__74084\ : std_logic;
signal \N__74081\ : std_logic;
signal \N__74078\ : std_logic;
signal \N__74075\ : std_logic;
signal \N__74072\ : std_logic;
signal \N__74071\ : std_logic;
signal \N__74070\ : std_logic;
signal \N__74069\ : std_logic;
signal \N__74068\ : std_logic;
signal \N__74067\ : std_logic;
signal \N__74066\ : std_logic;
signal \N__74065\ : std_logic;
signal \N__74062\ : std_logic;
signal \N__74061\ : std_logic;
signal \N__74058\ : std_logic;
signal \N__74053\ : std_logic;
signal \N__74050\ : std_logic;
signal \N__74045\ : std_logic;
signal \N__74042\ : std_logic;
signal \N__74039\ : std_logic;
signal \N__74038\ : std_logic;
signal \N__74037\ : std_logic;
signal \N__74034\ : std_logic;
signal \N__74031\ : std_logic;
signal \N__74024\ : std_logic;
signal \N__74023\ : std_logic;
signal \N__74020\ : std_logic;
signal \N__74017\ : std_logic;
signal \N__74012\ : std_logic;
signal \N__74011\ : std_logic;
signal \N__74008\ : std_logic;
signal \N__74007\ : std_logic;
signal \N__74004\ : std_logic;
signal \N__74001\ : std_logic;
signal \N__73998\ : std_logic;
signal \N__73997\ : std_logic;
signal \N__73994\ : std_logic;
signal \N__73989\ : std_logic;
signal \N__73986\ : std_logic;
signal \N__73983\ : std_logic;
signal \N__73980\ : std_logic;
signal \N__73977\ : std_logic;
signal \N__73972\ : std_logic;
signal \N__73969\ : std_logic;
signal \N__73964\ : std_logic;
signal \N__73959\ : std_logic;
signal \N__73946\ : std_logic;
signal \N__73945\ : std_logic;
signal \N__73942\ : std_logic;
signal \N__73937\ : std_logic;
signal \N__73934\ : std_logic;
signal \N__73931\ : std_logic;
signal \N__73928\ : std_logic;
signal \N__73925\ : std_logic;
signal \N__73922\ : std_logic;
signal \N__73919\ : std_logic;
signal \N__73918\ : std_logic;
signal \N__73915\ : std_logic;
signal \N__73912\ : std_logic;
signal \N__73911\ : std_logic;
signal \N__73906\ : std_logic;
signal \N__73905\ : std_logic;
signal \N__73902\ : std_logic;
signal \N__73899\ : std_logic;
signal \N__73896\ : std_logic;
signal \N__73893\ : std_logic;
signal \N__73892\ : std_logic;
signal \N__73891\ : std_logic;
signal \N__73886\ : std_logic;
signal \N__73883\ : std_logic;
signal \N__73880\ : std_logic;
signal \N__73877\ : std_logic;
signal \N__73874\ : std_logic;
signal \N__73873\ : std_logic;
signal \N__73870\ : std_logic;
signal \N__73867\ : std_logic;
signal \N__73864\ : std_logic;
signal \N__73861\ : std_logic;
signal \N__73858\ : std_logic;
signal \N__73857\ : std_logic;
signal \N__73852\ : std_logic;
signal \N__73849\ : std_logic;
signal \N__73846\ : std_logic;
signal \N__73841\ : std_logic;
signal \N__73838\ : std_logic;
signal \N__73829\ : std_logic;
signal \N__73826\ : std_logic;
signal \N__73823\ : std_logic;
signal \N__73820\ : std_logic;
signal \N__73817\ : std_logic;
signal \N__73814\ : std_logic;
signal \N__73813\ : std_logic;
signal \N__73812\ : std_logic;
signal \N__73811\ : std_logic;
signal \N__73810\ : std_logic;
signal \N__73809\ : std_logic;
signal \N__73808\ : std_logic;
signal \N__73805\ : std_logic;
signal \N__73800\ : std_logic;
signal \N__73797\ : std_logic;
signal \N__73794\ : std_logic;
signal \N__73791\ : std_logic;
signal \N__73788\ : std_logic;
signal \N__73787\ : std_logic;
signal \N__73784\ : std_logic;
signal \N__73781\ : std_logic;
signal \N__73778\ : std_logic;
signal \N__73773\ : std_logic;
signal \N__73770\ : std_logic;
signal \N__73767\ : std_logic;
signal \N__73766\ : std_logic;
signal \N__73761\ : std_logic;
signal \N__73752\ : std_logic;
signal \N__73749\ : std_logic;
signal \N__73742\ : std_logic;
signal \N__73741\ : std_logic;
signal \N__73740\ : std_logic;
signal \N__73737\ : std_logic;
signal \N__73734\ : std_logic;
signal \N__73731\ : std_logic;
signal \N__73730\ : std_logic;
signal \N__73729\ : std_logic;
signal \N__73728\ : std_logic;
signal \N__73725\ : std_logic;
signal \N__73722\ : std_logic;
signal \N__73721\ : std_logic;
signal \N__73720\ : std_logic;
signal \N__73719\ : std_logic;
signal \N__73716\ : std_logic;
signal \N__73713\ : std_logic;
signal \N__73712\ : std_logic;
signal \N__73707\ : std_logic;
signal \N__73702\ : std_logic;
signal \N__73697\ : std_logic;
signal \N__73694\ : std_logic;
signal \N__73691\ : std_logic;
signal \N__73688\ : std_logic;
signal \N__73687\ : std_logic;
signal \N__73686\ : std_logic;
signal \N__73683\ : std_logic;
signal \N__73680\ : std_logic;
signal \N__73679\ : std_logic;
signal \N__73678\ : std_logic;
signal \N__73677\ : std_logic;
signal \N__73672\ : std_logic;
signal \N__73669\ : std_logic;
signal \N__73668\ : std_logic;
signal \N__73665\ : std_logic;
signal \N__73662\ : std_logic;
signal \N__73661\ : std_logic;
signal \N__73658\ : std_logic;
signal \N__73655\ : std_logic;
signal \N__73652\ : std_logic;
signal \N__73649\ : std_logic;
signal \N__73642\ : std_logic;
signal \N__73637\ : std_logic;
signal \N__73636\ : std_logic;
signal \N__73633\ : std_logic;
signal \N__73628\ : std_logic;
signal \N__73627\ : std_logic;
signal \N__73624\ : std_logic;
signal \N__73619\ : std_logic;
signal \N__73614\ : std_logic;
signal \N__73611\ : std_logic;
signal \N__73608\ : std_logic;
signal \N__73605\ : std_logic;
signal \N__73600\ : std_logic;
signal \N__73595\ : std_logic;
signal \N__73588\ : std_logic;
signal \N__73585\ : std_logic;
signal \N__73574\ : std_logic;
signal \N__73573\ : std_logic;
signal \N__73572\ : std_logic;
signal \N__73569\ : std_logic;
signal \N__73566\ : std_logic;
signal \N__73565\ : std_logic;
signal \N__73562\ : std_logic;
signal \N__73559\ : std_logic;
signal \N__73554\ : std_logic;
signal \N__73553\ : std_logic;
signal \N__73552\ : std_logic;
signal \N__73549\ : std_logic;
signal \N__73546\ : std_logic;
signal \N__73543\ : std_logic;
signal \N__73542\ : std_logic;
signal \N__73539\ : std_logic;
signal \N__73536\ : std_logic;
signal \N__73533\ : std_logic;
signal \N__73530\ : std_logic;
signal \N__73527\ : std_logic;
signal \N__73524\ : std_logic;
signal \N__73519\ : std_logic;
signal \N__73516\ : std_logic;
signal \N__73505\ : std_logic;
signal \N__73504\ : std_logic;
signal \N__73503\ : std_logic;
signal \N__73498\ : std_logic;
signal \N__73495\ : std_logic;
signal \N__73492\ : std_logic;
signal \N__73491\ : std_logic;
signal \N__73488\ : std_logic;
signal \N__73485\ : std_logic;
signal \N__73482\ : std_logic;
signal \N__73475\ : std_logic;
signal \N__73472\ : std_logic;
signal \N__73469\ : std_logic;
signal \N__73466\ : std_logic;
signal \N__73463\ : std_logic;
signal \N__73460\ : std_logic;
signal \N__73457\ : std_logic;
signal \N__73454\ : std_logic;
signal \N__73451\ : std_logic;
signal \N__73448\ : std_logic;
signal \N__73445\ : std_logic;
signal \N__73442\ : std_logic;
signal \N__73439\ : std_logic;
signal \N__73436\ : std_logic;
signal \N__73433\ : std_logic;
signal \N__73430\ : std_logic;
signal \N__73427\ : std_logic;
signal \N__73424\ : std_logic;
signal \N__73421\ : std_logic;
signal \N__73418\ : std_logic;
signal \N__73415\ : std_logic;
signal \N__73412\ : std_logic;
signal \N__73409\ : std_logic;
signal \N__73406\ : std_logic;
signal \N__73403\ : std_logic;
signal \N__73400\ : std_logic;
signal \N__73397\ : std_logic;
signal \N__73394\ : std_logic;
signal \N__73391\ : std_logic;
signal \N__73388\ : std_logic;
signal \N__73385\ : std_logic;
signal \N__73382\ : std_logic;
signal \N__73379\ : std_logic;
signal \N__73376\ : std_logic;
signal \N__73373\ : std_logic;
signal \N__73370\ : std_logic;
signal \N__73367\ : std_logic;
signal \N__73364\ : std_logic;
signal \N__73361\ : std_logic;
signal \N__73358\ : std_logic;
signal \N__73355\ : std_logic;
signal \N__73352\ : std_logic;
signal \N__73349\ : std_logic;
signal \N__73348\ : std_logic;
signal \N__73345\ : std_logic;
signal \N__73342\ : std_logic;
signal \N__73339\ : std_logic;
signal \N__73336\ : std_logic;
signal \N__73333\ : std_logic;
signal \N__73330\ : std_logic;
signal \N__73327\ : std_logic;
signal \N__73324\ : std_logic;
signal \N__73319\ : std_logic;
signal \N__73316\ : std_logic;
signal \N__73313\ : std_logic;
signal \N__73310\ : std_logic;
signal \N__73307\ : std_logic;
signal \N__73304\ : std_logic;
signal \N__73303\ : std_logic;
signal \N__73302\ : std_logic;
signal \N__73299\ : std_logic;
signal \N__73294\ : std_logic;
signal \N__73293\ : std_logic;
signal \N__73292\ : std_logic;
signal \N__73291\ : std_logic;
signal \N__73290\ : std_logic;
signal \N__73287\ : std_logic;
signal \N__73286\ : std_logic;
signal \N__73283\ : std_logic;
signal \N__73282\ : std_logic;
signal \N__73281\ : std_logic;
signal \N__73280\ : std_logic;
signal \N__73279\ : std_logic;
signal \N__73278\ : std_logic;
signal \N__73277\ : std_logic;
signal \N__73276\ : std_logic;
signal \N__73275\ : std_logic;
signal \N__73274\ : std_logic;
signal \N__73273\ : std_logic;
signal \N__73272\ : std_logic;
signal \N__73271\ : std_logic;
signal \N__73270\ : std_logic;
signal \N__73269\ : std_logic;
signal \N__73268\ : std_logic;
signal \N__73267\ : std_logic;
signal \N__73266\ : std_logic;
signal \N__73265\ : std_logic;
signal \N__73264\ : std_logic;
signal \N__73263\ : std_logic;
signal \N__73262\ : std_logic;
signal \N__73261\ : std_logic;
signal \N__73260\ : std_logic;
signal \N__73259\ : std_logic;
signal \N__73258\ : std_logic;
signal \N__73257\ : std_logic;
signal \N__73256\ : std_logic;
signal \N__73255\ : std_logic;
signal \N__73254\ : std_logic;
signal \N__73253\ : std_logic;
signal \N__73252\ : std_logic;
signal \N__73251\ : std_logic;
signal \N__73250\ : std_logic;
signal \N__73249\ : std_logic;
signal \N__73248\ : std_logic;
signal \N__73247\ : std_logic;
signal \N__73246\ : std_logic;
signal \N__73245\ : std_logic;
signal \N__73244\ : std_logic;
signal \N__73243\ : std_logic;
signal \N__73242\ : std_logic;
signal \N__73241\ : std_logic;
signal \N__73240\ : std_logic;
signal \N__73239\ : std_logic;
signal \N__73238\ : std_logic;
signal \N__73237\ : std_logic;
signal \N__73236\ : std_logic;
signal \N__73235\ : std_logic;
signal \N__73234\ : std_logic;
signal \N__73233\ : std_logic;
signal \N__73232\ : std_logic;
signal \N__73231\ : std_logic;
signal \N__73230\ : std_logic;
signal \N__73229\ : std_logic;
signal \N__73228\ : std_logic;
signal \N__73227\ : std_logic;
signal \N__73226\ : std_logic;
signal \N__73225\ : std_logic;
signal \N__73224\ : std_logic;
signal \N__73223\ : std_logic;
signal \N__73222\ : std_logic;
signal \N__73221\ : std_logic;
signal \N__73220\ : std_logic;
signal \N__73219\ : std_logic;
signal \N__73218\ : std_logic;
signal \N__73217\ : std_logic;
signal \N__73216\ : std_logic;
signal \N__73215\ : std_logic;
signal \N__73214\ : std_logic;
signal \N__73213\ : std_logic;
signal \N__73212\ : std_logic;
signal \N__73211\ : std_logic;
signal \N__73210\ : std_logic;
signal \N__73209\ : std_logic;
signal \N__73208\ : std_logic;
signal \N__73207\ : std_logic;
signal \N__73206\ : std_logic;
signal \N__73205\ : std_logic;
signal \N__73204\ : std_logic;
signal \N__73203\ : std_logic;
signal \N__73202\ : std_logic;
signal \N__73201\ : std_logic;
signal \N__73200\ : std_logic;
signal \N__73199\ : std_logic;
signal \N__73198\ : std_logic;
signal \N__73197\ : std_logic;
signal \N__73196\ : std_logic;
signal \N__73195\ : std_logic;
signal \N__73194\ : std_logic;
signal \N__73193\ : std_logic;
signal \N__73192\ : std_logic;
signal \N__73191\ : std_logic;
signal \N__73190\ : std_logic;
signal \N__73189\ : std_logic;
signal \N__73188\ : std_logic;
signal \N__73187\ : std_logic;
signal \N__73186\ : std_logic;
signal \N__73185\ : std_logic;
signal \N__73184\ : std_logic;
signal \N__73183\ : std_logic;
signal \N__73182\ : std_logic;
signal \N__73181\ : std_logic;
signal \N__73180\ : std_logic;
signal \N__73179\ : std_logic;
signal \N__73178\ : std_logic;
signal \N__73177\ : std_logic;
signal \N__73176\ : std_logic;
signal \N__73175\ : std_logic;
signal \N__73174\ : std_logic;
signal \N__73173\ : std_logic;
signal \N__73172\ : std_logic;
signal \N__73171\ : std_logic;
signal \N__73170\ : std_logic;
signal \N__73169\ : std_logic;
signal \N__73168\ : std_logic;
signal \N__73167\ : std_logic;
signal \N__73166\ : std_logic;
signal \N__73165\ : std_logic;
signal \N__73164\ : std_logic;
signal \N__73163\ : std_logic;
signal \N__73162\ : std_logic;
signal \N__73161\ : std_logic;
signal \N__73160\ : std_logic;
signal \N__73159\ : std_logic;
signal \N__73158\ : std_logic;
signal \N__73157\ : std_logic;
signal \N__73156\ : std_logic;
signal \N__73155\ : std_logic;
signal \N__73154\ : std_logic;
signal \N__73153\ : std_logic;
signal \N__73152\ : std_logic;
signal \N__73151\ : std_logic;
signal \N__73150\ : std_logic;
signal \N__73149\ : std_logic;
signal \N__73148\ : std_logic;
signal \N__73147\ : std_logic;
signal \N__73146\ : std_logic;
signal \N__73145\ : std_logic;
signal \N__73144\ : std_logic;
signal \N__73143\ : std_logic;
signal \N__73142\ : std_logic;
signal \N__73141\ : std_logic;
signal \N__73140\ : std_logic;
signal \N__73139\ : std_logic;
signal \N__73138\ : std_logic;
signal \N__72833\ : std_logic;
signal \N__72830\ : std_logic;
signal \N__72827\ : std_logic;
signal \N__72824\ : std_logic;
signal \N__72821\ : std_logic;
signal \N__72818\ : std_logic;
signal \N__72815\ : std_logic;
signal \N__72812\ : std_logic;
signal \N__72809\ : std_logic;
signal \N__72806\ : std_logic;
signal \N__72803\ : std_logic;
signal \N__72800\ : std_logic;
signal \N__72797\ : std_logic;
signal \N__72794\ : std_logic;
signal \N__72791\ : std_logic;
signal \N__72790\ : std_logic;
signal \N__72789\ : std_logic;
signal \N__72786\ : std_logic;
signal \N__72785\ : std_logic;
signal \N__72784\ : std_logic;
signal \N__72781\ : std_logic;
signal \N__72778\ : std_logic;
signal \N__72777\ : std_logic;
signal \N__72776\ : std_logic;
signal \N__72775\ : std_logic;
signal \N__72774\ : std_logic;
signal \N__72773\ : std_logic;
signal \N__72772\ : std_logic;
signal \N__72771\ : std_logic;
signal \N__72770\ : std_logic;
signal \N__72769\ : std_logic;
signal \N__72768\ : std_logic;
signal \N__72761\ : std_logic;
signal \N__72752\ : std_logic;
signal \N__72749\ : std_logic;
signal \N__72746\ : std_logic;
signal \N__72743\ : std_logic;
signal \N__72742\ : std_logic;
signal \N__72741\ : std_logic;
signal \N__72738\ : std_logic;
signal \N__72737\ : std_logic;
signal \N__72732\ : std_logic;
signal \N__72731\ : std_logic;
signal \N__72730\ : std_logic;
signal \N__72729\ : std_logic;
signal \N__72728\ : std_logic;
signal \N__72727\ : std_logic;
signal \N__72726\ : std_logic;
signal \N__72725\ : std_logic;
signal \N__72724\ : std_logic;
signal \N__72723\ : std_logic;
signal \N__72722\ : std_logic;
signal \N__72721\ : std_logic;
signal \N__72720\ : std_logic;
signal \N__72717\ : std_logic;
signal \N__72714\ : std_logic;
signal \N__72713\ : std_logic;
signal \N__72712\ : std_logic;
signal \N__72707\ : std_logic;
signal \N__72704\ : std_logic;
signal \N__72699\ : std_logic;
signal \N__72698\ : std_logic;
signal \N__72697\ : std_logic;
signal \N__72696\ : std_logic;
signal \N__72695\ : std_logic;
signal \N__72694\ : std_logic;
signal \N__72693\ : std_logic;
signal \N__72692\ : std_logic;
signal \N__72691\ : std_logic;
signal \N__72690\ : std_logic;
signal \N__72689\ : std_logic;
signal \N__72688\ : std_logic;
signal \N__72685\ : std_logic;
signal \N__72684\ : std_logic;
signal \N__72683\ : std_logic;
signal \N__72682\ : std_logic;
signal \N__72681\ : std_logic;
signal \N__72676\ : std_logic;
signal \N__72673\ : std_logic;
signal \N__72672\ : std_logic;
signal \N__72669\ : std_logic;
signal \N__72666\ : std_logic;
signal \N__72657\ : std_logic;
signal \N__72656\ : std_logic;
signal \N__72655\ : std_logic;
signal \N__72652\ : std_logic;
signal \N__72649\ : std_logic;
signal \N__72648\ : std_logic;
signal \N__72637\ : std_logic;
signal \N__72630\ : std_logic;
signal \N__72627\ : std_logic;
signal \N__72626\ : std_logic;
signal \N__72619\ : std_logic;
signal \N__72618\ : std_logic;
signal \N__72615\ : std_logic;
signal \N__72612\ : std_logic;
signal \N__72609\ : std_logic;
signal \N__72608\ : std_logic;
signal \N__72607\ : std_logic;
signal \N__72606\ : std_logic;
signal \N__72603\ : std_logic;
signal \N__72600\ : std_logic;
signal \N__72597\ : std_logic;
signal \N__72588\ : std_logic;
signal \N__72583\ : std_logic;
signal \N__72580\ : std_logic;
signal \N__72577\ : std_logic;
signal \N__72572\ : std_logic;
signal \N__72567\ : std_logic;
signal \N__72564\ : std_logic;
signal \N__72563\ : std_logic;
signal \N__72560\ : std_logic;
signal \N__72557\ : std_logic;
signal \N__72554\ : std_logic;
signal \N__72549\ : std_logic;
signal \N__72546\ : std_logic;
signal \N__72541\ : std_logic;
signal \N__72538\ : std_logic;
signal \N__72535\ : std_logic;
signal \N__72532\ : std_logic;
signal \N__72529\ : std_logic;
signal \N__72526\ : std_logic;
signal \N__72523\ : std_logic;
signal \N__72520\ : std_logic;
signal \N__72515\ : std_logic;
signal \N__72512\ : std_logic;
signal \N__72511\ : std_logic;
signal \N__72508\ : std_logic;
signal \N__72505\ : std_logic;
signal \N__72504\ : std_logic;
signal \N__72503\ : std_logic;
signal \N__72500\ : std_logic;
signal \N__72495\ : std_logic;
signal \N__72490\ : std_logic;
signal \N__72485\ : std_logic;
signal \N__72480\ : std_logic;
signal \N__72475\ : std_logic;
signal \N__72470\ : std_logic;
signal \N__72461\ : std_logic;
signal \N__72454\ : std_logic;
signal \N__72451\ : std_logic;
signal \N__72446\ : std_logic;
signal \N__72439\ : std_logic;
signal \N__72436\ : std_logic;
signal \N__72433\ : std_logic;
signal \N__72430\ : std_logic;
signal \N__72427\ : std_logic;
signal \N__72424\ : std_logic;
signal \N__72415\ : std_logic;
signal \N__72404\ : std_logic;
signal \N__72383\ : std_logic;
signal \N__72380\ : std_logic;
signal \N__72377\ : std_logic;
signal \N__72376\ : std_logic;
signal \N__72373\ : std_logic;
signal \N__72370\ : std_logic;
signal \N__72367\ : std_logic;
signal \N__72364\ : std_logic;
signal \N__72361\ : std_logic;
signal \N__72358\ : std_logic;
signal \N__72353\ : std_logic;
signal \N__72352\ : std_logic;
signal \N__72349\ : std_logic;
signal \N__72348\ : std_logic;
signal \N__72345\ : std_logic;
signal \N__72342\ : std_logic;
signal \N__72339\ : std_logic;
signal \N__72336\ : std_logic;
signal \N__72331\ : std_logic;
signal \N__72328\ : std_logic;
signal \N__72325\ : std_logic;
signal \N__72320\ : std_logic;
signal \N__72319\ : std_logic;
signal \N__72318\ : std_logic;
signal \N__72317\ : std_logic;
signal \N__72316\ : std_logic;
signal \N__72315\ : std_logic;
signal \N__72312\ : std_logic;
signal \N__72311\ : std_logic;
signal \N__72308\ : std_logic;
signal \N__72307\ : std_logic;
signal \N__72306\ : std_logic;
signal \N__72305\ : std_logic;
signal \N__72304\ : std_logic;
signal \N__72301\ : std_logic;
signal \N__72300\ : std_logic;
signal \N__72299\ : std_logic;
signal \N__72298\ : std_logic;
signal \N__72297\ : std_logic;
signal \N__72294\ : std_logic;
signal \N__72293\ : std_logic;
signal \N__72290\ : std_logic;
signal \N__72289\ : std_logic;
signal \N__72288\ : std_logic;
signal \N__72285\ : std_logic;
signal \N__72284\ : std_logic;
signal \N__72281\ : std_logic;
signal \N__72274\ : std_logic;
signal \N__72273\ : std_logic;
signal \N__72272\ : std_logic;
signal \N__72271\ : std_logic;
signal \N__72268\ : std_logic;
signal \N__72265\ : std_logic;
signal \N__72264\ : std_logic;
signal \N__72263\ : std_logic;
signal \N__72262\ : std_logic;
signal \N__72261\ : std_logic;
signal \N__72260\ : std_logic;
signal \N__72257\ : std_logic;
signal \N__72256\ : std_logic;
signal \N__72253\ : std_logic;
signal \N__72252\ : std_logic;
signal \N__72251\ : std_logic;
signal \N__72250\ : std_logic;
signal \N__72249\ : std_logic;
signal \N__72248\ : std_logic;
signal \N__72247\ : std_logic;
signal \N__72244\ : std_logic;
signal \N__72239\ : std_logic;
signal \N__72236\ : std_logic;
signal \N__72231\ : std_logic;
signal \N__72228\ : std_logic;
signal \N__72227\ : std_logic;
signal \N__72226\ : std_logic;
signal \N__72225\ : std_logic;
signal \N__72224\ : std_logic;
signal \N__72223\ : std_logic;
signal \N__72222\ : std_logic;
signal \N__72221\ : std_logic;
signal \N__72220\ : std_logic;
signal \N__72217\ : std_logic;
signal \N__72214\ : std_logic;
signal \N__72213\ : std_logic;
signal \N__72212\ : std_logic;
signal \N__72209\ : std_logic;
signal \N__72206\ : std_logic;
signal \N__72201\ : std_logic;
signal \N__72198\ : std_logic;
signal \N__72195\ : std_logic;
signal \N__72194\ : std_logic;
signal \N__72193\ : std_logic;
signal \N__72192\ : std_logic;
signal \N__72191\ : std_logic;
signal \N__72190\ : std_logic;
signal \N__72189\ : std_logic;
signal \N__72188\ : std_logic;
signal \N__72185\ : std_logic;
signal \N__72182\ : std_logic;
signal \N__72181\ : std_logic;
signal \N__72180\ : std_logic;
signal \N__72179\ : std_logic;
signal \N__72178\ : std_logic;
signal \N__72177\ : std_logic;
signal \N__72176\ : std_logic;
signal \N__72171\ : std_logic;
signal \N__72166\ : std_logic;
signal \N__72161\ : std_logic;
signal \N__72158\ : std_logic;
signal \N__72155\ : std_logic;
signal \N__72152\ : std_logic;
signal \N__72149\ : std_logic;
signal \N__72146\ : std_logic;
signal \N__72141\ : std_logic;
signal \N__72140\ : std_logic;
signal \N__72137\ : std_logic;
signal \N__72134\ : std_logic;
signal \N__72133\ : std_logic;
signal \N__72132\ : std_logic;
signal \N__72131\ : std_logic;
signal \N__72130\ : std_logic;
signal \N__72129\ : std_logic;
signal \N__72128\ : std_logic;
signal \N__72123\ : std_logic;
signal \N__72118\ : std_logic;
signal \N__72115\ : std_logic;
signal \N__72110\ : std_logic;
signal \N__72105\ : std_logic;
signal \N__72104\ : std_logic;
signal \N__72103\ : std_logic;
signal \N__72102\ : std_logic;
signal \N__72101\ : std_logic;
signal \N__72100\ : std_logic;
signal \N__72097\ : std_logic;
signal \N__72092\ : std_logic;
signal \N__72081\ : std_logic;
signal \N__72078\ : std_logic;
signal \N__72075\ : std_logic;
signal \N__72068\ : std_logic;
signal \N__72061\ : std_logic;
signal \N__72052\ : std_logic;
signal \N__72047\ : std_logic;
signal \N__72044\ : std_logic;
signal \N__72033\ : std_logic;
signal \N__72026\ : std_logic;
signal \N__72013\ : std_logic;
signal \N__72010\ : std_logic;
signal \N__72009\ : std_logic;
signal \N__72008\ : std_logic;
signal \N__72005\ : std_logic;
signal \N__72002\ : std_logic;
signal \N__71997\ : std_logic;
signal \N__71994\ : std_logic;
signal \N__71987\ : std_logic;
signal \N__71976\ : std_logic;
signal \N__71973\ : std_logic;
signal \N__71968\ : std_logic;
signal \N__71963\ : std_logic;
signal \N__71960\ : std_logic;
signal \N__71951\ : std_logic;
signal \N__71948\ : std_logic;
signal \N__71935\ : std_logic;
signal \N__71932\ : std_logic;
signal \N__71925\ : std_logic;
signal \N__71922\ : std_logic;
signal \N__71915\ : std_logic;
signal \N__71910\ : std_logic;
signal \N__71895\ : std_logic;
signal \N__71892\ : std_logic;
signal \N__71879\ : std_logic;
signal \N__71876\ : std_logic;
signal \N__71875\ : std_logic;
signal \N__71874\ : std_logic;
signal \N__71873\ : std_logic;
signal \N__71872\ : std_logic;
signal \N__71871\ : std_logic;
signal \N__71870\ : std_logic;
signal \N__71869\ : std_logic;
signal \N__71868\ : std_logic;
signal \N__71867\ : std_logic;
signal \N__71866\ : std_logic;
signal \N__71863\ : std_logic;
signal \N__71860\ : std_logic;
signal \N__71855\ : std_logic;
signal \N__71854\ : std_logic;
signal \N__71853\ : std_logic;
signal \N__71852\ : std_logic;
signal \N__71849\ : std_logic;
signal \N__71842\ : std_logic;
signal \N__71835\ : std_logic;
signal \N__71832\ : std_logic;
signal \N__71831\ : std_logic;
signal \N__71830\ : std_logic;
signal \N__71829\ : std_logic;
signal \N__71828\ : std_logic;
signal \N__71827\ : std_logic;
signal \N__71826\ : std_logic;
signal \N__71825\ : std_logic;
signal \N__71824\ : std_logic;
signal \N__71823\ : std_logic;
signal \N__71822\ : std_logic;
signal \N__71821\ : std_logic;
signal \N__71820\ : std_logic;
signal \N__71819\ : std_logic;
signal \N__71816\ : std_logic;
signal \N__71813\ : std_logic;
signal \N__71810\ : std_logic;
signal \N__71807\ : std_logic;
signal \N__71806\ : std_logic;
signal \N__71805\ : std_logic;
signal \N__71804\ : std_logic;
signal \N__71803\ : std_logic;
signal \N__71802\ : std_logic;
signal \N__71799\ : std_logic;
signal \N__71792\ : std_logic;
signal \N__71789\ : std_logic;
signal \N__71786\ : std_logic;
signal \N__71783\ : std_logic;
signal \N__71776\ : std_logic;
signal \N__71765\ : std_logic;
signal \N__71762\ : std_logic;
signal \N__71759\ : std_logic;
signal \N__71758\ : std_logic;
signal \N__71755\ : std_logic;
signal \N__71752\ : std_logic;
signal \N__71749\ : std_logic;
signal \N__71746\ : std_logic;
signal \N__71745\ : std_logic;
signal \N__71742\ : std_logic;
signal \N__71739\ : std_logic;
signal \N__71730\ : std_logic;
signal \N__71727\ : std_logic;
signal \N__71722\ : std_logic;
signal \N__71715\ : std_logic;
signal \N__71712\ : std_logic;
signal \N__71709\ : std_logic;
signal \N__71706\ : std_logic;
signal \N__71701\ : std_logic;
signal \N__71698\ : std_logic;
signal \N__71693\ : std_logic;
signal \N__71690\ : std_logic;
signal \N__71683\ : std_logic;
signal \N__71676\ : std_logic;
signal \N__71657\ : std_logic;
signal \N__71654\ : std_logic;
signal \N__71651\ : std_logic;
signal \N__71648\ : std_logic;
signal \N__71645\ : std_logic;
signal \N__71642\ : std_logic;
signal \N__71639\ : std_logic;
signal \N__71636\ : std_logic;
signal \N__71633\ : std_logic;
signal \N__71630\ : std_logic;
signal \N__71627\ : std_logic;
signal \N__71624\ : std_logic;
signal \N__71621\ : std_logic;
signal \N__71618\ : std_logic;
signal \N__71615\ : std_logic;
signal \N__71612\ : std_logic;
signal \N__71609\ : std_logic;
signal \N__71606\ : std_logic;
signal \N__71603\ : std_logic;
signal \N__71600\ : std_logic;
signal \N__71597\ : std_logic;
signal \N__71594\ : std_logic;
signal \N__71591\ : std_logic;
signal \N__71588\ : std_logic;
signal \N__71585\ : std_logic;
signal \N__71582\ : std_logic;
signal \N__71579\ : std_logic;
signal \N__71578\ : std_logic;
signal \N__71573\ : std_logic;
signal \N__71570\ : std_logic;
signal \N__71567\ : std_logic;
signal \N__71564\ : std_logic;
signal \N__71561\ : std_logic;
signal \N__71558\ : std_logic;
signal \N__71555\ : std_logic;
signal \N__71554\ : std_logic;
signal \N__71553\ : std_logic;
signal \N__71550\ : std_logic;
signal \N__71547\ : std_logic;
signal \N__71544\ : std_logic;
signal \N__71539\ : std_logic;
signal \N__71536\ : std_logic;
signal \N__71533\ : std_logic;
signal \N__71530\ : std_logic;
signal \N__71527\ : std_logic;
signal \N__71522\ : std_logic;
signal \N__71519\ : std_logic;
signal \N__71516\ : std_logic;
signal \N__71515\ : std_logic;
signal \N__71512\ : std_logic;
signal \N__71509\ : std_logic;
signal \N__71504\ : std_logic;
signal \N__71501\ : std_logic;
signal \N__71500\ : std_logic;
signal \N__71495\ : std_logic;
signal \N__71492\ : std_logic;
signal \N__71491\ : std_logic;
signal \N__71490\ : std_logic;
signal \N__71487\ : std_logic;
signal \N__71484\ : std_logic;
signal \N__71481\ : std_logic;
signal \N__71478\ : std_logic;
signal \N__71471\ : std_logic;
signal \N__71470\ : std_logic;
signal \N__71469\ : std_logic;
signal \N__71468\ : std_logic;
signal \N__71467\ : std_logic;
signal \N__71464\ : std_logic;
signal \N__71463\ : std_logic;
signal \N__71460\ : std_logic;
signal \N__71455\ : std_logic;
signal \N__71454\ : std_logic;
signal \N__71453\ : std_logic;
signal \N__71452\ : std_logic;
signal \N__71451\ : std_logic;
signal \N__71450\ : std_logic;
signal \N__71449\ : std_logic;
signal \N__71448\ : std_logic;
signal \N__71445\ : std_logic;
signal \N__71442\ : std_logic;
signal \N__71441\ : std_logic;
signal \N__71440\ : std_logic;
signal \N__71437\ : std_logic;
signal \N__71436\ : std_logic;
signal \N__71435\ : std_logic;
signal \N__71432\ : std_logic;
signal \N__71429\ : std_logic;
signal \N__71426\ : std_logic;
signal \N__71425\ : std_logic;
signal \N__71424\ : std_logic;
signal \N__71423\ : std_logic;
signal \N__71418\ : std_logic;
signal \N__71411\ : std_logic;
signal \N__71410\ : std_logic;
signal \N__71407\ : std_logic;
signal \N__71402\ : std_logic;
signal \N__71401\ : std_logic;
signal \N__71400\ : std_logic;
signal \N__71399\ : std_logic;
signal \N__71396\ : std_logic;
signal \N__71395\ : std_logic;
signal \N__71394\ : std_logic;
signal \N__71391\ : std_logic;
signal \N__71388\ : std_logic;
signal \N__71385\ : std_logic;
signal \N__71384\ : std_logic;
signal \N__71381\ : std_logic;
signal \N__71380\ : std_logic;
signal \N__71377\ : std_logic;
signal \N__71372\ : std_logic;
signal \N__71367\ : std_logic;
signal \N__71364\ : std_logic;
signal \N__71361\ : std_logic;
signal \N__71358\ : std_logic;
signal \N__71353\ : std_logic;
signal \N__71350\ : std_logic;
signal \N__71347\ : std_logic;
signal \N__71344\ : std_logic;
signal \N__71341\ : std_logic;
signal \N__71338\ : std_logic;
signal \N__71333\ : std_logic;
signal \N__71330\ : std_logic;
signal \N__71327\ : std_logic;
signal \N__71324\ : std_logic;
signal \N__71321\ : std_logic;
signal \N__71320\ : std_logic;
signal \N__71315\ : std_logic;
signal \N__71314\ : std_logic;
signal \N__71309\ : std_logic;
signal \N__71304\ : std_logic;
signal \N__71297\ : std_logic;
signal \N__71292\ : std_logic;
signal \N__71289\ : std_logic;
signal \N__71282\ : std_logic;
signal \N__71279\ : std_logic;
signal \N__71274\ : std_logic;
signal \N__71269\ : std_logic;
signal \N__71266\ : std_logic;
signal \N__71263\ : std_logic;
signal \N__71260\ : std_logic;
signal \N__71257\ : std_logic;
signal \N__71254\ : std_logic;
signal \N__71251\ : std_logic;
signal \N__71248\ : std_logic;
signal \N__71245\ : std_logic;
signal \N__71236\ : std_logic;
signal \N__71219\ : std_logic;
signal \N__71216\ : std_logic;
signal \N__71215\ : std_logic;
signal \N__71214\ : std_logic;
signal \N__71213\ : std_logic;
signal \N__71212\ : std_logic;
signal \N__71211\ : std_logic;
signal \N__71208\ : std_logic;
signal \N__71207\ : std_logic;
signal \N__71204\ : std_logic;
signal \N__71201\ : std_logic;
signal \N__71200\ : std_logic;
signal \N__71199\ : std_logic;
signal \N__71198\ : std_logic;
signal \N__71197\ : std_logic;
signal \N__71194\ : std_logic;
signal \N__71193\ : std_logic;
signal \N__71190\ : std_logic;
signal \N__71189\ : std_logic;
signal \N__71186\ : std_logic;
signal \N__71183\ : std_logic;
signal \N__71180\ : std_logic;
signal \N__71177\ : std_logic;
signal \N__71176\ : std_logic;
signal \N__71173\ : std_logic;
signal \N__71170\ : std_logic;
signal \N__71167\ : std_logic;
signal \N__71164\ : std_logic;
signal \N__71163\ : std_logic;
signal \N__71160\ : std_logic;
signal \N__71157\ : std_logic;
signal \N__71154\ : std_logic;
signal \N__71151\ : std_logic;
signal \N__71148\ : std_logic;
signal \N__71145\ : std_logic;
signal \N__71140\ : std_logic;
signal \N__71137\ : std_logic;
signal \N__71134\ : std_logic;
signal \N__71131\ : std_logic;
signal \N__71128\ : std_logic;
signal \N__71125\ : std_logic;
signal \N__71122\ : std_logic;
signal \N__71119\ : std_logic;
signal \N__71116\ : std_logic;
signal \N__71113\ : std_logic;
signal \N__71110\ : std_logic;
signal \N__71105\ : std_logic;
signal \N__71102\ : std_logic;
signal \N__71097\ : std_logic;
signal \N__71094\ : std_logic;
signal \N__71089\ : std_logic;
signal \N__71084\ : std_logic;
signal \N__71081\ : std_logic;
signal \N__71076\ : std_logic;
signal \N__71071\ : std_logic;
signal \N__71066\ : std_logic;
signal \N__71063\ : std_logic;
signal \N__71060\ : std_logic;
signal \N__71057\ : std_logic;
signal \N__71052\ : std_logic;
signal \N__71049\ : std_logic;
signal \N__71046\ : std_logic;
signal \N__71043\ : std_logic;
signal \N__71038\ : std_logic;
signal \N__71035\ : std_logic;
signal \N__71030\ : std_logic;
signal \N__71021\ : std_logic;
signal \N__71020\ : std_logic;
signal \N__71019\ : std_logic;
signal \N__71012\ : std_logic;
signal \N__71009\ : std_logic;
signal \N__71008\ : std_logic;
signal \N__71007\ : std_logic;
signal \N__71006\ : std_logic;
signal \N__70997\ : std_logic;
signal \N__70994\ : std_logic;
signal \N__70993\ : std_logic;
signal \N__70990\ : std_logic;
signal \N__70987\ : std_logic;
signal \N__70986\ : std_logic;
signal \N__70983\ : std_logic;
signal \N__70980\ : std_logic;
signal \N__70977\ : std_logic;
signal \N__70974\ : std_logic;
signal \N__70971\ : std_logic;
signal \N__70968\ : std_logic;
signal \N__70965\ : std_logic;
signal \N__70962\ : std_logic;
signal \N__70959\ : std_logic;
signal \N__70956\ : std_logic;
signal \N__70953\ : std_logic;
signal \N__70948\ : std_logic;
signal \N__70943\ : std_logic;
signal \N__70942\ : std_logic;
signal \N__70941\ : std_logic;
signal \N__70940\ : std_logic;
signal \N__70937\ : std_logic;
signal \N__70936\ : std_logic;
signal \N__70935\ : std_logic;
signal \N__70932\ : std_logic;
signal \N__70931\ : std_logic;
signal \N__70922\ : std_logic;
signal \N__70915\ : std_logic;
signal \N__70914\ : std_logic;
signal \N__70913\ : std_logic;
signal \N__70908\ : std_logic;
signal \N__70905\ : std_logic;
signal \N__70902\ : std_logic;
signal \N__70897\ : std_logic;
signal \N__70892\ : std_logic;
signal \N__70891\ : std_logic;
signal \N__70890\ : std_logic;
signal \N__70889\ : std_logic;
signal \N__70888\ : std_logic;
signal \N__70887\ : std_logic;
signal \N__70884\ : std_logic;
signal \N__70883\ : std_logic;
signal \N__70882\ : std_logic;
signal \N__70875\ : std_logic;
signal \N__70866\ : std_logic;
signal \N__70865\ : std_logic;
signal \N__70862\ : std_logic;
signal \N__70859\ : std_logic;
signal \N__70856\ : std_logic;
signal \N__70853\ : std_logic;
signal \N__70844\ : std_logic;
signal \N__70841\ : std_logic;
signal \N__70838\ : std_logic;
signal \N__70835\ : std_logic;
signal \N__70832\ : std_logic;
signal \N__70829\ : std_logic;
signal \N__70828\ : std_logic;
signal \N__70825\ : std_logic;
signal \N__70822\ : std_logic;
signal \N__70819\ : std_logic;
signal \N__70816\ : std_logic;
signal \N__70815\ : std_logic;
signal \N__70812\ : std_logic;
signal \N__70809\ : std_logic;
signal \N__70806\ : std_logic;
signal \N__70799\ : std_logic;
signal \N__70798\ : std_logic;
signal \N__70797\ : std_logic;
signal \N__70796\ : std_logic;
signal \N__70795\ : std_logic;
signal \N__70794\ : std_logic;
signal \N__70791\ : std_logic;
signal \N__70790\ : std_logic;
signal \N__70789\ : std_logic;
signal \N__70788\ : std_logic;
signal \N__70787\ : std_logic;
signal \N__70786\ : std_logic;
signal \N__70785\ : std_logic;
signal \N__70782\ : std_logic;
signal \N__70779\ : std_logic;
signal \N__70776\ : std_logic;
signal \N__70773\ : std_logic;
signal \N__70770\ : std_logic;
signal \N__70767\ : std_logic;
signal \N__70766\ : std_logic;
signal \N__70765\ : std_logic;
signal \N__70764\ : std_logic;
signal \N__70763\ : std_logic;
signal \N__70762\ : std_logic;
signal \N__70761\ : std_logic;
signal \N__70760\ : std_logic;
signal \N__70759\ : std_logic;
signal \N__70758\ : std_logic;
signal \N__70757\ : std_logic;
signal \N__70756\ : std_logic;
signal \N__70755\ : std_logic;
signal \N__70754\ : std_logic;
signal \N__70751\ : std_logic;
signal \N__70746\ : std_logic;
signal \N__70733\ : std_logic;
signal \N__70730\ : std_logic;
signal \N__70727\ : std_logic;
signal \N__70724\ : std_logic;
signal \N__70723\ : std_logic;
signal \N__70722\ : std_logic;
signal \N__70721\ : std_logic;
signal \N__70718\ : std_logic;
signal \N__70715\ : std_logic;
signal \N__70712\ : std_logic;
signal \N__70711\ : std_logic;
signal \N__70710\ : std_logic;
signal \N__70709\ : std_logic;
signal \N__70708\ : std_logic;
signal \N__70703\ : std_logic;
signal \N__70700\ : std_logic;
signal \N__70693\ : std_logic;
signal \N__70690\ : std_logic;
signal \N__70683\ : std_logic;
signal \N__70678\ : std_logic;
signal \N__70671\ : std_logic;
signal \N__70668\ : std_logic;
signal \N__70661\ : std_logic;
signal \N__70646\ : std_logic;
signal \N__70643\ : std_logic;
signal \N__70640\ : std_logic;
signal \N__70631\ : std_logic;
signal \N__70626\ : std_logic;
signal \N__70613\ : std_logic;
signal \N__70610\ : std_logic;
signal \N__70607\ : std_logic;
signal \N__70604\ : std_logic;
signal \N__70603\ : std_logic;
signal \N__70600\ : std_logic;
signal \N__70597\ : std_logic;
signal \N__70594\ : std_logic;
signal \N__70591\ : std_logic;
signal \N__70586\ : std_logic;
signal \N__70585\ : std_logic;
signal \N__70582\ : std_logic;
signal \N__70579\ : std_logic;
signal \N__70576\ : std_logic;
signal \N__70573\ : std_logic;
signal \N__70570\ : std_logic;
signal \N__70567\ : std_logic;
signal \N__70564\ : std_logic;
signal \N__70561\ : std_logic;
signal \N__70556\ : std_logic;
signal \N__70553\ : std_logic;
signal \N__70552\ : std_logic;
signal \N__70551\ : std_logic;
signal \N__70550\ : std_logic;
signal \N__70549\ : std_logic;
signal \N__70548\ : std_logic;
signal \N__70545\ : std_logic;
signal \N__70544\ : std_logic;
signal \N__70543\ : std_logic;
signal \N__70542\ : std_logic;
signal \N__70541\ : std_logic;
signal \N__70540\ : std_logic;
signal \N__70539\ : std_logic;
signal \N__70536\ : std_logic;
signal \N__70535\ : std_logic;
signal \N__70528\ : std_logic;
signal \N__70527\ : std_logic;
signal \N__70526\ : std_logic;
signal \N__70525\ : std_logic;
signal \N__70524\ : std_logic;
signal \N__70523\ : std_logic;
signal \N__70522\ : std_logic;
signal \N__70521\ : std_logic;
signal \N__70518\ : std_logic;
signal \N__70515\ : std_logic;
signal \N__70514\ : std_logic;
signal \N__70511\ : std_logic;
signal \N__70500\ : std_logic;
signal \N__70497\ : std_logic;
signal \N__70494\ : std_logic;
signal \N__70491\ : std_logic;
signal \N__70478\ : std_logic;
signal \N__70475\ : std_logic;
signal \N__70472\ : std_logic;
signal \N__70469\ : std_logic;
signal \N__70468\ : std_logic;
signal \N__70467\ : std_logic;
signal \N__70466\ : std_logic;
signal \N__70463\ : std_logic;
signal \N__70462\ : std_logic;
signal \N__70461\ : std_logic;
signal \N__70460\ : std_logic;
signal \N__70459\ : std_logic;
signal \N__70458\ : std_logic;
signal \N__70457\ : std_logic;
signal \N__70456\ : std_logic;
signal \N__70455\ : std_logic;
signal \N__70452\ : std_logic;
signal \N__70445\ : std_logic;
signal \N__70442\ : std_logic;
signal \N__70437\ : std_logic;
signal \N__70432\ : std_logic;
signal \N__70425\ : std_logic;
signal \N__70422\ : std_logic;
signal \N__70417\ : std_logic;
signal \N__70404\ : std_logic;
signal \N__70401\ : std_logic;
signal \N__70398\ : std_logic;
signal \N__70395\ : std_logic;
signal \N__70390\ : std_logic;
signal \N__70373\ : std_logic;
signal \N__70370\ : std_logic;
signal \N__70369\ : std_logic;
signal \N__70366\ : std_logic;
signal \N__70363\ : std_logic;
signal \N__70360\ : std_logic;
signal \N__70357\ : std_logic;
signal \N__70354\ : std_logic;
signal \N__70351\ : std_logic;
signal \N__70348\ : std_logic;
signal \N__70345\ : std_logic;
signal \N__70340\ : std_logic;
signal \N__70337\ : std_logic;
signal \N__70334\ : std_logic;
signal \N__70331\ : std_logic;
signal \N__70330\ : std_logic;
signal \N__70329\ : std_logic;
signal \N__70328\ : std_logic;
signal \N__70325\ : std_logic;
signal \N__70322\ : std_logic;
signal \N__70319\ : std_logic;
signal \N__70318\ : std_logic;
signal \N__70317\ : std_logic;
signal \N__70314\ : std_logic;
signal \N__70309\ : std_logic;
signal \N__70306\ : std_logic;
signal \N__70303\ : std_logic;
signal \N__70300\ : std_logic;
signal \N__70297\ : std_logic;
signal \N__70292\ : std_logic;
signal \N__70285\ : std_logic;
signal \N__70282\ : std_logic;
signal \N__70279\ : std_logic;
signal \N__70276\ : std_logic;
signal \N__70271\ : std_logic;
signal \N__70268\ : std_logic;
signal \N__70265\ : std_logic;
signal \N__70262\ : std_logic;
signal \N__70259\ : std_logic;
signal \N__70256\ : std_logic;
signal \N__70253\ : std_logic;
signal \N__70250\ : std_logic;
signal \N__70249\ : std_logic;
signal \N__70246\ : std_logic;
signal \N__70243\ : std_logic;
signal \N__70240\ : std_logic;
signal \N__70239\ : std_logic;
signal \N__70236\ : std_logic;
signal \N__70233\ : std_logic;
signal \N__70230\ : std_logic;
signal \N__70227\ : std_logic;
signal \N__70224\ : std_logic;
signal \N__70221\ : std_logic;
signal \N__70218\ : std_logic;
signal \N__70215\ : std_logic;
signal \N__70212\ : std_logic;
signal \N__70209\ : std_logic;
signal \N__70206\ : std_logic;
signal \N__70199\ : std_logic;
signal \N__70198\ : std_logic;
signal \N__70197\ : std_logic;
signal \N__70192\ : std_logic;
signal \N__70191\ : std_logic;
signal \N__70188\ : std_logic;
signal \N__70187\ : std_logic;
signal \N__70186\ : std_logic;
signal \N__70185\ : std_logic;
signal \N__70184\ : std_logic;
signal \N__70181\ : std_logic;
signal \N__70178\ : std_logic;
signal \N__70175\ : std_logic;
signal \N__70172\ : std_logic;
signal \N__70171\ : std_logic;
signal \N__70170\ : std_logic;
signal \N__70169\ : std_logic;
signal \N__70168\ : std_logic;
signal \N__70167\ : std_logic;
signal \N__70160\ : std_logic;
signal \N__70159\ : std_logic;
signal \N__70158\ : std_logic;
signal \N__70157\ : std_logic;
signal \N__70154\ : std_logic;
signal \N__70147\ : std_logic;
signal \N__70140\ : std_logic;
signal \N__70139\ : std_logic;
signal \N__70134\ : std_logic;
signal \N__70131\ : std_logic;
signal \N__70128\ : std_logic;
signal \N__70123\ : std_logic;
signal \N__70118\ : std_logic;
signal \N__70117\ : std_logic;
signal \N__70114\ : std_logic;
signal \N__70111\ : std_logic;
signal \N__70106\ : std_logic;
signal \N__70103\ : std_logic;
signal \N__70100\ : std_logic;
signal \N__70097\ : std_logic;
signal \N__70096\ : std_logic;
signal \N__70095\ : std_logic;
signal \N__70094\ : std_logic;
signal \N__70091\ : std_logic;
signal \N__70090\ : std_logic;
signal \N__70089\ : std_logic;
signal \N__70088\ : std_logic;
signal \N__70085\ : std_logic;
signal \N__70080\ : std_logic;
signal \N__70075\ : std_logic;
signal \N__70072\ : std_logic;
signal \N__70065\ : std_logic;
signal \N__70062\ : std_logic;
signal \N__70055\ : std_logic;
signal \N__70054\ : std_logic;
signal \N__70047\ : std_logic;
signal \N__70042\ : std_logic;
signal \N__70037\ : std_logic;
signal \N__70034\ : std_logic;
signal \N__70031\ : std_logic;
signal \N__70028\ : std_logic;
signal \N__70025\ : std_logic;
signal \N__70016\ : std_logic;
signal \N__70013\ : std_logic;
signal \N__70012\ : std_logic;
signal \N__70011\ : std_logic;
signal \N__70008\ : std_logic;
signal \N__70007\ : std_logic;
signal \N__70004\ : std_logic;
signal \N__70001\ : std_logic;
signal \N__70000\ : std_logic;
signal \N__69999\ : std_logic;
signal \N__69998\ : std_logic;
signal \N__69995\ : std_logic;
signal \N__69992\ : std_logic;
signal \N__69989\ : std_logic;
signal \N__69988\ : std_logic;
signal \N__69983\ : std_logic;
signal \N__69978\ : std_logic;
signal \N__69977\ : std_logic;
signal \N__69974\ : std_logic;
signal \N__69973\ : std_logic;
signal \N__69972\ : std_logic;
signal \N__69969\ : std_logic;
signal \N__69968\ : std_logic;
signal \N__69967\ : std_logic;
signal \N__69966\ : std_logic;
signal \N__69965\ : std_logic;
signal \N__69962\ : std_logic;
signal \N__69959\ : std_logic;
signal \N__69954\ : std_logic;
signal \N__69951\ : std_logic;
signal \N__69948\ : std_logic;
signal \N__69945\ : std_logic;
signal \N__69944\ : std_logic;
signal \N__69943\ : std_logic;
signal \N__69940\ : std_logic;
signal \N__69937\ : std_logic;
signal \N__69932\ : std_logic;
signal \N__69929\ : std_logic;
signal \N__69928\ : std_logic;
signal \N__69925\ : std_logic;
signal \N__69922\ : std_logic;
signal \N__69919\ : std_logic;
signal \N__69914\ : std_logic;
signal \N__69909\ : std_logic;
signal \N__69908\ : std_logic;
signal \N__69907\ : std_logic;
signal \N__69904\ : std_logic;
signal \N__69901\ : std_logic;
signal \N__69898\ : std_logic;
signal \N__69891\ : std_logic;
signal \N__69886\ : std_logic;
signal \N__69885\ : std_logic;
signal \N__69882\ : std_logic;
signal \N__69879\ : std_logic;
signal \N__69876\ : std_logic;
signal \N__69873\ : std_logic;
signal \N__69868\ : std_logic;
signal \N__69863\ : std_logic;
signal \N__69860\ : std_logic;
signal \N__69855\ : std_logic;
signal \N__69852\ : std_logic;
signal \N__69849\ : std_logic;
signal \N__69846\ : std_logic;
signal \N__69839\ : std_logic;
signal \N__69836\ : std_logic;
signal \N__69833\ : std_logic;
signal \N__69830\ : std_logic;
signal \N__69827\ : std_logic;
signal \N__69822\ : std_logic;
signal \N__69819\ : std_logic;
signal \N__69812\ : std_logic;
signal \N__69803\ : std_logic;
signal \N__69800\ : std_logic;
signal \N__69799\ : std_logic;
signal \N__69798\ : std_logic;
signal \N__69791\ : std_logic;
signal \N__69790\ : std_logic;
signal \N__69789\ : std_logic;
signal \N__69786\ : std_logic;
signal \N__69783\ : std_logic;
signal \N__69780\ : std_logic;
signal \N__69773\ : std_logic;
signal \N__69770\ : std_logic;
signal \N__69767\ : std_logic;
signal \N__69766\ : std_logic;
signal \N__69763\ : std_logic;
signal \N__69760\ : std_logic;
signal \N__69757\ : std_logic;
signal \N__69752\ : std_logic;
signal \N__69749\ : std_logic;
signal \N__69748\ : std_logic;
signal \N__69747\ : std_logic;
signal \N__69746\ : std_logic;
signal \N__69745\ : std_logic;
signal \N__69744\ : std_logic;
signal \N__69739\ : std_logic;
signal \N__69736\ : std_logic;
signal \N__69733\ : std_logic;
signal \N__69730\ : std_logic;
signal \N__69729\ : std_logic;
signal \N__69726\ : std_logic;
signal \N__69723\ : std_logic;
signal \N__69720\ : std_logic;
signal \N__69717\ : std_logic;
signal \N__69716\ : std_logic;
signal \N__69715\ : std_logic;
signal \N__69712\ : std_logic;
signal \N__69707\ : std_logic;
signal \N__69700\ : std_logic;
signal \N__69699\ : std_logic;
signal \N__69698\ : std_logic;
signal \N__69697\ : std_logic;
signal \N__69694\ : std_logic;
signal \N__69691\ : std_logic;
signal \N__69690\ : std_logic;
signal \N__69689\ : std_logic;
signal \N__69684\ : std_logic;
signal \N__69681\ : std_logic;
signal \N__69680\ : std_logic;
signal \N__69679\ : std_logic;
signal \N__69678\ : std_logic;
signal \N__69675\ : std_logic;
signal \N__69672\ : std_logic;
signal \N__69667\ : std_logic;
signal \N__69666\ : std_logic;
signal \N__69661\ : std_logic;
signal \N__69658\ : std_logic;
signal \N__69655\ : std_logic;
signal \N__69652\ : std_logic;
signal \N__69651\ : std_logic;
signal \N__69648\ : std_logic;
signal \N__69647\ : std_logic;
signal \N__69646\ : std_logic;
signal \N__69645\ : std_logic;
signal \N__69642\ : std_logic;
signal \N__69641\ : std_logic;
signal \N__69640\ : std_logic;
signal \N__69637\ : std_logic;
signal \N__69634\ : std_logic;
signal \N__69631\ : std_logic;
signal \N__69628\ : std_logic;
signal \N__69627\ : std_logic;
signal \N__69624\ : std_logic;
signal \N__69621\ : std_logic;
signal \N__69618\ : std_logic;
signal \N__69613\ : std_logic;
signal \N__69610\ : std_logic;
signal \N__69603\ : std_logic;
signal \N__69596\ : std_logic;
signal \N__69593\ : std_logic;
signal \N__69590\ : std_logic;
signal \N__69583\ : std_logic;
signal \N__69580\ : std_logic;
signal \N__69577\ : std_logic;
signal \N__69574\ : std_logic;
signal \N__69563\ : std_logic;
signal \N__69560\ : std_logic;
signal \N__69555\ : std_logic;
signal \N__69552\ : std_logic;
signal \N__69547\ : std_logic;
signal \N__69544\ : std_logic;
signal \N__69539\ : std_logic;
signal \N__69530\ : std_logic;
signal \N__69529\ : std_logic;
signal \N__69526\ : std_logic;
signal \N__69523\ : std_logic;
signal \N__69520\ : std_logic;
signal \N__69519\ : std_logic;
signal \N__69514\ : std_logic;
signal \N__69513\ : std_logic;
signal \N__69512\ : std_logic;
signal \N__69509\ : std_logic;
signal \N__69506\ : std_logic;
signal \N__69503\ : std_logic;
signal \N__69500\ : std_logic;
signal \N__69497\ : std_logic;
signal \N__69496\ : std_logic;
signal \N__69493\ : std_logic;
signal \N__69490\ : std_logic;
signal \N__69487\ : std_logic;
signal \N__69484\ : std_logic;
signal \N__69481\ : std_logic;
signal \N__69478\ : std_logic;
signal \N__69473\ : std_logic;
signal \N__69470\ : std_logic;
signal \N__69467\ : std_logic;
signal \N__69458\ : std_logic;
signal \N__69455\ : std_logic;
signal \N__69454\ : std_logic;
signal \N__69453\ : std_logic;
signal \N__69452\ : std_logic;
signal \N__69451\ : std_logic;
signal \N__69450\ : std_logic;
signal \N__69449\ : std_logic;
signal \N__69446\ : std_logic;
signal \N__69443\ : std_logic;
signal \N__69440\ : std_logic;
signal \N__69437\ : std_logic;
signal \N__69434\ : std_logic;
signal \N__69431\ : std_logic;
signal \N__69428\ : std_logic;
signal \N__69425\ : std_logic;
signal \N__69422\ : std_logic;
signal \N__69419\ : std_logic;
signal \N__69416\ : std_logic;
signal \N__69413\ : std_logic;
signal \N__69408\ : std_logic;
signal \N__69405\ : std_logic;
signal \N__69402\ : std_logic;
signal \N__69399\ : std_logic;
signal \N__69396\ : std_logic;
signal \N__69393\ : std_logic;
signal \N__69390\ : std_logic;
signal \N__69387\ : std_logic;
signal \N__69382\ : std_logic;
signal \N__69379\ : std_logic;
signal \N__69376\ : std_logic;
signal \N__69373\ : std_logic;
signal \N__69370\ : std_logic;
signal \N__69359\ : std_logic;
signal \N__69356\ : std_logic;
signal \N__69353\ : std_logic;
signal \N__69350\ : std_logic;
signal \N__69347\ : std_logic;
signal \N__69344\ : std_logic;
signal \N__69341\ : std_logic;
signal \N__69338\ : std_logic;
signal \N__69337\ : std_logic;
signal \N__69334\ : std_logic;
signal \N__69333\ : std_logic;
signal \N__69332\ : std_logic;
signal \N__69331\ : std_logic;
signal \N__69324\ : std_logic;
signal \N__69319\ : std_logic;
signal \N__69318\ : std_logic;
signal \N__69317\ : std_logic;
signal \N__69312\ : std_logic;
signal \N__69309\ : std_logic;
signal \N__69306\ : std_logic;
signal \N__69303\ : std_logic;
signal \N__69298\ : std_logic;
signal \N__69295\ : std_logic;
signal \N__69292\ : std_logic;
signal \N__69289\ : std_logic;
signal \N__69284\ : std_logic;
signal \N__69283\ : std_logic;
signal \N__69282\ : std_logic;
signal \N__69281\ : std_logic;
signal \N__69276\ : std_logic;
signal \N__69271\ : std_logic;
signal \N__69270\ : std_logic;
signal \N__69267\ : std_logic;
signal \N__69264\ : std_logic;
signal \N__69261\ : std_logic;
signal \N__69258\ : std_logic;
signal \N__69255\ : std_logic;
signal \N__69248\ : std_logic;
signal \N__69245\ : std_logic;
signal \N__69244\ : std_logic;
signal \N__69243\ : std_logic;
signal \N__69240\ : std_logic;
signal \N__69237\ : std_logic;
signal \N__69234\ : std_logic;
signal \N__69231\ : std_logic;
signal \N__69228\ : std_logic;
signal \N__69225\ : std_logic;
signal \N__69222\ : std_logic;
signal \N__69219\ : std_logic;
signal \N__69216\ : std_logic;
signal \N__69213\ : std_logic;
signal \N__69210\ : std_logic;
signal \N__69207\ : std_logic;
signal \N__69204\ : std_logic;
signal \N__69201\ : std_logic;
signal \N__69198\ : std_logic;
signal \N__69195\ : std_logic;
signal \N__69188\ : std_logic;
signal \N__69185\ : std_logic;
signal \N__69182\ : std_logic;
signal \N__69179\ : std_logic;
signal \N__69176\ : std_logic;
signal \N__69173\ : std_logic;
signal \N__69170\ : std_logic;
signal \N__69169\ : std_logic;
signal \N__69168\ : std_logic;
signal \N__69165\ : std_logic;
signal \N__69162\ : std_logic;
signal \N__69161\ : std_logic;
signal \N__69160\ : std_logic;
signal \N__69157\ : std_logic;
signal \N__69156\ : std_logic;
signal \N__69151\ : std_logic;
signal \N__69150\ : std_logic;
signal \N__69149\ : std_logic;
signal \N__69146\ : std_logic;
signal \N__69143\ : std_logic;
signal \N__69140\ : std_logic;
signal \N__69137\ : std_logic;
signal \N__69134\ : std_logic;
signal \N__69131\ : std_logic;
signal \N__69128\ : std_logic;
signal \N__69121\ : std_logic;
signal \N__69118\ : std_logic;
signal \N__69117\ : std_logic;
signal \N__69112\ : std_logic;
signal \N__69107\ : std_logic;
signal \N__69106\ : std_logic;
signal \N__69103\ : std_logic;
signal \N__69100\ : std_logic;
signal \N__69095\ : std_logic;
signal \N__69092\ : std_logic;
signal \N__69089\ : std_logic;
signal \N__69084\ : std_logic;
signal \N__69077\ : std_logic;
signal \N__69074\ : std_logic;
signal \N__69071\ : std_logic;
signal \N__69070\ : std_logic;
signal \N__69067\ : std_logic;
signal \N__69064\ : std_logic;
signal \N__69061\ : std_logic;
signal \N__69058\ : std_logic;
signal \N__69057\ : std_logic;
signal \N__69054\ : std_logic;
signal \N__69051\ : std_logic;
signal \N__69048\ : std_logic;
signal \N__69045\ : std_logic;
signal \N__69042\ : std_logic;
signal \N__69039\ : std_logic;
signal \N__69036\ : std_logic;
signal \N__69033\ : std_logic;
signal \N__69030\ : std_logic;
signal \N__69027\ : std_logic;
signal \N__69024\ : std_logic;
signal \N__69021\ : std_logic;
signal \N__69014\ : std_logic;
signal \N__69013\ : std_logic;
signal \N__69012\ : std_logic;
signal \N__69011\ : std_logic;
signal \N__69010\ : std_logic;
signal \N__69009\ : std_logic;
signal \N__69006\ : std_logic;
signal \N__69003\ : std_logic;
signal \N__69002\ : std_logic;
signal \N__68999\ : std_logic;
signal \N__68996\ : std_logic;
signal \N__68993\ : std_logic;
signal \N__68990\ : std_logic;
signal \N__68989\ : std_logic;
signal \N__68986\ : std_logic;
signal \N__68983\ : std_logic;
signal \N__68980\ : std_logic;
signal \N__68977\ : std_logic;
signal \N__68970\ : std_logic;
signal \N__68967\ : std_logic;
signal \N__68962\ : std_logic;
signal \N__68955\ : std_logic;
signal \N__68950\ : std_logic;
signal \N__68945\ : std_logic;
signal \N__68944\ : std_logic;
signal \N__68943\ : std_logic;
signal \N__68942\ : std_logic;
signal \N__68941\ : std_logic;
signal \N__68940\ : std_logic;
signal \N__68939\ : std_logic;
signal \N__68936\ : std_logic;
signal \N__68935\ : std_logic;
signal \N__68934\ : std_logic;
signal \N__68933\ : std_logic;
signal \N__68932\ : std_logic;
signal \N__68931\ : std_logic;
signal \N__68930\ : std_logic;
signal \N__68929\ : std_logic;
signal \N__68928\ : std_logic;
signal \N__68927\ : std_logic;
signal \N__68926\ : std_logic;
signal \N__68925\ : std_logic;
signal \N__68924\ : std_logic;
signal \N__68923\ : std_logic;
signal \N__68922\ : std_logic;
signal \N__68921\ : std_logic;
signal \N__68920\ : std_logic;
signal \N__68919\ : std_logic;
signal \N__68918\ : std_logic;
signal \N__68917\ : std_logic;
signal \N__68914\ : std_logic;
signal \N__68911\ : std_logic;
signal \N__68910\ : std_logic;
signal \N__68909\ : std_logic;
signal \N__68908\ : std_logic;
signal \N__68901\ : std_logic;
signal \N__68898\ : std_logic;
signal \N__68897\ : std_logic;
signal \N__68896\ : std_logic;
signal \N__68895\ : std_logic;
signal \N__68894\ : std_logic;
signal \N__68891\ : std_logic;
signal \N__68886\ : std_logic;
signal \N__68883\ : std_logic;
signal \N__68880\ : std_logic;
signal \N__68875\ : std_logic;
signal \N__68872\ : std_logic;
signal \N__68867\ : std_logic;
signal \N__68860\ : std_logic;
signal \N__68855\ : std_logic;
signal \N__68852\ : std_logic;
signal \N__68847\ : std_logic;
signal \N__68846\ : std_logic;
signal \N__68845\ : std_logic;
signal \N__68844\ : std_logic;
signal \N__68843\ : std_logic;
signal \N__68842\ : std_logic;
signal \N__68841\ : std_logic;
signal \N__68836\ : std_logic;
signal \N__68831\ : std_logic;
signal \N__68826\ : std_logic;
signal \N__68825\ : std_logic;
signal \N__68824\ : std_logic;
signal \N__68823\ : std_logic;
signal \N__68822\ : std_logic;
signal \N__68819\ : std_logic;
signal \N__68816\ : std_logic;
signal \N__68813\ : std_logic;
signal \N__68812\ : std_logic;
signal \N__68811\ : std_logic;
signal \N__68810\ : std_logic;
signal \N__68809\ : std_logic;
signal \N__68804\ : std_logic;
signal \N__68799\ : std_logic;
signal \N__68796\ : std_logic;
signal \N__68791\ : std_logic;
signal \N__68790\ : std_logic;
signal \N__68789\ : std_logic;
signal \N__68786\ : std_logic;
signal \N__68783\ : std_logic;
signal \N__68774\ : std_logic;
signal \N__68769\ : std_logic;
signal \N__68762\ : std_logic;
signal \N__68755\ : std_logic;
signal \N__68752\ : std_logic;
signal \N__68747\ : std_logic;
signal \N__68746\ : std_logic;
signal \N__68745\ : std_logic;
signal \N__68744\ : std_logic;
signal \N__68741\ : std_logic;
signal \N__68734\ : std_logic;
signal \N__68733\ : std_logic;
signal \N__68730\ : std_logic;
signal \N__68729\ : std_logic;
signal \N__68728\ : std_logic;
signal \N__68727\ : std_logic;
signal \N__68722\ : std_logic;
signal \N__68721\ : std_logic;
signal \N__68720\ : std_logic;
signal \N__68719\ : std_logic;
signal \N__68712\ : std_logic;
signal \N__68709\ : std_logic;
signal \N__68706\ : std_logic;
signal \N__68703\ : std_logic;
signal \N__68698\ : std_logic;
signal \N__68693\ : std_logic;
signal \N__68690\ : std_logic;
signal \N__68679\ : std_logic;
signal \N__68674\ : std_logic;
signal \N__68667\ : std_logic;
signal \N__68662\ : std_logic;
signal \N__68661\ : std_logic;
signal \N__68660\ : std_logic;
signal \N__68659\ : std_logic;
signal \N__68658\ : std_logic;
signal \N__68655\ : std_logic;
signal \N__68652\ : std_logic;
signal \N__68649\ : std_logic;
signal \N__68646\ : std_logic;
signal \N__68643\ : std_logic;
signal \N__68640\ : std_logic;
signal \N__68637\ : std_logic;
signal \N__68632\ : std_logic;
signal \N__68619\ : std_logic;
signal \N__68614\ : std_logic;
signal \N__68607\ : std_logic;
signal \N__68600\ : std_logic;
signal \N__68595\ : std_logic;
signal \N__68588\ : std_logic;
signal \N__68567\ : std_logic;
signal \N__68566\ : std_logic;
signal \N__68565\ : std_logic;
signal \N__68560\ : std_logic;
signal \N__68557\ : std_logic;
signal \N__68556\ : std_logic;
signal \N__68553\ : std_logic;
signal \N__68550\ : std_logic;
signal \N__68547\ : std_logic;
signal \N__68544\ : std_logic;
signal \N__68541\ : std_logic;
signal \N__68538\ : std_logic;
signal \N__68531\ : std_logic;
signal \N__68530\ : std_logic;
signal \N__68529\ : std_logic;
signal \N__68528\ : std_logic;
signal \N__68527\ : std_logic;
signal \N__68526\ : std_logic;
signal \N__68525\ : std_logic;
signal \N__68524\ : std_logic;
signal \N__68523\ : std_logic;
signal \N__68522\ : std_logic;
signal \N__68521\ : std_logic;
signal \N__68518\ : std_logic;
signal \N__68517\ : std_logic;
signal \N__68516\ : std_logic;
signal \N__68515\ : std_logic;
signal \N__68512\ : std_logic;
signal \N__68511\ : std_logic;
signal \N__68510\ : std_logic;
signal \N__68509\ : std_logic;
signal \N__68508\ : std_logic;
signal \N__68507\ : std_logic;
signal \N__68506\ : std_logic;
signal \N__68505\ : std_logic;
signal \N__68502\ : std_logic;
signal \N__68499\ : std_logic;
signal \N__68494\ : std_logic;
signal \N__68491\ : std_logic;
signal \N__68490\ : std_logic;
signal \N__68485\ : std_logic;
signal \N__68484\ : std_logic;
signal \N__68483\ : std_logic;
signal \N__68482\ : std_logic;
signal \N__68481\ : std_logic;
signal \N__68480\ : std_logic;
signal \N__68479\ : std_logic;
signal \N__68472\ : std_logic;
signal \N__68469\ : std_logic;
signal \N__68468\ : std_logic;
signal \N__68465\ : std_logic;
signal \N__68464\ : std_logic;
signal \N__68461\ : std_logic;
signal \N__68460\ : std_logic;
signal \N__68459\ : std_logic;
signal \N__68458\ : std_logic;
signal \N__68455\ : std_logic;
signal \N__68452\ : std_logic;
signal \N__68445\ : std_logic;
signal \N__68442\ : std_logic;
signal \N__68441\ : std_logic;
signal \N__68440\ : std_logic;
signal \N__68439\ : std_logic;
signal \N__68438\ : std_logic;
signal \N__68435\ : std_logic;
signal \N__68432\ : std_logic;
signal \N__68431\ : std_logic;
signal \N__68426\ : std_logic;
signal \N__68423\ : std_logic;
signal \N__68420\ : std_logic;
signal \N__68417\ : std_logic;
signal \N__68414\ : std_logic;
signal \N__68411\ : std_logic;
signal \N__68404\ : std_logic;
signal \N__68399\ : std_logic;
signal \N__68396\ : std_logic;
signal \N__68395\ : std_logic;
signal \N__68394\ : std_logic;
signal \N__68391\ : std_logic;
signal \N__68388\ : std_logic;
signal \N__68385\ : std_logic;
signal \N__68382\ : std_logic;
signal \N__68379\ : std_logic;
signal \N__68378\ : std_logic;
signal \N__68375\ : std_logic;
signal \N__68374\ : std_logic;
signal \N__68371\ : std_logic;
signal \N__68368\ : std_logic;
signal \N__68359\ : std_logic;
signal \N__68352\ : std_logic;
signal \N__68349\ : std_logic;
signal \N__68346\ : std_logic;
signal \N__68343\ : std_logic;
signal \N__68340\ : std_logic;
signal \N__68329\ : std_logic;
signal \N__68322\ : std_logic;
signal \N__68319\ : std_logic;
signal \N__68316\ : std_logic;
signal \N__68315\ : std_logic;
signal \N__68312\ : std_logic;
signal \N__68309\ : std_logic;
signal \N__68306\ : std_logic;
signal \N__68299\ : std_logic;
signal \N__68292\ : std_logic;
signal \N__68285\ : std_logic;
signal \N__68282\ : std_logic;
signal \N__68281\ : std_logic;
signal \N__68280\ : std_logic;
signal \N__68271\ : std_logic;
signal \N__68270\ : std_logic;
signal \N__68267\ : std_logic;
signal \N__68260\ : std_logic;
signal \N__68257\ : std_logic;
signal \N__68256\ : std_logic;
signal \N__68253\ : std_logic;
signal \N__68240\ : std_logic;
signal \N__68237\ : std_logic;
signal \N__68234\ : std_logic;
signal \N__68233\ : std_logic;
signal \N__68232\ : std_logic;
signal \N__68231\ : std_logic;
signal \N__68230\ : std_logic;
signal \N__68229\ : std_logic;
signal \N__68228\ : std_logic;
signal \N__68225\ : std_logic;
signal \N__68222\ : std_logic;
signal \N__68215\ : std_logic;
signal \N__68212\ : std_logic;
signal \N__68205\ : std_logic;
signal \N__68196\ : std_logic;
signal \N__68189\ : std_logic;
signal \N__68174\ : std_logic;
signal \N__68171\ : std_logic;
signal \N__68168\ : std_logic;
signal \N__68167\ : std_logic;
signal \N__68166\ : std_logic;
signal \N__68163\ : std_logic;
signal \N__68158\ : std_logic;
signal \N__68153\ : std_logic;
signal \N__68150\ : std_logic;
signal \N__68147\ : std_logic;
signal \N__68144\ : std_logic;
signal \N__68141\ : std_logic;
signal \N__68140\ : std_logic;
signal \N__68139\ : std_logic;
signal \N__68138\ : std_logic;
signal \N__68137\ : std_logic;
signal \N__68136\ : std_logic;
signal \N__68133\ : std_logic;
signal \N__68130\ : std_logic;
signal \N__68127\ : std_logic;
signal \N__68124\ : std_logic;
signal \N__68123\ : std_logic;
signal \N__68122\ : std_logic;
signal \N__68119\ : std_logic;
signal \N__68116\ : std_logic;
signal \N__68109\ : std_logic;
signal \N__68106\ : std_logic;
signal \N__68103\ : std_logic;
signal \N__68100\ : std_logic;
signal \N__68087\ : std_logic;
signal \N__68086\ : std_logic;
signal \N__68083\ : std_logic;
signal \N__68080\ : std_logic;
signal \N__68079\ : std_logic;
signal \N__68078\ : std_logic;
signal \N__68077\ : std_logic;
signal \N__68076\ : std_logic;
signal \N__68071\ : std_logic;
signal \N__68068\ : std_logic;
signal \N__68065\ : std_logic;
signal \N__68062\ : std_logic;
signal \N__68059\ : std_logic;
signal \N__68058\ : std_logic;
signal \N__68057\ : std_logic;
signal \N__68054\ : std_logic;
signal \N__68049\ : std_logic;
signal \N__68046\ : std_logic;
signal \N__68043\ : std_logic;
signal \N__68040\ : std_logic;
signal \N__68037\ : std_logic;
signal \N__68034\ : std_logic;
signal \N__68023\ : std_logic;
signal \N__68020\ : std_logic;
signal \N__68017\ : std_logic;
signal \N__68012\ : std_logic;
signal \N__68011\ : std_logic;
signal \N__68008\ : std_logic;
signal \N__68005\ : std_logic;
signal \N__68004\ : std_logic;
signal \N__68003\ : std_logic;
signal \N__68002\ : std_logic;
signal \N__68001\ : std_logic;
signal \N__68000\ : std_logic;
signal \N__67997\ : std_logic;
signal \N__67994\ : std_logic;
signal \N__67991\ : std_logic;
signal \N__67988\ : std_logic;
signal \N__67985\ : std_logic;
signal \N__67982\ : std_logic;
signal \N__67979\ : std_logic;
signal \N__67964\ : std_logic;
signal \N__67963\ : std_logic;
signal \N__67960\ : std_logic;
signal \N__67957\ : std_logic;
signal \N__67952\ : std_logic;
signal \N__67949\ : std_logic;
signal \N__67946\ : std_logic;
signal \N__67943\ : std_logic;
signal \N__67942\ : std_logic;
signal \N__67939\ : std_logic;
signal \N__67938\ : std_logic;
signal \N__67935\ : std_logic;
signal \N__67932\ : std_logic;
signal \N__67931\ : std_logic;
signal \N__67928\ : std_logic;
signal \N__67925\ : std_logic;
signal \N__67922\ : std_logic;
signal \N__67921\ : std_logic;
signal \N__67918\ : std_logic;
signal \N__67915\ : std_logic;
signal \N__67912\ : std_logic;
signal \N__67909\ : std_logic;
signal \N__67906\ : std_logic;
signal \N__67903\ : std_logic;
signal \N__67900\ : std_logic;
signal \N__67897\ : std_logic;
signal \N__67894\ : std_logic;
signal \N__67891\ : std_logic;
signal \N__67888\ : std_logic;
signal \N__67885\ : std_logic;
signal \N__67880\ : std_logic;
signal \N__67871\ : std_logic;
signal \N__67868\ : std_logic;
signal \N__67865\ : std_logic;
signal \N__67864\ : std_logic;
signal \N__67861\ : std_logic;
signal \N__67860\ : std_logic;
signal \N__67857\ : std_logic;
signal \N__67854\ : std_logic;
signal \N__67851\ : std_logic;
signal \N__67848\ : std_logic;
signal \N__67845\ : std_logic;
signal \N__67842\ : std_logic;
signal \N__67839\ : std_logic;
signal \N__67836\ : std_logic;
signal \N__67833\ : std_logic;
signal \N__67830\ : std_logic;
signal \N__67827\ : std_logic;
signal \N__67820\ : std_logic;
signal \N__67817\ : std_logic;
signal \N__67814\ : std_logic;
signal \N__67811\ : std_logic;
signal \N__67808\ : std_logic;
signal \N__67805\ : std_logic;
signal \N__67802\ : std_logic;
signal \N__67799\ : std_logic;
signal \N__67796\ : std_logic;
signal \N__67793\ : std_logic;
signal \N__67790\ : std_logic;
signal \N__67787\ : std_logic;
signal \N__67784\ : std_logic;
signal \N__67783\ : std_logic;
signal \N__67780\ : std_logic;
signal \N__67777\ : std_logic;
signal \N__67774\ : std_logic;
signal \N__67771\ : std_logic;
signal \N__67766\ : std_logic;
signal \N__67763\ : std_logic;
signal \N__67760\ : std_logic;
signal \N__67757\ : std_logic;
signal \N__67756\ : std_logic;
signal \N__67755\ : std_logic;
signal \N__67754\ : std_logic;
signal \N__67753\ : std_logic;
signal \N__67750\ : std_logic;
signal \N__67747\ : std_logic;
signal \N__67744\ : std_logic;
signal \N__67743\ : std_logic;
signal \N__67742\ : std_logic;
signal \N__67741\ : std_logic;
signal \N__67738\ : std_logic;
signal \N__67735\ : std_logic;
signal \N__67732\ : std_logic;
signal \N__67729\ : std_logic;
signal \N__67726\ : std_logic;
signal \N__67723\ : std_logic;
signal \N__67720\ : std_logic;
signal \N__67717\ : std_logic;
signal \N__67712\ : std_logic;
signal \N__67707\ : std_logic;
signal \N__67704\ : std_logic;
signal \N__67691\ : std_logic;
signal \N__67688\ : std_logic;
signal \N__67687\ : std_logic;
signal \N__67686\ : std_logic;
signal \N__67685\ : std_logic;
signal \N__67682\ : std_logic;
signal \N__67679\ : std_logic;
signal \N__67676\ : std_logic;
signal \N__67673\ : std_logic;
signal \N__67672\ : std_logic;
signal \N__67669\ : std_logic;
signal \N__67668\ : std_logic;
signal \N__67665\ : std_logic;
signal \N__67662\ : std_logic;
signal \N__67659\ : std_logic;
signal \N__67656\ : std_logic;
signal \N__67655\ : std_logic;
signal \N__67654\ : std_logic;
signal \N__67651\ : std_logic;
signal \N__67648\ : std_logic;
signal \N__67639\ : std_logic;
signal \N__67636\ : std_logic;
signal \N__67633\ : std_logic;
signal \N__67622\ : std_logic;
signal \N__67621\ : std_logic;
signal \N__67618\ : std_logic;
signal \N__67617\ : std_logic;
signal \N__67614\ : std_logic;
signal \N__67611\ : std_logic;
signal \N__67610\ : std_logic;
signal \N__67607\ : std_logic;
signal \N__67604\ : std_logic;
signal \N__67603\ : std_logic;
signal \N__67602\ : std_logic;
signal \N__67599\ : std_logic;
signal \N__67596\ : std_logic;
signal \N__67595\ : std_logic;
signal \N__67590\ : std_logic;
signal \N__67587\ : std_logic;
signal \N__67584\ : std_logic;
signal \N__67581\ : std_logic;
signal \N__67578\ : std_logic;
signal \N__67575\ : std_logic;
signal \N__67570\ : std_logic;
signal \N__67567\ : std_logic;
signal \N__67556\ : std_logic;
signal \N__67553\ : std_logic;
signal \N__67550\ : std_logic;
signal \N__67549\ : std_logic;
signal \N__67546\ : std_logic;
signal \N__67543\ : std_logic;
signal \N__67538\ : std_logic;
signal \N__67535\ : std_logic;
signal \N__67532\ : std_logic;
signal \N__67529\ : std_logic;
signal \N__67526\ : std_logic;
signal \N__67523\ : std_logic;
signal \N__67520\ : std_logic;
signal \N__67517\ : std_logic;
signal \N__67516\ : std_logic;
signal \N__67513\ : std_logic;
signal \N__67512\ : std_logic;
signal \N__67509\ : std_logic;
signal \N__67508\ : std_logic;
signal \N__67505\ : std_logic;
signal \N__67504\ : std_logic;
signal \N__67501\ : std_logic;
signal \N__67498\ : std_logic;
signal \N__67495\ : std_logic;
signal \N__67494\ : std_logic;
signal \N__67493\ : std_logic;
signal \N__67490\ : std_logic;
signal \N__67487\ : std_logic;
signal \N__67484\ : std_logic;
signal \N__67479\ : std_logic;
signal \N__67476\ : std_logic;
signal \N__67473\ : std_logic;
signal \N__67460\ : std_logic;
signal \N__67459\ : std_logic;
signal \N__67456\ : std_logic;
signal \N__67455\ : std_logic;
signal \N__67452\ : std_logic;
signal \N__67451\ : std_logic;
signal \N__67450\ : std_logic;
signal \N__67449\ : std_logic;
signal \N__67446\ : std_logic;
signal \N__67443\ : std_logic;
signal \N__67442\ : std_logic;
signal \N__67439\ : std_logic;
signal \N__67436\ : std_logic;
signal \N__67433\ : std_logic;
signal \N__67432\ : std_logic;
signal \N__67429\ : std_logic;
signal \N__67424\ : std_logic;
signal \N__67421\ : std_logic;
signal \N__67414\ : std_logic;
signal \N__67411\ : std_logic;
signal \N__67400\ : std_logic;
signal \N__67399\ : std_logic;
signal \N__67396\ : std_logic;
signal \N__67393\ : std_logic;
signal \N__67392\ : std_logic;
signal \N__67391\ : std_logic;
signal \N__67390\ : std_logic;
signal \N__67389\ : std_logic;
signal \N__67388\ : std_logic;
signal \N__67385\ : std_logic;
signal \N__67382\ : std_logic;
signal \N__67379\ : std_logic;
signal \N__67376\ : std_logic;
signal \N__67373\ : std_logic;
signal \N__67370\ : std_logic;
signal \N__67367\ : std_logic;
signal \N__67352\ : std_logic;
signal \N__67349\ : std_logic;
signal \N__67348\ : std_logic;
signal \N__67345\ : std_logic;
signal \N__67342\ : std_logic;
signal \N__67339\ : std_logic;
signal \N__67336\ : std_logic;
signal \N__67333\ : std_logic;
signal \N__67330\ : std_logic;
signal \N__67327\ : std_logic;
signal \N__67324\ : std_logic;
signal \N__67321\ : std_logic;
signal \N__67316\ : std_logic;
signal \N__67313\ : std_logic;
signal \N__67312\ : std_logic;
signal \N__67309\ : std_logic;
signal \N__67306\ : std_logic;
signal \N__67303\ : std_logic;
signal \N__67300\ : std_logic;
signal \N__67297\ : std_logic;
signal \N__67294\ : std_logic;
signal \N__67289\ : std_logic;
signal \N__67286\ : std_logic;
signal \N__67283\ : std_logic;
signal \N__67282\ : std_logic;
signal \N__67277\ : std_logic;
signal \N__67274\ : std_logic;
signal \N__67273\ : std_logic;
signal \N__67272\ : std_logic;
signal \N__67271\ : std_logic;
signal \N__67270\ : std_logic;
signal \N__67269\ : std_logic;
signal \N__67268\ : std_logic;
signal \N__67267\ : std_logic;
signal \N__67266\ : std_logic;
signal \N__67263\ : std_logic;
signal \N__67256\ : std_logic;
signal \N__67255\ : std_logic;
signal \N__67254\ : std_logic;
signal \N__67253\ : std_logic;
signal \N__67252\ : std_logic;
signal \N__67251\ : std_logic;
signal \N__67250\ : std_logic;
signal \N__67249\ : std_logic;
signal \N__67248\ : std_logic;
signal \N__67245\ : std_logic;
signal \N__67244\ : std_logic;
signal \N__67243\ : std_logic;
signal \N__67242\ : std_logic;
signal \N__67239\ : std_logic;
signal \N__67236\ : std_logic;
signal \N__67233\ : std_logic;
signal \N__67232\ : std_logic;
signal \N__67231\ : std_logic;
signal \N__67230\ : std_logic;
signal \N__67227\ : std_logic;
signal \N__67226\ : std_logic;
signal \N__67225\ : std_logic;
signal \N__67220\ : std_logic;
signal \N__67219\ : std_logic;
signal \N__67218\ : std_logic;
signal \N__67217\ : std_logic;
signal \N__67216\ : std_logic;
signal \N__67215\ : std_logic;
signal \N__67214\ : std_logic;
signal \N__67213\ : std_logic;
signal \N__67212\ : std_logic;
signal \N__67209\ : std_logic;
signal \N__67208\ : std_logic;
signal \N__67207\ : std_logic;
signal \N__67206\ : std_logic;
signal \N__67205\ : std_logic;
signal \N__67204\ : std_logic;
signal \N__67197\ : std_logic;
signal \N__67184\ : std_logic;
signal \N__67183\ : std_logic;
signal \N__67180\ : std_logic;
signal \N__67179\ : std_logic;
signal \N__67176\ : std_logic;
signal \N__67173\ : std_logic;
signal \N__67170\ : std_logic;
signal \N__67165\ : std_logic;
signal \N__67164\ : std_logic;
signal \N__67161\ : std_logic;
signal \N__67158\ : std_logic;
signal \N__67151\ : std_logic;
signal \N__67148\ : std_logic;
signal \N__67145\ : std_logic;
signal \N__67138\ : std_logic;
signal \N__67135\ : std_logic;
signal \N__67130\ : std_logic;
signal \N__67123\ : std_logic;
signal \N__67116\ : std_logic;
signal \N__67115\ : std_logic;
signal \N__67112\ : std_logic;
signal \N__67107\ : std_logic;
signal \N__67100\ : std_logic;
signal \N__67097\ : std_logic;
signal \N__67090\ : std_logic;
signal \N__67087\ : std_logic;
signal \N__67066\ : std_logic;
signal \N__67065\ : std_logic;
signal \N__67064\ : std_logic;
signal \N__67061\ : std_logic;
signal \N__67060\ : std_logic;
signal \N__67057\ : std_logic;
signal \N__67054\ : std_logic;
signal \N__67053\ : std_logic;
signal \N__67052\ : std_logic;
signal \N__67051\ : std_logic;
signal \N__67048\ : std_logic;
signal \N__67047\ : std_logic;
signal \N__67046\ : std_logic;
signal \N__67045\ : std_logic;
signal \N__67044\ : std_logic;
signal \N__67043\ : std_logic;
signal \N__67042\ : std_logic;
signal \N__67039\ : std_logic;
signal \N__67036\ : std_logic;
signal \N__67033\ : std_logic;
signal \N__67030\ : std_logic;
signal \N__67027\ : std_logic;
signal \N__67020\ : std_logic;
signal \N__67017\ : std_logic;
signal \N__67014\ : std_logic;
signal \N__67007\ : std_logic;
signal \N__67004\ : std_logic;
signal \N__66997\ : std_logic;
signal \N__66994\ : std_logic;
signal \N__66991\ : std_logic;
signal \N__66988\ : std_logic;
signal \N__66985\ : std_logic;
signal \N__66982\ : std_logic;
signal \N__66977\ : std_logic;
signal \N__66976\ : std_logic;
signal \N__66973\ : std_logic;
signal \N__66970\ : std_logic;
signal \N__66963\ : std_logic;
signal \N__66958\ : std_logic;
signal \N__66951\ : std_logic;
signal \N__66948\ : std_logic;
signal \N__66945\ : std_logic;
signal \N__66942\ : std_logic;
signal \N__66939\ : std_logic;
signal \N__66930\ : std_logic;
signal \N__66927\ : std_logic;
signal \N__66920\ : std_logic;
signal \N__66915\ : std_logic;
signal \N__66910\ : std_logic;
signal \N__66907\ : std_logic;
signal \N__66902\ : std_logic;
signal \N__66901\ : std_logic;
signal \N__66898\ : std_logic;
signal \N__66897\ : std_logic;
signal \N__66896\ : std_logic;
signal \N__66891\ : std_logic;
signal \N__66888\ : std_logic;
signal \N__66885\ : std_logic;
signal \N__66882\ : std_logic;
signal \N__66879\ : std_logic;
signal \N__66876\ : std_logic;
signal \N__66873\ : std_logic;
signal \N__66870\ : std_logic;
signal \N__66865\ : std_logic;
signal \N__66860\ : std_logic;
signal \N__66857\ : std_logic;
signal \N__66856\ : std_logic;
signal \N__66853\ : std_logic;
signal \N__66850\ : std_logic;
signal \N__66845\ : std_logic;
signal \N__66844\ : std_logic;
signal \N__66843\ : std_logic;
signal \N__66840\ : std_logic;
signal \N__66837\ : std_logic;
signal \N__66834\ : std_logic;
signal \N__66833\ : std_logic;
signal \N__66832\ : std_logic;
signal \N__66831\ : std_logic;
signal \N__66828\ : std_logic;
signal \N__66827\ : std_logic;
signal \N__66822\ : std_logic;
signal \N__66819\ : std_logic;
signal \N__66816\ : std_logic;
signal \N__66813\ : std_logic;
signal \N__66810\ : std_logic;
signal \N__66807\ : std_logic;
signal \N__66806\ : std_logic;
signal \N__66801\ : std_logic;
signal \N__66796\ : std_logic;
signal \N__66791\ : std_logic;
signal \N__66788\ : std_logic;
signal \N__66785\ : std_logic;
signal \N__66778\ : std_logic;
signal \N__66773\ : std_logic;
signal \N__66772\ : std_logic;
signal \N__66769\ : std_logic;
signal \N__66768\ : std_logic;
signal \N__66767\ : std_logic;
signal \N__66766\ : std_logic;
signal \N__66765\ : std_logic;
signal \N__66764\ : std_logic;
signal \N__66763\ : std_logic;
signal \N__66762\ : std_logic;
signal \N__66761\ : std_logic;
signal \N__66758\ : std_logic;
signal \N__66757\ : std_logic;
signal \N__66756\ : std_logic;
signal \N__66755\ : std_logic;
signal \N__66754\ : std_logic;
signal \N__66753\ : std_logic;
signal \N__66750\ : std_logic;
signal \N__66747\ : std_logic;
signal \N__66746\ : std_logic;
signal \N__66743\ : std_logic;
signal \N__66742\ : std_logic;
signal \N__66737\ : std_logic;
signal \N__66736\ : std_logic;
signal \N__66735\ : std_logic;
signal \N__66734\ : std_logic;
signal \N__66733\ : std_logic;
signal \N__66730\ : std_logic;
signal \N__66727\ : std_logic;
signal \N__66722\ : std_logic;
signal \N__66721\ : std_logic;
signal \N__66720\ : std_logic;
signal \N__66719\ : std_logic;
signal \N__66718\ : std_logic;
signal \N__66717\ : std_logic;
signal \N__66716\ : std_logic;
signal \N__66715\ : std_logic;
signal \N__66714\ : std_logic;
signal \N__66713\ : std_logic;
signal \N__66710\ : std_logic;
signal \N__66705\ : std_logic;
signal \N__66704\ : std_logic;
signal \N__66703\ : std_logic;
signal \N__66702\ : std_logic;
signal \N__66701\ : std_logic;
signal \N__66700\ : std_logic;
signal \N__66699\ : std_logic;
signal \N__66698\ : std_logic;
signal \N__66697\ : std_logic;
signal \N__66696\ : std_logic;
signal \N__66693\ : std_logic;
signal \N__66690\ : std_logic;
signal \N__66687\ : std_logic;
signal \N__66686\ : std_logic;
signal \N__66685\ : std_logic;
signal \N__66684\ : std_logic;
signal \N__66683\ : std_logic;
signal \N__66682\ : std_logic;
signal \N__66677\ : std_logic;
signal \N__66672\ : std_logic;
signal \N__66669\ : std_logic;
signal \N__66666\ : std_logic;
signal \N__66663\ : std_logic;
signal \N__66662\ : std_logic;
signal \N__66659\ : std_logic;
signal \N__66654\ : std_logic;
signal \N__66653\ : std_logic;
signal \N__66652\ : std_logic;
signal \N__66647\ : std_logic;
signal \N__66644\ : std_logic;
signal \N__66641\ : std_logic;
signal \N__66634\ : std_logic;
signal \N__66631\ : std_logic;
signal \N__66630\ : std_logic;
signal \N__66629\ : std_logic;
signal \N__66626\ : std_logic;
signal \N__66623\ : std_logic;
signal \N__66618\ : std_logic;
signal \N__66615\ : std_logic;
signal \N__66612\ : std_logic;
signal \N__66609\ : std_logic;
signal \N__66604\ : std_logic;
signal \N__66603\ : std_logic;
signal \N__66602\ : std_logic;
signal \N__66601\ : std_logic;
signal \N__66600\ : std_logic;
signal \N__66599\ : std_logic;
signal \N__66598\ : std_logic;
signal \N__66597\ : std_logic;
signal \N__66596\ : std_logic;
signal \N__66591\ : std_logic;
signal \N__66586\ : std_logic;
signal \N__66583\ : std_logic;
signal \N__66582\ : std_logic;
signal \N__66581\ : std_logic;
signal \N__66580\ : std_logic;
signal \N__66579\ : std_logic;
signal \N__66578\ : std_logic;
signal \N__66577\ : std_logic;
signal \N__66574\ : std_logic;
signal \N__66571\ : std_logic;
signal \N__66570\ : std_logic;
signal \N__66569\ : std_logic;
signal \N__66564\ : std_logic;
signal \N__66559\ : std_logic;
signal \N__66552\ : std_logic;
signal \N__66547\ : std_logic;
signal \N__66540\ : std_logic;
signal \N__66537\ : std_logic;
signal \N__66532\ : std_logic;
signal \N__66529\ : std_logic;
signal \N__66526\ : std_logic;
signal \N__66523\ : std_logic;
signal \N__66516\ : std_logic;
signal \N__66513\ : std_logic;
signal \N__66508\ : std_logic;
signal \N__66501\ : std_logic;
signal \N__66492\ : std_logic;
signal \N__66487\ : std_logic;
signal \N__66482\ : std_logic;
signal \N__66473\ : std_logic;
signal \N__66468\ : std_logic;
signal \N__66465\ : std_logic;
signal \N__66462\ : std_logic;
signal \N__66451\ : std_logic;
signal \N__66448\ : std_logic;
signal \N__66445\ : std_logic;
signal \N__66442\ : std_logic;
signal \N__66441\ : std_logic;
signal \N__66438\ : std_logic;
signal \N__66435\ : std_logic;
signal \N__66426\ : std_logic;
signal \N__66421\ : std_logic;
signal \N__66418\ : std_logic;
signal \N__66415\ : std_logic;
signal \N__66410\ : std_logic;
signal \N__66401\ : std_logic;
signal \N__66394\ : std_logic;
signal \N__66385\ : std_logic;
signal \N__66378\ : std_logic;
signal \N__66377\ : std_logic;
signal \N__66376\ : std_logic;
signal \N__66375\ : std_logic;
signal \N__66372\ : std_logic;
signal \N__66369\ : std_logic;
signal \N__66362\ : std_logic;
signal \N__66355\ : std_logic;
signal \N__66350\ : std_logic;
signal \N__66345\ : std_logic;
signal \N__66340\ : std_logic;
signal \N__66337\ : std_logic;
signal \N__66320\ : std_logic;
signal \N__66317\ : std_logic;
signal \N__66316\ : std_logic;
signal \N__66315\ : std_logic;
signal \N__66314\ : std_logic;
signal \N__66313\ : std_logic;
signal \N__66312\ : std_logic;
signal \N__66309\ : std_logic;
signal \N__66304\ : std_logic;
signal \N__66303\ : std_logic;
signal \N__66300\ : std_logic;
signal \N__66299\ : std_logic;
signal \N__66298\ : std_logic;
signal \N__66297\ : std_logic;
signal \N__66296\ : std_logic;
signal \N__66293\ : std_logic;
signal \N__66292\ : std_logic;
signal \N__66289\ : std_logic;
signal \N__66288\ : std_logic;
signal \N__66287\ : std_logic;
signal \N__66284\ : std_logic;
signal \N__66281\ : std_logic;
signal \N__66278\ : std_logic;
signal \N__66275\ : std_logic;
signal \N__66272\ : std_logic;
signal \N__66271\ : std_logic;
signal \N__66270\ : std_logic;
signal \N__66269\ : std_logic;
signal \N__66266\ : std_logic;
signal \N__66263\ : std_logic;
signal \N__66260\ : std_logic;
signal \N__66257\ : std_logic;
signal \N__66254\ : std_logic;
signal \N__66253\ : std_logic;
signal \N__66252\ : std_logic;
signal \N__66251\ : std_logic;
signal \N__66250\ : std_logic;
signal \N__66249\ : std_logic;
signal \N__66248\ : std_logic;
signal \N__66245\ : std_logic;
signal \N__66242\ : std_logic;
signal \N__66241\ : std_logic;
signal \N__66240\ : std_logic;
signal \N__66237\ : std_logic;
signal \N__66230\ : std_logic;
signal \N__66229\ : std_logic;
signal \N__66228\ : std_logic;
signal \N__66225\ : std_logic;
signal \N__66222\ : std_logic;
signal \N__66215\ : std_logic;
signal \N__66208\ : std_logic;
signal \N__66203\ : std_logic;
signal \N__66198\ : std_logic;
signal \N__66195\ : std_logic;
signal \N__66188\ : std_logic;
signal \N__66183\ : std_logic;
signal \N__66180\ : std_logic;
signal \N__66177\ : std_logic;
signal \N__66176\ : std_logic;
signal \N__66175\ : std_logic;
signal \N__66174\ : std_logic;
signal \N__66169\ : std_logic;
signal \N__66164\ : std_logic;
signal \N__66161\ : std_logic;
signal \N__66154\ : std_logic;
signal \N__66151\ : std_logic;
signal \N__66140\ : std_logic;
signal \N__66137\ : std_logic;
signal \N__66134\ : std_logic;
signal \N__66131\ : std_logic;
signal \N__66128\ : std_logic;
signal \N__66127\ : std_logic;
signal \N__66124\ : std_logic;
signal \N__66117\ : std_logic;
signal \N__66112\ : std_logic;
signal \N__66103\ : std_logic;
signal \N__66100\ : std_logic;
signal \N__66089\ : std_logic;
signal \N__66086\ : std_logic;
signal \N__66085\ : std_logic;
signal \N__66084\ : std_logic;
signal \N__66083\ : std_logic;
signal \N__66082\ : std_logic;
signal \N__66081\ : std_logic;
signal \N__66080\ : std_logic;
signal \N__66079\ : std_logic;
signal \N__66078\ : std_logic;
signal \N__66077\ : std_logic;
signal \N__66076\ : std_logic;
signal \N__66075\ : std_logic;
signal \N__66074\ : std_logic;
signal \N__66073\ : std_logic;
signal \N__66068\ : std_logic;
signal \N__66067\ : std_logic;
signal \N__66066\ : std_logic;
signal \N__66065\ : std_logic;
signal \N__66064\ : std_logic;
signal \N__66063\ : std_logic;
signal \N__66062\ : std_logic;
signal \N__66061\ : std_logic;
signal \N__66060\ : std_logic;
signal \N__66059\ : std_logic;
signal \N__66058\ : std_logic;
signal \N__66055\ : std_logic;
signal \N__66052\ : std_logic;
signal \N__66051\ : std_logic;
signal \N__66050\ : std_logic;
signal \N__66049\ : std_logic;
signal \N__66048\ : std_logic;
signal \N__66047\ : std_logic;
signal \N__66046\ : std_logic;
signal \N__66045\ : std_logic;
signal \N__66040\ : std_logic;
signal \N__66037\ : std_logic;
signal \N__66030\ : std_logic;
signal \N__66029\ : std_logic;
signal \N__66028\ : std_logic;
signal \N__66027\ : std_logic;
signal \N__66026\ : std_logic;
signal \N__66023\ : std_logic;
signal \N__66020\ : std_logic;
signal \N__66015\ : std_logic;
signal \N__66014\ : std_logic;
signal \N__66013\ : std_logic;
signal \N__66012\ : std_logic;
signal \N__66011\ : std_logic;
signal \N__66010\ : std_logic;
signal \N__66007\ : std_logic;
signal \N__66000\ : std_logic;
signal \N__65991\ : std_logic;
signal \N__65990\ : std_logic;
signal \N__65989\ : std_logic;
signal \N__65986\ : std_logic;
signal \N__65981\ : std_logic;
signal \N__65978\ : std_logic;
signal \N__65969\ : std_logic;
signal \N__65968\ : std_logic;
signal \N__65967\ : std_logic;
signal \N__65966\ : std_logic;
signal \N__65965\ : std_logic;
signal \N__65964\ : std_logic;
signal \N__65963\ : std_logic;
signal \N__65962\ : std_logic;
signal \N__65959\ : std_logic;
signal \N__65958\ : std_logic;
signal \N__65957\ : std_logic;
signal \N__65956\ : std_logic;
signal \N__65955\ : std_logic;
signal \N__65954\ : std_logic;
signal \N__65953\ : std_logic;
signal \N__65952\ : std_logic;
signal \N__65951\ : std_logic;
signal \N__65944\ : std_logic;
signal \N__65937\ : std_logic;
signal \N__65936\ : std_logic;
signal \N__65935\ : std_logic;
signal \N__65932\ : std_logic;
signal \N__65931\ : std_logic;
signal \N__65930\ : std_logic;
signal \N__65929\ : std_logic;
signal \N__65928\ : std_logic;
signal \N__65927\ : std_logic;
signal \N__65926\ : std_logic;
signal \N__65921\ : std_logic;
signal \N__65918\ : std_logic;
signal \N__65911\ : std_logic;
signal \N__65906\ : std_logic;
signal \N__65905\ : std_logic;
signal \N__65904\ : std_logic;
signal \N__65903\ : std_logic;
signal \N__65902\ : std_logic;
signal \N__65899\ : std_logic;
signal \N__65896\ : std_logic;
signal \N__65893\ : std_logic;
signal \N__65890\ : std_logic;
signal \N__65887\ : std_logic;
signal \N__65884\ : std_logic;
signal \N__65881\ : std_logic;
signal \N__65878\ : std_logic;
signal \N__65873\ : std_logic;
signal \N__65868\ : std_logic;
signal \N__65861\ : std_logic;
signal \N__65852\ : std_logic;
signal \N__65849\ : std_logic;
signal \N__65840\ : std_logic;
signal \N__65837\ : std_logic;
signal \N__65834\ : std_logic;
signal \N__65829\ : std_logic;
signal \N__65828\ : std_logic;
signal \N__65827\ : std_logic;
signal \N__65826\ : std_logic;
signal \N__65823\ : std_logic;
signal \N__65820\ : std_logic;
signal \N__65817\ : std_logic;
signal \N__65814\ : std_logic;
signal \N__65811\ : std_logic;
signal \N__65808\ : std_logic;
signal \N__65805\ : std_logic;
signal \N__65802\ : std_logic;
signal \N__65799\ : std_logic;
signal \N__65794\ : std_logic;
signal \N__65789\ : std_logic;
signal \N__65784\ : std_logic;
signal \N__65779\ : std_logic;
signal \N__65774\ : std_logic;
signal \N__65771\ : std_logic;
signal \N__65766\ : std_logic;
signal \N__65759\ : std_logic;
signal \N__65756\ : std_logic;
signal \N__65755\ : std_logic;
signal \N__65754\ : std_logic;
signal \N__65753\ : std_logic;
signal \N__65750\ : std_logic;
signal \N__65743\ : std_logic;
signal \N__65740\ : std_logic;
signal \N__65737\ : std_logic;
signal \N__65734\ : std_logic;
signal \N__65727\ : std_logic;
signal \N__65724\ : std_logic;
signal \N__65721\ : std_logic;
signal \N__65720\ : std_logic;
signal \N__65719\ : std_logic;
signal \N__65718\ : std_logic;
signal \N__65717\ : std_logic;
signal \N__65716\ : std_logic;
signal \N__65715\ : std_logic;
signal \N__65712\ : std_logic;
signal \N__65711\ : std_logic;
signal \N__65710\ : std_logic;
signal \N__65701\ : std_logic;
signal \N__65698\ : std_logic;
signal \N__65695\ : std_logic;
signal \N__65690\ : std_logic;
signal \N__65687\ : std_logic;
signal \N__65676\ : std_logic;
signal \N__65667\ : std_logic;
signal \N__65660\ : std_logic;
signal \N__65655\ : std_logic;
signal \N__65652\ : std_logic;
signal \N__65647\ : std_logic;
signal \N__65642\ : std_logic;
signal \N__65635\ : std_logic;
signal \N__65628\ : std_logic;
signal \N__65619\ : std_logic;
signal \N__65610\ : std_logic;
signal \N__65585\ : std_logic;
signal \N__65584\ : std_logic;
signal \N__65581\ : std_logic;
signal \N__65576\ : std_logic;
signal \N__65575\ : std_logic;
signal \N__65574\ : std_logic;
signal \N__65571\ : std_logic;
signal \N__65570\ : std_logic;
signal \N__65569\ : std_logic;
signal \N__65566\ : std_logic;
signal \N__65565\ : std_logic;
signal \N__65564\ : std_logic;
signal \N__65563\ : std_logic;
signal \N__65562\ : std_logic;
signal \N__65559\ : std_logic;
signal \N__65558\ : std_logic;
signal \N__65557\ : std_logic;
signal \N__65556\ : std_logic;
signal \N__65553\ : std_logic;
signal \N__65552\ : std_logic;
signal \N__65551\ : std_logic;
signal \N__65550\ : std_logic;
signal \N__65547\ : std_logic;
signal \N__65546\ : std_logic;
signal \N__65545\ : std_logic;
signal \N__65544\ : std_logic;
signal \N__65543\ : std_logic;
signal \N__65542\ : std_logic;
signal \N__65541\ : std_logic;
signal \N__65540\ : std_logic;
signal \N__65539\ : std_logic;
signal \N__65538\ : std_logic;
signal \N__65537\ : std_logic;
signal \N__65536\ : std_logic;
signal \N__65531\ : std_logic;
signal \N__65528\ : std_logic;
signal \N__65527\ : std_logic;
signal \N__65526\ : std_logic;
signal \N__65523\ : std_logic;
signal \N__65522\ : std_logic;
signal \N__65521\ : std_logic;
signal \N__65520\ : std_logic;
signal \N__65517\ : std_logic;
signal \N__65514\ : std_logic;
signal \N__65511\ : std_logic;
signal \N__65508\ : std_logic;
signal \N__65505\ : std_logic;
signal \N__65502\ : std_logic;
signal \N__65499\ : std_logic;
signal \N__65494\ : std_logic;
signal \N__65493\ : std_logic;
signal \N__65490\ : std_logic;
signal \N__65487\ : std_logic;
signal \N__65484\ : std_logic;
signal \N__65483\ : std_logic;
signal \N__65482\ : std_logic;
signal \N__65481\ : std_logic;
signal \N__65480\ : std_logic;
signal \N__65479\ : std_logic;
signal \N__65474\ : std_logic;
signal \N__65469\ : std_logic;
signal \N__65464\ : std_logic;
signal \N__65461\ : std_logic;
signal \N__65458\ : std_logic;
signal \N__65455\ : std_logic;
signal \N__65452\ : std_logic;
signal \N__65447\ : std_logic;
signal \N__65446\ : std_logic;
signal \N__65445\ : std_logic;
signal \N__65444\ : std_logic;
signal \N__65439\ : std_logic;
signal \N__65434\ : std_logic;
signal \N__65431\ : std_logic;
signal \N__65428\ : std_logic;
signal \N__65423\ : std_logic;
signal \N__65418\ : std_logic;
signal \N__65409\ : std_logic;
signal \N__65408\ : std_logic;
signal \N__65407\ : std_logic;
signal \N__65404\ : std_logic;
signal \N__65399\ : std_logic;
signal \N__65386\ : std_logic;
signal \N__65379\ : std_logic;
signal \N__65374\ : std_logic;
signal \N__65369\ : std_logic;
signal \N__65366\ : std_logic;
signal \N__65359\ : std_logic;
signal \N__65352\ : std_logic;
signal \N__65351\ : std_logic;
signal \N__65348\ : std_logic;
signal \N__65343\ : std_logic;
signal \N__65340\ : std_logic;
signal \N__65335\ : std_logic;
signal \N__65326\ : std_logic;
signal \N__65319\ : std_logic;
signal \N__65316\ : std_logic;
signal \N__65313\ : std_logic;
signal \N__65310\ : std_logic;
signal \N__65305\ : std_logic;
signal \N__65298\ : std_logic;
signal \N__65285\ : std_logic;
signal \N__65282\ : std_logic;
signal \N__65279\ : std_logic;
signal \N__65276\ : std_logic;
signal \N__65273\ : std_logic;
signal \N__65272\ : std_logic;
signal \N__65269\ : std_logic;
signal \N__65266\ : std_logic;
signal \N__65263\ : std_logic;
signal \N__65260\ : std_logic;
signal \N__65255\ : std_logic;
signal \N__65252\ : std_logic;
signal \N__65249\ : std_logic;
signal \N__65246\ : std_logic;
signal \N__65243\ : std_logic;
signal \N__65240\ : std_logic;
signal \N__65237\ : std_logic;
signal \N__65236\ : std_logic;
signal \N__65233\ : std_logic;
signal \N__65228\ : std_logic;
signal \N__65225\ : std_logic;
signal \N__65222\ : std_logic;
signal \N__65219\ : std_logic;
signal \N__65216\ : std_logic;
signal \N__65213\ : std_logic;
signal \N__65210\ : std_logic;
signal \N__65207\ : std_logic;
signal \N__65204\ : std_logic;
signal \N__65201\ : std_logic;
signal \N__65198\ : std_logic;
signal \N__65195\ : std_logic;
signal \N__65192\ : std_logic;
signal \N__65189\ : std_logic;
signal \N__65186\ : std_logic;
signal \N__65183\ : std_logic;
signal \N__65180\ : std_logic;
signal \N__65177\ : std_logic;
signal \N__65174\ : std_logic;
signal \N__65171\ : std_logic;
signal \N__65168\ : std_logic;
signal \N__65165\ : std_logic;
signal \N__65162\ : std_logic;
signal \N__65159\ : std_logic;
signal \N__65156\ : std_logic;
signal \N__65153\ : std_logic;
signal \N__65150\ : std_logic;
signal \N__65149\ : std_logic;
signal \N__65146\ : std_logic;
signal \N__65143\ : std_logic;
signal \N__65140\ : std_logic;
signal \N__65137\ : std_logic;
signal \N__65134\ : std_logic;
signal \N__65131\ : std_logic;
signal \N__65126\ : std_logic;
signal \N__65123\ : std_logic;
signal \N__65120\ : std_logic;
signal \N__65117\ : std_logic;
signal \N__65114\ : std_logic;
signal \N__65111\ : std_logic;
signal \N__65108\ : std_logic;
signal \N__65105\ : std_logic;
signal \N__65102\ : std_logic;
signal \N__65099\ : std_logic;
signal \N__65096\ : std_logic;
signal \N__65093\ : std_logic;
signal \N__65090\ : std_logic;
signal \N__65089\ : std_logic;
signal \N__65086\ : std_logic;
signal \N__65083\ : std_logic;
signal \N__65078\ : std_logic;
signal \N__65075\ : std_logic;
signal \N__65072\ : std_logic;
signal \N__65069\ : std_logic;
signal \N__65066\ : std_logic;
signal \N__65063\ : std_logic;
signal \N__65060\ : std_logic;
signal \N__65057\ : std_logic;
signal \N__65056\ : std_logic;
signal \N__65053\ : std_logic;
signal \N__65050\ : std_logic;
signal \N__65047\ : std_logic;
signal \N__65044\ : std_logic;
signal \N__65041\ : std_logic;
signal \N__65038\ : std_logic;
signal \N__65033\ : std_logic;
signal \N__65030\ : std_logic;
signal \N__65029\ : std_logic;
signal \N__65026\ : std_logic;
signal \N__65023\ : std_logic;
signal \N__65020\ : std_logic;
signal \N__65017\ : std_logic;
signal \N__65014\ : std_logic;
signal \N__65013\ : std_logic;
signal \N__65010\ : std_logic;
signal \N__65007\ : std_logic;
signal \N__65004\ : std_logic;
signal \N__65001\ : std_logic;
signal \N__64998\ : std_logic;
signal \N__64995\ : std_logic;
signal \N__64992\ : std_logic;
signal \N__64989\ : std_logic;
signal \N__64984\ : std_logic;
signal \N__64981\ : std_logic;
signal \N__64976\ : std_logic;
signal \N__64973\ : std_logic;
signal \N__64970\ : std_logic;
signal \N__64967\ : std_logic;
signal \N__64966\ : std_logic;
signal \N__64965\ : std_logic;
signal \N__64964\ : std_logic;
signal \N__64961\ : std_logic;
signal \N__64958\ : std_logic;
signal \N__64955\ : std_logic;
signal \N__64952\ : std_logic;
signal \N__64949\ : std_logic;
signal \N__64946\ : std_logic;
signal \N__64941\ : std_logic;
signal \N__64940\ : std_logic;
signal \N__64933\ : std_logic;
signal \N__64930\ : std_logic;
signal \N__64925\ : std_logic;
signal \N__64922\ : std_logic;
signal \N__64919\ : std_logic;
signal \N__64916\ : std_logic;
signal \N__64913\ : std_logic;
signal \N__64910\ : std_logic;
signal \N__64907\ : std_logic;
signal \N__64904\ : std_logic;
signal \N__64901\ : std_logic;
signal \N__64900\ : std_logic;
signal \N__64897\ : std_logic;
signal \N__64894\ : std_logic;
signal \N__64891\ : std_logic;
signal \N__64888\ : std_logic;
signal \N__64885\ : std_logic;
signal \N__64882\ : std_logic;
signal \N__64877\ : std_logic;
signal \N__64876\ : std_logic;
signal \N__64875\ : std_logic;
signal \N__64872\ : std_logic;
signal \N__64871\ : std_logic;
signal \N__64870\ : std_logic;
signal \N__64867\ : std_logic;
signal \N__64864\ : std_logic;
signal \N__64863\ : std_logic;
signal \N__64862\ : std_logic;
signal \N__64861\ : std_logic;
signal \N__64858\ : std_logic;
signal \N__64855\ : std_logic;
signal \N__64852\ : std_logic;
signal \N__64849\ : std_logic;
signal \N__64844\ : std_logic;
signal \N__64841\ : std_logic;
signal \N__64838\ : std_logic;
signal \N__64837\ : std_logic;
signal \N__64834\ : std_logic;
signal \N__64831\ : std_logic;
signal \N__64828\ : std_logic;
signal \N__64825\ : std_logic;
signal \N__64822\ : std_logic;
signal \N__64819\ : std_logic;
signal \N__64814\ : std_logic;
signal \N__64809\ : std_logic;
signal \N__64804\ : std_logic;
signal \N__64793\ : std_logic;
signal \N__64790\ : std_logic;
signal \N__64789\ : std_logic;
signal \N__64786\ : std_logic;
signal \N__64783\ : std_logic;
signal \N__64778\ : std_logic;
signal \N__64775\ : std_logic;
signal \N__64772\ : std_logic;
signal \N__64769\ : std_logic;
signal \N__64766\ : std_logic;
signal \N__64763\ : std_logic;
signal \N__64760\ : std_logic;
signal \N__64757\ : std_logic;
signal \N__64754\ : std_logic;
signal \N__64751\ : std_logic;
signal \N__64748\ : std_logic;
signal \N__64747\ : std_logic;
signal \N__64742\ : std_logic;
signal \N__64741\ : std_logic;
signal \N__64740\ : std_logic;
signal \N__64737\ : std_logic;
signal \N__64734\ : std_logic;
signal \N__64731\ : std_logic;
signal \N__64728\ : std_logic;
signal \N__64725\ : std_logic;
signal \N__64722\ : std_logic;
signal \N__64715\ : std_logic;
signal \N__64712\ : std_logic;
signal \N__64711\ : std_logic;
signal \N__64710\ : std_logic;
signal \N__64705\ : std_logic;
signal \N__64702\ : std_logic;
signal \N__64699\ : std_logic;
signal \N__64698\ : std_logic;
signal \N__64695\ : std_logic;
signal \N__64694\ : std_logic;
signal \N__64693\ : std_logic;
signal \N__64692\ : std_logic;
signal \N__64689\ : std_logic;
signal \N__64686\ : std_logic;
signal \N__64683\ : std_logic;
signal \N__64680\ : std_logic;
signal \N__64675\ : std_logic;
signal \N__64664\ : std_logic;
signal \N__64663\ : std_logic;
signal \N__64662\ : std_logic;
signal \N__64659\ : std_logic;
signal \N__64656\ : std_logic;
signal \N__64655\ : std_logic;
signal \N__64652\ : std_logic;
signal \N__64649\ : std_logic;
signal \N__64646\ : std_logic;
signal \N__64643\ : std_logic;
signal \N__64642\ : std_logic;
signal \N__64641\ : std_logic;
signal \N__64638\ : std_logic;
signal \N__64635\ : std_logic;
signal \N__64632\ : std_logic;
signal \N__64629\ : std_logic;
signal \N__64626\ : std_logic;
signal \N__64623\ : std_logic;
signal \N__64620\ : std_logic;
signal \N__64619\ : std_logic;
signal \N__64616\ : std_logic;
signal \N__64611\ : std_logic;
signal \N__64608\ : std_logic;
signal \N__64605\ : std_logic;
signal \N__64602\ : std_logic;
signal \N__64599\ : std_logic;
signal \N__64598\ : std_logic;
signal \N__64597\ : std_logic;
signal \N__64596\ : std_logic;
signal \N__64595\ : std_logic;
signal \N__64594\ : std_logic;
signal \N__64591\ : std_logic;
signal \N__64588\ : std_logic;
signal \N__64583\ : std_logic;
signal \N__64580\ : std_logic;
signal \N__64577\ : std_logic;
signal \N__64574\ : std_logic;
signal \N__64569\ : std_logic;
signal \N__64566\ : std_logic;
signal \N__64563\ : std_logic;
signal \N__64544\ : std_logic;
signal \N__64541\ : std_logic;
signal \N__64538\ : std_logic;
signal \N__64535\ : std_logic;
signal \N__64532\ : std_logic;
signal \N__64531\ : std_logic;
signal \N__64528\ : std_logic;
signal \N__64525\ : std_logic;
signal \N__64524\ : std_logic;
signal \N__64521\ : std_logic;
signal \N__64518\ : std_logic;
signal \N__64515\ : std_logic;
signal \N__64512\ : std_logic;
signal \N__64509\ : std_logic;
signal \N__64506\ : std_logic;
signal \N__64503\ : std_logic;
signal \N__64500\ : std_logic;
signal \N__64497\ : std_logic;
signal \N__64492\ : std_logic;
signal \N__64487\ : std_logic;
signal \N__64486\ : std_logic;
signal \N__64485\ : std_logic;
signal \N__64482\ : std_logic;
signal \N__64479\ : std_logic;
signal \N__64476\ : std_logic;
signal \N__64473\ : std_logic;
signal \N__64470\ : std_logic;
signal \N__64467\ : std_logic;
signal \N__64466\ : std_logic;
signal \N__64465\ : std_logic;
signal \N__64462\ : std_logic;
signal \N__64459\ : std_logic;
signal \N__64456\ : std_logic;
signal \N__64451\ : std_logic;
signal \N__64442\ : std_logic;
signal \N__64439\ : std_logic;
signal \N__64436\ : std_logic;
signal \N__64433\ : std_logic;
signal \N__64430\ : std_logic;
signal \N__64427\ : std_logic;
signal \N__64424\ : std_logic;
signal \N__64421\ : std_logic;
signal \N__64418\ : std_logic;
signal \N__64415\ : std_logic;
signal \N__64412\ : std_logic;
signal \N__64409\ : std_logic;
signal \N__64406\ : std_logic;
signal \N__64403\ : std_logic;
signal \N__64400\ : std_logic;
signal \N__64397\ : std_logic;
signal \N__64396\ : std_logic;
signal \N__64393\ : std_logic;
signal \N__64390\ : std_logic;
signal \N__64387\ : std_logic;
signal \N__64382\ : std_logic;
signal \N__64379\ : std_logic;
signal \N__64376\ : std_logic;
signal \N__64373\ : std_logic;
signal \N__64370\ : std_logic;
signal \N__64367\ : std_logic;
signal \N__64364\ : std_logic;
signal \N__64361\ : std_logic;
signal \N__64358\ : std_logic;
signal \N__64355\ : std_logic;
signal \N__64352\ : std_logic;
signal \N__64349\ : std_logic;
signal \N__64346\ : std_logic;
signal \N__64343\ : std_logic;
signal \N__64340\ : std_logic;
signal \N__64337\ : std_logic;
signal \N__64334\ : std_logic;
signal \N__64331\ : std_logic;
signal \N__64328\ : std_logic;
signal \N__64325\ : std_logic;
signal \N__64324\ : std_logic;
signal \N__64323\ : std_logic;
signal \N__64320\ : std_logic;
signal \N__64317\ : std_logic;
signal \N__64314\ : std_logic;
signal \N__64311\ : std_logic;
signal \N__64308\ : std_logic;
signal \N__64305\ : std_logic;
signal \N__64298\ : std_logic;
signal \N__64295\ : std_logic;
signal \N__64292\ : std_logic;
signal \N__64289\ : std_logic;
signal \N__64286\ : std_logic;
signal \N__64283\ : std_logic;
signal \N__64280\ : std_logic;
signal \N__64277\ : std_logic;
signal \N__64274\ : std_logic;
signal \N__64271\ : std_logic;
signal \N__64268\ : std_logic;
signal \N__64265\ : std_logic;
signal \N__64262\ : std_logic;
signal \N__64261\ : std_logic;
signal \N__64258\ : std_logic;
signal \N__64255\ : std_logic;
signal \N__64254\ : std_logic;
signal \N__64251\ : std_logic;
signal \N__64250\ : std_logic;
signal \N__64247\ : std_logic;
signal \N__64246\ : std_logic;
signal \N__64245\ : std_logic;
signal \N__64242\ : std_logic;
signal \N__64239\ : std_logic;
signal \N__64236\ : std_logic;
signal \N__64235\ : std_logic;
signal \N__64232\ : std_logic;
signal \N__64229\ : std_logic;
signal \N__64226\ : std_logic;
signal \N__64223\ : std_logic;
signal \N__64218\ : std_logic;
signal \N__64215\ : std_logic;
signal \N__64202\ : std_logic;
signal \N__64199\ : std_logic;
signal \N__64196\ : std_logic;
signal \N__64193\ : std_logic;
signal \N__64190\ : std_logic;
signal \N__64187\ : std_logic;
signal \N__64184\ : std_logic;
signal \N__64181\ : std_logic;
signal \N__64178\ : std_logic;
signal \N__64175\ : std_logic;
signal \N__64172\ : std_logic;
signal \N__64169\ : std_logic;
signal \N__64166\ : std_logic;
signal \N__64163\ : std_logic;
signal \N__64160\ : std_logic;
signal \N__64157\ : std_logic;
signal \N__64154\ : std_logic;
signal \N__64151\ : std_logic;
signal \N__64148\ : std_logic;
signal \N__64145\ : std_logic;
signal \N__64142\ : std_logic;
signal \N__64139\ : std_logic;
signal \N__64136\ : std_logic;
signal \N__64133\ : std_logic;
signal \N__64130\ : std_logic;
signal \N__64127\ : std_logic;
signal \N__64124\ : std_logic;
signal \N__64123\ : std_logic;
signal \N__64120\ : std_logic;
signal \N__64117\ : std_logic;
signal \N__64112\ : std_logic;
signal \N__64109\ : std_logic;
signal \N__64108\ : std_logic;
signal \N__64107\ : std_logic;
signal \N__64106\ : std_logic;
signal \N__64105\ : std_logic;
signal \N__64102\ : std_logic;
signal \N__64099\ : std_logic;
signal \N__64092\ : std_logic;
signal \N__64085\ : std_logic;
signal \N__64084\ : std_logic;
signal \N__64083\ : std_logic;
signal \N__64080\ : std_logic;
signal \N__64075\ : std_logic;
signal \N__64070\ : std_logic;
signal \N__64067\ : std_logic;
signal \N__64064\ : std_logic;
signal \N__64061\ : std_logic;
signal \N__64058\ : std_logic;
signal \N__64057\ : std_logic;
signal \N__64054\ : std_logic;
signal \N__64049\ : std_logic;
signal \N__64046\ : std_logic;
signal \N__64043\ : std_logic;
signal \N__64040\ : std_logic;
signal \N__64037\ : std_logic;
signal \N__64034\ : std_logic;
signal \N__64031\ : std_logic;
signal \N__64028\ : std_logic;
signal \N__64025\ : std_logic;
signal \N__64022\ : std_logic;
signal \N__64019\ : std_logic;
signal \N__64018\ : std_logic;
signal \N__64017\ : std_logic;
signal \N__64014\ : std_logic;
signal \N__64011\ : std_logic;
signal \N__64008\ : std_logic;
signal \N__64007\ : std_logic;
signal \N__64004\ : std_logic;
signal \N__64001\ : std_logic;
signal \N__63998\ : std_logic;
signal \N__63995\ : std_logic;
signal \N__63992\ : std_logic;
signal \N__63987\ : std_logic;
signal \N__63984\ : std_logic;
signal \N__63981\ : std_logic;
signal \N__63978\ : std_logic;
signal \N__63975\ : std_logic;
signal \N__63968\ : std_logic;
signal \N__63967\ : std_logic;
signal \N__63964\ : std_logic;
signal \N__63959\ : std_logic;
signal \N__63956\ : std_logic;
signal \N__63953\ : std_logic;
signal \N__63950\ : std_logic;
signal \N__63947\ : std_logic;
signal \N__63944\ : std_logic;
signal \N__63941\ : std_logic;
signal \N__63938\ : std_logic;
signal \N__63935\ : std_logic;
signal \N__63932\ : std_logic;
signal \N__63929\ : std_logic;
signal \N__63926\ : std_logic;
signal \N__63923\ : std_logic;
signal \N__63920\ : std_logic;
signal \N__63917\ : std_logic;
signal \N__63914\ : std_logic;
signal \N__63911\ : std_logic;
signal \N__63908\ : std_logic;
signal \N__63905\ : std_logic;
signal \N__63902\ : std_logic;
signal \N__63899\ : std_logic;
signal \N__63896\ : std_logic;
signal \N__63893\ : std_logic;
signal \N__63890\ : std_logic;
signal \N__63887\ : std_logic;
signal \N__63884\ : std_logic;
signal \N__63881\ : std_logic;
signal \N__63878\ : std_logic;
signal \N__63875\ : std_logic;
signal \N__63872\ : std_logic;
signal \N__63869\ : std_logic;
signal \N__63866\ : std_logic;
signal \N__63863\ : std_logic;
signal \N__63860\ : std_logic;
signal \N__63857\ : std_logic;
signal \N__63854\ : std_logic;
signal \N__63853\ : std_logic;
signal \N__63852\ : std_logic;
signal \N__63849\ : std_logic;
signal \N__63848\ : std_logic;
signal \N__63847\ : std_logic;
signal \N__63844\ : std_logic;
signal \N__63843\ : std_logic;
signal \N__63842\ : std_logic;
signal \N__63839\ : std_logic;
signal \N__63836\ : std_logic;
signal \N__63835\ : std_logic;
signal \N__63832\ : std_logic;
signal \N__63829\ : std_logic;
signal \N__63826\ : std_logic;
signal \N__63823\ : std_logic;
signal \N__63820\ : std_logic;
signal \N__63819\ : std_logic;
signal \N__63816\ : std_logic;
signal \N__63813\ : std_logic;
signal \N__63810\ : std_logic;
signal \N__63809\ : std_logic;
signal \N__63806\ : std_logic;
signal \N__63803\ : std_logic;
signal \N__63802\ : std_logic;
signal \N__63797\ : std_logic;
signal \N__63794\ : std_logic;
signal \N__63791\ : std_logic;
signal \N__63788\ : std_logic;
signal \N__63783\ : std_logic;
signal \N__63780\ : std_logic;
signal \N__63779\ : std_logic;
signal \N__63778\ : std_logic;
signal \N__63775\ : std_logic;
signal \N__63774\ : std_logic;
signal \N__63771\ : std_logic;
signal \N__63768\ : std_logic;
signal \N__63763\ : std_logic;
signal \N__63760\ : std_logic;
signal \N__63753\ : std_logic;
signal \N__63748\ : std_logic;
signal \N__63745\ : std_logic;
signal \N__63742\ : std_logic;
signal \N__63739\ : std_logic;
signal \N__63734\ : std_logic;
signal \N__63731\ : std_logic;
signal \N__63728\ : std_logic;
signal \N__63721\ : std_logic;
signal \N__63716\ : std_logic;
signal \N__63711\ : std_logic;
signal \N__63706\ : std_logic;
signal \N__63701\ : std_logic;
signal \N__63700\ : std_logic;
signal \N__63699\ : std_logic;
signal \N__63694\ : std_logic;
signal \N__63691\ : std_logic;
signal \N__63688\ : std_logic;
signal \N__63683\ : std_logic;
signal \N__63680\ : std_logic;
signal \N__63677\ : std_logic;
signal \N__63674\ : std_logic;
signal \N__63671\ : std_logic;
signal \N__63670\ : std_logic;
signal \N__63669\ : std_logic;
signal \N__63668\ : std_logic;
signal \N__63665\ : std_logic;
signal \N__63662\ : std_logic;
signal \N__63659\ : std_logic;
signal \N__63658\ : std_logic;
signal \N__63655\ : std_logic;
signal \N__63652\ : std_logic;
signal \N__63649\ : std_logic;
signal \N__63646\ : std_logic;
signal \N__63645\ : std_logic;
signal \N__63644\ : std_logic;
signal \N__63641\ : std_logic;
signal \N__63640\ : std_logic;
signal \N__63639\ : std_logic;
signal \N__63638\ : std_logic;
signal \N__63635\ : std_logic;
signal \N__63628\ : std_logic;
signal \N__63625\ : std_logic;
signal \N__63622\ : std_logic;
signal \N__63619\ : std_logic;
signal \N__63616\ : std_logic;
signal \N__63615\ : std_logic;
signal \N__63614\ : std_logic;
signal \N__63613\ : std_logic;
signal \N__63612\ : std_logic;
signal \N__63607\ : std_logic;
signal \N__63598\ : std_logic;
signal \N__63595\ : std_logic;
signal \N__63594\ : std_logic;
signal \N__63593\ : std_logic;
signal \N__63592\ : std_logic;
signal \N__63589\ : std_logic;
signal \N__63586\ : std_logic;
signal \N__63583\ : std_logic;
signal \N__63582\ : std_logic;
signal \N__63579\ : std_logic;
signal \N__63576\ : std_logic;
signal \N__63571\ : std_logic;
signal \N__63568\ : std_logic;
signal \N__63561\ : std_logic;
signal \N__63558\ : std_logic;
signal \N__63555\ : std_logic;
signal \N__63548\ : std_logic;
signal \N__63545\ : std_logic;
signal \N__63542\ : std_logic;
signal \N__63537\ : std_logic;
signal \N__63524\ : std_logic;
signal \N__63523\ : std_logic;
signal \N__63520\ : std_logic;
signal \N__63517\ : std_logic;
signal \N__63516\ : std_logic;
signal \N__63513\ : std_logic;
signal \N__63512\ : std_logic;
signal \N__63509\ : std_logic;
signal \N__63506\ : std_logic;
signal \N__63503\ : std_logic;
signal \N__63500\ : std_logic;
signal \N__63497\ : std_logic;
signal \N__63488\ : std_logic;
signal \N__63485\ : std_logic;
signal \N__63482\ : std_logic;
signal \N__63481\ : std_logic;
signal \N__63478\ : std_logic;
signal \N__63475\ : std_logic;
signal \N__63472\ : std_logic;
signal \N__63469\ : std_logic;
signal \N__63464\ : std_logic;
signal \N__63463\ : std_logic;
signal \N__63462\ : std_logic;
signal \N__63461\ : std_logic;
signal \N__63460\ : std_logic;
signal \N__63459\ : std_logic;
signal \N__63456\ : std_logic;
signal \N__63453\ : std_logic;
signal \N__63448\ : std_logic;
signal \N__63443\ : std_logic;
signal \N__63442\ : std_logic;
signal \N__63435\ : std_logic;
signal \N__63432\ : std_logic;
signal \N__63429\ : std_logic;
signal \N__63426\ : std_logic;
signal \N__63423\ : std_logic;
signal \N__63418\ : std_logic;
signal \N__63415\ : std_logic;
signal \N__63414\ : std_logic;
signal \N__63411\ : std_logic;
signal \N__63408\ : std_logic;
signal \N__63405\ : std_logic;
signal \N__63402\ : std_logic;
signal \N__63399\ : std_logic;
signal \N__63392\ : std_logic;
signal \N__63389\ : std_logic;
signal \N__63386\ : std_logic;
signal \N__63383\ : std_logic;
signal \N__63380\ : std_logic;
signal \N__63377\ : std_logic;
signal \N__63374\ : std_logic;
signal \N__63371\ : std_logic;
signal \N__63370\ : std_logic;
signal \N__63367\ : std_logic;
signal \N__63364\ : std_logic;
signal \N__63361\ : std_logic;
signal \N__63360\ : std_logic;
signal \N__63357\ : std_logic;
signal \N__63354\ : std_logic;
signal \N__63351\ : std_logic;
signal \N__63348\ : std_logic;
signal \N__63343\ : std_logic;
signal \N__63340\ : std_logic;
signal \N__63337\ : std_logic;
signal \N__63334\ : std_logic;
signal \N__63331\ : std_logic;
signal \N__63328\ : std_logic;
signal \N__63325\ : std_logic;
signal \N__63320\ : std_logic;
signal \N__63319\ : std_logic;
signal \N__63314\ : std_logic;
signal \N__63311\ : std_logic;
signal \N__63308\ : std_logic;
signal \N__63305\ : std_logic;
signal \N__63302\ : std_logic;
signal \N__63301\ : std_logic;
signal \N__63300\ : std_logic;
signal \N__63299\ : std_logic;
signal \N__63298\ : std_logic;
signal \N__63297\ : std_logic;
signal \N__63294\ : std_logic;
signal \N__63293\ : std_logic;
signal \N__63292\ : std_logic;
signal \N__63291\ : std_logic;
signal \N__63290\ : std_logic;
signal \N__63289\ : std_logic;
signal \N__63280\ : std_logic;
signal \N__63277\ : std_logic;
signal \N__63276\ : std_logic;
signal \N__63275\ : std_logic;
signal \N__63274\ : std_logic;
signal \N__63273\ : std_logic;
signal \N__63270\ : std_logic;
signal \N__63269\ : std_logic;
signal \N__63266\ : std_logic;
signal \N__63265\ : std_logic;
signal \N__63262\ : std_logic;
signal \N__63261\ : std_logic;
signal \N__63260\ : std_logic;
signal \N__63257\ : std_logic;
signal \N__63256\ : std_logic;
signal \N__63255\ : std_logic;
signal \N__63254\ : std_logic;
signal \N__63253\ : std_logic;
signal \N__63250\ : std_logic;
signal \N__63249\ : std_logic;
signal \N__63248\ : std_logic;
signal \N__63247\ : std_logic;
signal \N__63246\ : std_logic;
signal \N__63243\ : std_logic;
signal \N__63242\ : std_logic;
signal \N__63241\ : std_logic;
signal \N__63240\ : std_logic;
signal \N__63239\ : std_logic;
signal \N__63238\ : std_logic;
signal \N__63235\ : std_logic;
signal \N__63232\ : std_logic;
signal \N__63229\ : std_logic;
signal \N__63226\ : std_logic;
signal \N__63225\ : std_logic;
signal \N__63222\ : std_logic;
signal \N__63219\ : std_logic;
signal \N__63218\ : std_logic;
signal \N__63217\ : std_logic;
signal \N__63214\ : std_logic;
signal \N__63209\ : std_logic;
signal \N__63204\ : std_logic;
signal \N__63199\ : std_logic;
signal \N__63196\ : std_logic;
signal \N__63193\ : std_logic;
signal \N__63188\ : std_logic;
signal \N__63185\ : std_logic;
signal \N__63178\ : std_logic;
signal \N__63173\ : std_logic;
signal \N__63170\ : std_logic;
signal \N__63163\ : std_logic;
signal \N__63158\ : std_logic;
signal \N__63151\ : std_logic;
signal \N__63150\ : std_logic;
signal \N__63147\ : std_logic;
signal \N__63142\ : std_logic;
signal \N__63135\ : std_logic;
signal \N__63132\ : std_logic;
signal \N__63125\ : std_logic;
signal \N__63122\ : std_logic;
signal \N__63117\ : std_logic;
signal \N__63116\ : std_logic;
signal \N__63115\ : std_logic;
signal \N__63114\ : std_logic;
signal \N__63113\ : std_logic;
signal \N__63112\ : std_logic;
signal \N__63109\ : std_logic;
signal \N__63106\ : std_logic;
signal \N__63103\ : std_logic;
signal \N__63100\ : std_logic;
signal \N__63093\ : std_logic;
signal \N__63090\ : std_logic;
signal \N__63087\ : std_logic;
signal \N__63082\ : std_logic;
signal \N__63077\ : std_logic;
signal \N__63076\ : std_logic;
signal \N__63075\ : std_logic;
signal \N__63070\ : std_logic;
signal \N__63067\ : std_logic;
signal \N__63062\ : std_logic;
signal \N__63059\ : std_logic;
signal \N__63056\ : std_logic;
signal \N__63053\ : std_logic;
signal \N__63050\ : std_logic;
signal \N__63047\ : std_logic;
signal \N__63044\ : std_logic;
signal \N__63041\ : std_logic;
signal \N__63036\ : std_logic;
signal \N__63031\ : std_logic;
signal \N__63030\ : std_logic;
signal \N__63027\ : std_logic;
signal \N__63026\ : std_logic;
signal \N__63023\ : std_logic;
signal \N__63022\ : std_logic;
signal \N__63009\ : std_logic;
signal \N__63004\ : std_logic;
signal \N__63001\ : std_logic;
signal \N__62998\ : std_logic;
signal \N__62993\ : std_logic;
signal \N__62986\ : std_logic;
signal \N__62981\ : std_logic;
signal \N__62978\ : std_logic;
signal \N__62973\ : std_logic;
signal \N__62968\ : std_logic;
signal \N__62957\ : std_logic;
signal \N__62956\ : std_logic;
signal \N__62953\ : std_logic;
signal \N__62950\ : std_logic;
signal \N__62949\ : std_logic;
signal \N__62946\ : std_logic;
signal \N__62943\ : std_logic;
signal \N__62940\ : std_logic;
signal \N__62939\ : std_logic;
signal \N__62936\ : std_logic;
signal \N__62933\ : std_logic;
signal \N__62928\ : std_logic;
signal \N__62927\ : std_logic;
signal \N__62922\ : std_logic;
signal \N__62919\ : std_logic;
signal \N__62916\ : std_logic;
signal \N__62913\ : std_logic;
signal \N__62910\ : std_logic;
signal \N__62907\ : std_logic;
signal \N__62904\ : std_logic;
signal \N__62899\ : std_logic;
signal \N__62894\ : std_logic;
signal \N__62891\ : std_logic;
signal \N__62890\ : std_logic;
signal \N__62889\ : std_logic;
signal \N__62888\ : std_logic;
signal \N__62887\ : std_logic;
signal \N__62886\ : std_logic;
signal \N__62885\ : std_logic;
signal \N__62884\ : std_logic;
signal \N__62883\ : std_logic;
signal \N__62882\ : std_logic;
signal \N__62881\ : std_logic;
signal \N__62878\ : std_logic;
signal \N__62875\ : std_logic;
signal \N__62874\ : std_logic;
signal \N__62873\ : std_logic;
signal \N__62872\ : std_logic;
signal \N__62871\ : std_logic;
signal \N__62868\ : std_logic;
signal \N__62863\ : std_logic;
signal \N__62860\ : std_logic;
signal \N__62859\ : std_logic;
signal \N__62856\ : std_logic;
signal \N__62849\ : std_logic;
signal \N__62846\ : std_logic;
signal \N__62845\ : std_logic;
signal \N__62842\ : std_logic;
signal \N__62839\ : std_logic;
signal \N__62836\ : std_logic;
signal \N__62833\ : std_logic;
signal \N__62830\ : std_logic;
signal \N__62829\ : std_logic;
signal \N__62826\ : std_logic;
signal \N__62821\ : std_logic;
signal \N__62820\ : std_logic;
signal \N__62819\ : std_logic;
signal \N__62818\ : std_logic;
signal \N__62815\ : std_logic;
signal \N__62812\ : std_logic;
signal \N__62811\ : std_logic;
signal \N__62806\ : std_logic;
signal \N__62805\ : std_logic;
signal \N__62802\ : std_logic;
signal \N__62801\ : std_logic;
signal \N__62798\ : std_logic;
signal \N__62793\ : std_logic;
signal \N__62786\ : std_logic;
signal \N__62785\ : std_logic;
signal \N__62782\ : std_logic;
signal \N__62777\ : std_logic;
signal \N__62774\ : std_logic;
signal \N__62769\ : std_logic;
signal \N__62766\ : std_logic;
signal \N__62765\ : std_logic;
signal \N__62764\ : std_logic;
signal \N__62761\ : std_logic;
signal \N__62758\ : std_logic;
signal \N__62755\ : std_logic;
signal \N__62752\ : std_logic;
signal \N__62749\ : std_logic;
signal \N__62746\ : std_logic;
signal \N__62739\ : std_logic;
signal \N__62736\ : std_logic;
signal \N__62733\ : std_logic;
signal \N__62726\ : std_logic;
signal \N__62723\ : std_logic;
signal \N__62718\ : std_logic;
signal \N__62709\ : std_logic;
signal \N__62704\ : std_logic;
signal \N__62701\ : std_logic;
signal \N__62698\ : std_logic;
signal \N__62693\ : std_logic;
signal \N__62688\ : std_logic;
signal \N__62685\ : std_logic;
signal \N__62672\ : std_logic;
signal \N__62669\ : std_logic;
signal \N__62666\ : std_logic;
signal \N__62663\ : std_logic;
signal \N__62660\ : std_logic;
signal \N__62657\ : std_logic;
signal \N__62656\ : std_logic;
signal \N__62655\ : std_logic;
signal \N__62652\ : std_logic;
signal \N__62649\ : std_logic;
signal \N__62648\ : std_logic;
signal \N__62645\ : std_logic;
signal \N__62642\ : std_logic;
signal \N__62639\ : std_logic;
signal \N__62636\ : std_logic;
signal \N__62627\ : std_logic;
signal \N__62624\ : std_logic;
signal \N__62621\ : std_logic;
signal \N__62618\ : std_logic;
signal \N__62615\ : std_logic;
signal \N__62612\ : std_logic;
signal \N__62609\ : std_logic;
signal \N__62608\ : std_logic;
signal \N__62603\ : std_logic;
signal \N__62600\ : std_logic;
signal \N__62597\ : std_logic;
signal \N__62594\ : std_logic;
signal \N__62591\ : std_logic;
signal \N__62588\ : std_logic;
signal \N__62587\ : std_logic;
signal \N__62586\ : std_logic;
signal \N__62585\ : std_logic;
signal \N__62584\ : std_logic;
signal \N__62583\ : std_logic;
signal \N__62580\ : std_logic;
signal \N__62579\ : std_logic;
signal \N__62576\ : std_logic;
signal \N__62573\ : std_logic;
signal \N__62572\ : std_logic;
signal \N__62571\ : std_logic;
signal \N__62570\ : std_logic;
signal \N__62567\ : std_logic;
signal \N__62564\ : std_logic;
signal \N__62559\ : std_logic;
signal \N__62558\ : std_logic;
signal \N__62557\ : std_logic;
signal \N__62556\ : std_logic;
signal \N__62553\ : std_logic;
signal \N__62552\ : std_logic;
signal \N__62551\ : std_logic;
signal \N__62550\ : std_logic;
signal \N__62547\ : std_logic;
signal \N__62544\ : std_logic;
signal \N__62541\ : std_logic;
signal \N__62538\ : std_logic;
signal \N__62535\ : std_logic;
signal \N__62530\ : std_logic;
signal \N__62527\ : std_logic;
signal \N__62524\ : std_logic;
signal \N__62523\ : std_logic;
signal \N__62520\ : std_logic;
signal \N__62519\ : std_logic;
signal \N__62518\ : std_logic;
signal \N__62515\ : std_logic;
signal \N__62512\ : std_logic;
signal \N__62507\ : std_logic;
signal \N__62506\ : std_logic;
signal \N__62505\ : std_logic;
signal \N__62504\ : std_logic;
signal \N__62503\ : std_logic;
signal \N__62502\ : std_logic;
signal \N__62499\ : std_logic;
signal \N__62496\ : std_logic;
signal \N__62493\ : std_logic;
signal \N__62490\ : std_logic;
signal \N__62487\ : std_logic;
signal \N__62482\ : std_logic;
signal \N__62479\ : std_logic;
signal \N__62476\ : std_logic;
signal \N__62473\ : std_logic;
signal \N__62468\ : std_logic;
signal \N__62465\ : std_logic;
signal \N__62462\ : std_logic;
signal \N__62459\ : std_logic;
signal \N__62456\ : std_logic;
signal \N__62447\ : std_logic;
signal \N__62444\ : std_logic;
signal \N__62441\ : std_logic;
signal \N__62436\ : std_logic;
signal \N__62433\ : std_logic;
signal \N__62430\ : std_logic;
signal \N__62427\ : std_logic;
signal \N__62422\ : std_logic;
signal \N__62417\ : std_logic;
signal \N__62414\ : std_logic;
signal \N__62411\ : std_logic;
signal \N__62402\ : std_logic;
signal \N__62399\ : std_logic;
signal \N__62392\ : std_logic;
signal \N__62389\ : std_logic;
signal \N__62382\ : std_logic;
signal \N__62377\ : std_logic;
signal \N__62366\ : std_logic;
signal \N__62363\ : std_logic;
signal \N__62360\ : std_logic;
signal \N__62357\ : std_logic;
signal \N__62354\ : std_logic;
signal \N__62351\ : std_logic;
signal \N__62348\ : std_logic;
signal \N__62345\ : std_logic;
signal \N__62342\ : std_logic;
signal \N__62339\ : std_logic;
signal \N__62338\ : std_logic;
signal \N__62335\ : std_logic;
signal \N__62332\ : std_logic;
signal \N__62327\ : std_logic;
signal \N__62324\ : std_logic;
signal \N__62321\ : std_logic;
signal \N__62320\ : std_logic;
signal \N__62317\ : std_logic;
signal \N__62316\ : std_logic;
signal \N__62315\ : std_logic;
signal \N__62314\ : std_logic;
signal \N__62311\ : std_logic;
signal \N__62308\ : std_logic;
signal \N__62307\ : std_logic;
signal \N__62306\ : std_logic;
signal \N__62303\ : std_logic;
signal \N__62302\ : std_logic;
signal \N__62299\ : std_logic;
signal \N__62298\ : std_logic;
signal \N__62295\ : std_logic;
signal \N__62292\ : std_logic;
signal \N__62289\ : std_logic;
signal \N__62286\ : std_logic;
signal \N__62285\ : std_logic;
signal \N__62282\ : std_logic;
signal \N__62281\ : std_logic;
signal \N__62278\ : std_logic;
signal \N__62275\ : std_logic;
signal \N__62274\ : std_logic;
signal \N__62273\ : std_logic;
signal \N__62272\ : std_logic;
signal \N__62271\ : std_logic;
signal \N__62270\ : std_logic;
signal \N__62269\ : std_logic;
signal \N__62266\ : std_logic;
signal \N__62265\ : std_logic;
signal \N__62262\ : std_logic;
signal \N__62261\ : std_logic;
signal \N__62256\ : std_logic;
signal \N__62251\ : std_logic;
signal \N__62244\ : std_logic;
signal \N__62241\ : std_logic;
signal \N__62238\ : std_logic;
signal \N__62235\ : std_logic;
signal \N__62234\ : std_logic;
signal \N__62233\ : std_logic;
signal \N__62232\ : std_logic;
signal \N__62223\ : std_logic;
signal \N__62220\ : std_logic;
signal \N__62219\ : std_logic;
signal \N__62216\ : std_logic;
signal \N__62213\ : std_logic;
signal \N__62210\ : std_logic;
signal \N__62209\ : std_logic;
signal \N__62206\ : std_logic;
signal \N__62199\ : std_logic;
signal \N__62192\ : std_logic;
signal \N__62191\ : std_logic;
signal \N__62190\ : std_logic;
signal \N__62187\ : std_logic;
signal \N__62186\ : std_logic;
signal \N__62185\ : std_logic;
signal \N__62182\ : std_logic;
signal \N__62179\ : std_logic;
signal \N__62176\ : std_logic;
signal \N__62173\ : std_logic;
signal \N__62170\ : std_logic;
signal \N__62165\ : std_logic;
signal \N__62162\ : std_logic;
signal \N__62159\ : std_logic;
signal \N__62158\ : std_logic;
signal \N__62157\ : std_logic;
signal \N__62156\ : std_logic;
signal \N__62151\ : std_logic;
signal \N__62148\ : std_logic;
signal \N__62143\ : std_logic;
signal \N__62138\ : std_logic;
signal \N__62135\ : std_logic;
signal \N__62132\ : std_logic;
signal \N__62125\ : std_logic;
signal \N__62122\ : std_logic;
signal \N__62119\ : std_logic;
signal \N__62114\ : std_logic;
signal \N__62107\ : std_logic;
signal \N__62100\ : std_logic;
signal \N__62095\ : std_logic;
signal \N__62090\ : std_logic;
signal \N__62087\ : std_logic;
signal \N__62084\ : std_logic;
signal \N__62079\ : std_logic;
signal \N__62076\ : std_logic;
signal \N__62071\ : std_logic;
signal \N__62060\ : std_logic;
signal \N__62057\ : std_logic;
signal \N__62054\ : std_logic;
signal \N__62051\ : std_logic;
signal \N__62048\ : std_logic;
signal \N__62047\ : std_logic;
signal \N__62044\ : std_logic;
signal \N__62041\ : std_logic;
signal \N__62038\ : std_logic;
signal \N__62035\ : std_logic;
signal \N__62030\ : std_logic;
signal \N__62027\ : std_logic;
signal \N__62026\ : std_logic;
signal \N__62025\ : std_logic;
signal \N__62024\ : std_logic;
signal \N__62023\ : std_logic;
signal \N__62022\ : std_logic;
signal \N__62021\ : std_logic;
signal \N__62018\ : std_logic;
signal \N__62017\ : std_logic;
signal \N__62014\ : std_logic;
signal \N__62011\ : std_logic;
signal \N__62010\ : std_logic;
signal \N__62007\ : std_logic;
signal \N__62004\ : std_logic;
signal \N__62001\ : std_logic;
signal \N__62000\ : std_logic;
signal \N__61997\ : std_logic;
signal \N__61994\ : std_logic;
signal \N__61991\ : std_logic;
signal \N__61984\ : std_logic;
signal \N__61983\ : std_logic;
signal \N__61982\ : std_logic;
signal \N__61979\ : std_logic;
signal \N__61978\ : std_logic;
signal \N__61977\ : std_logic;
signal \N__61976\ : std_logic;
signal \N__61975\ : std_logic;
signal \N__61972\ : std_logic;
signal \N__61969\ : std_logic;
signal \N__61966\ : std_logic;
signal \N__61963\ : std_logic;
signal \N__61960\ : std_logic;
signal \N__61955\ : std_logic;
signal \N__61952\ : std_logic;
signal \N__61949\ : std_logic;
signal \N__61948\ : std_logic;
signal \N__61947\ : std_logic;
signal \N__61944\ : std_logic;
signal \N__61939\ : std_logic;
signal \N__61936\ : std_logic;
signal \N__61935\ : std_logic;
signal \N__61932\ : std_logic;
signal \N__61931\ : std_logic;
signal \N__61930\ : std_logic;
signal \N__61925\ : std_logic;
signal \N__61922\ : std_logic;
signal \N__61919\ : std_logic;
signal \N__61914\ : std_logic;
signal \N__61911\ : std_logic;
signal \N__61908\ : std_logic;
signal \N__61905\ : std_logic;
signal \N__61902\ : std_logic;
signal \N__61901\ : std_logic;
signal \N__61896\ : std_logic;
signal \N__61893\ : std_logic;
signal \N__61890\ : std_logic;
signal \N__61887\ : std_logic;
signal \N__61882\ : std_logic;
signal \N__61881\ : std_logic;
signal \N__61878\ : std_logic;
signal \N__61869\ : std_logic;
signal \N__61866\ : std_logic;
signal \N__61863\ : std_logic;
signal \N__61860\ : std_logic;
signal \N__61857\ : std_logic;
signal \N__61852\ : std_logic;
signal \N__61849\ : std_logic;
signal \N__61846\ : std_logic;
signal \N__61843\ : std_logic;
signal \N__61840\ : std_logic;
signal \N__61837\ : std_logic;
signal \N__61836\ : std_logic;
signal \N__61833\ : std_logic;
signal \N__61830\ : std_logic;
signal \N__61827\ : std_logic;
signal \N__61820\ : std_logic;
signal \N__61817\ : std_logic;
signal \N__61812\ : std_logic;
signal \N__61807\ : std_logic;
signal \N__61804\ : std_logic;
signal \N__61799\ : std_logic;
signal \N__61794\ : std_logic;
signal \N__61781\ : std_logic;
signal \N__61778\ : std_logic;
signal \N__61775\ : std_logic;
signal \N__61772\ : std_logic;
signal \N__61769\ : std_logic;
signal \N__61766\ : std_logic;
signal \N__61763\ : std_logic;
signal \N__61760\ : std_logic;
signal \N__61757\ : std_logic;
signal \N__61754\ : std_logic;
signal \N__61753\ : std_logic;
signal \N__61750\ : std_logic;
signal \N__61747\ : std_logic;
signal \N__61742\ : std_logic;
signal \N__61739\ : std_logic;
signal \N__61736\ : std_logic;
signal \N__61733\ : std_logic;
signal \N__61730\ : std_logic;
signal \N__61727\ : std_logic;
signal \N__61724\ : std_logic;
signal \N__61721\ : std_logic;
signal \N__61718\ : std_logic;
signal \N__61717\ : std_logic;
signal \N__61716\ : std_logic;
signal \N__61715\ : std_logic;
signal \N__61714\ : std_logic;
signal \N__61711\ : std_logic;
signal \N__61710\ : std_logic;
signal \N__61707\ : std_logic;
signal \N__61704\ : std_logic;
signal \N__61703\ : std_logic;
signal \N__61702\ : std_logic;
signal \N__61701\ : std_logic;
signal \N__61698\ : std_logic;
signal \N__61697\ : std_logic;
signal \N__61692\ : std_logic;
signal \N__61689\ : std_logic;
signal \N__61686\ : std_logic;
signal \N__61683\ : std_logic;
signal \N__61682\ : std_logic;
signal \N__61681\ : std_logic;
signal \N__61676\ : std_logic;
signal \N__61675\ : std_logic;
signal \N__61672\ : std_logic;
signal \N__61669\ : std_logic;
signal \N__61668\ : std_logic;
signal \N__61667\ : std_logic;
signal \N__61666\ : std_logic;
signal \N__61663\ : std_logic;
signal \N__61662\ : std_logic;
signal \N__61661\ : std_logic;
signal \N__61658\ : std_logic;
signal \N__61655\ : std_logic;
signal \N__61650\ : std_logic;
signal \N__61647\ : std_logic;
signal \N__61644\ : std_logic;
signal \N__61641\ : std_logic;
signal \N__61640\ : std_logic;
signal \N__61637\ : std_logic;
signal \N__61636\ : std_logic;
signal \N__61633\ : std_logic;
signal \N__61630\ : std_logic;
signal \N__61627\ : std_logic;
signal \N__61624\ : std_logic;
signal \N__61621\ : std_logic;
signal \N__61618\ : std_logic;
signal \N__61613\ : std_logic;
signal \N__61610\ : std_logic;
signal \N__61607\ : std_logic;
signal \N__61604\ : std_logic;
signal \N__61599\ : std_logic;
signal \N__61596\ : std_logic;
signal \N__61593\ : std_logic;
signal \N__61588\ : std_logic;
signal \N__61583\ : std_logic;
signal \N__61580\ : std_logic;
signal \N__61577\ : std_logic;
signal \N__61574\ : std_logic;
signal \N__61571\ : std_logic;
signal \N__61568\ : std_logic;
signal \N__61565\ : std_logic;
signal \N__61562\ : std_logic;
signal \N__61559\ : std_logic;
signal \N__61556\ : std_logic;
signal \N__61553\ : std_logic;
signal \N__61546\ : std_logic;
signal \N__61541\ : std_logic;
signal \N__61536\ : std_logic;
signal \N__61533\ : std_logic;
signal \N__61526\ : std_logic;
signal \N__61521\ : std_logic;
signal \N__61516\ : std_logic;
signal \N__61505\ : std_logic;
signal \N__61502\ : std_logic;
signal \N__61499\ : std_logic;
signal \N__61496\ : std_logic;
signal \N__61493\ : std_logic;
signal \N__61492\ : std_logic;
signal \N__61489\ : std_logic;
signal \N__61486\ : std_logic;
signal \N__61483\ : std_logic;
signal \N__61478\ : std_logic;
signal \N__61475\ : std_logic;
signal \N__61474\ : std_logic;
signal \N__61473\ : std_logic;
signal \N__61472\ : std_logic;
signal \N__61471\ : std_logic;
signal \N__61470\ : std_logic;
signal \N__61467\ : std_logic;
signal \N__61466\ : std_logic;
signal \N__61465\ : std_logic;
signal \N__61464\ : std_logic;
signal \N__61463\ : std_logic;
signal \N__61462\ : std_logic;
signal \N__61461\ : std_logic;
signal \N__61460\ : std_logic;
signal \N__61457\ : std_logic;
signal \N__61454\ : std_logic;
signal \N__61447\ : std_logic;
signal \N__61446\ : std_logic;
signal \N__61443\ : std_logic;
signal \N__61440\ : std_logic;
signal \N__61439\ : std_logic;
signal \N__61436\ : std_logic;
signal \N__61435\ : std_logic;
signal \N__61434\ : std_logic;
signal \N__61433\ : std_logic;
signal \N__61428\ : std_logic;
signal \N__61427\ : std_logic;
signal \N__61426\ : std_logic;
signal \N__61425\ : std_logic;
signal \N__61422\ : std_logic;
signal \N__61417\ : std_logic;
signal \N__61410\ : std_logic;
signal \N__61407\ : std_logic;
signal \N__61404\ : std_logic;
signal \N__61401\ : std_logic;
signal \N__61398\ : std_logic;
signal \N__61395\ : std_logic;
signal \N__61390\ : std_logic;
signal \N__61387\ : std_logic;
signal \N__61384\ : std_logic;
signal \N__61381\ : std_logic;
signal \N__61378\ : std_logic;
signal \N__61375\ : std_logic;
signal \N__61372\ : std_logic;
signal \N__61365\ : std_logic;
signal \N__61364\ : std_logic;
signal \N__61353\ : std_logic;
signal \N__61350\ : std_logic;
signal \N__61347\ : std_logic;
signal \N__61344\ : std_logic;
signal \N__61341\ : std_logic;
signal \N__61334\ : std_logic;
signal \N__61331\ : std_logic;
signal \N__61328\ : std_logic;
signal \N__61325\ : std_logic;
signal \N__61322\ : std_logic;
signal \N__61317\ : std_logic;
signal \N__61314\ : std_logic;
signal \N__61309\ : std_logic;
signal \N__61298\ : std_logic;
signal \N__61295\ : std_logic;
signal \N__61292\ : std_logic;
signal \N__61289\ : std_logic;
signal \N__61286\ : std_logic;
signal \N__61283\ : std_logic;
signal \N__61280\ : std_logic;
signal \N__61277\ : std_logic;
signal \N__61276\ : std_logic;
signal \N__61273\ : std_logic;
signal \N__61270\ : std_logic;
signal \N__61267\ : std_logic;
signal \N__61264\ : std_logic;
signal \N__61261\ : std_logic;
signal \N__61258\ : std_logic;
signal \N__61255\ : std_logic;
signal \N__61252\ : std_logic;
signal \N__61247\ : std_logic;
signal \N__61244\ : std_logic;
signal \N__61241\ : std_logic;
signal \N__61238\ : std_logic;
signal \N__61235\ : std_logic;
signal \N__61232\ : std_logic;
signal \N__61229\ : std_logic;
signal \N__61226\ : std_logic;
signal \N__61225\ : std_logic;
signal \N__61224\ : std_logic;
signal \N__61221\ : std_logic;
signal \N__61218\ : std_logic;
signal \N__61217\ : std_logic;
signal \N__61216\ : std_logic;
signal \N__61213\ : std_logic;
signal \N__61212\ : std_logic;
signal \N__61211\ : std_logic;
signal \N__61210\ : std_logic;
signal \N__61207\ : std_logic;
signal \N__61204\ : std_logic;
signal \N__61203\ : std_logic;
signal \N__61200\ : std_logic;
signal \N__61199\ : std_logic;
signal \N__61196\ : std_logic;
signal \N__61195\ : std_logic;
signal \N__61194\ : std_logic;
signal \N__61193\ : std_logic;
signal \N__61190\ : std_logic;
signal \N__61187\ : std_logic;
signal \N__61184\ : std_logic;
signal \N__61181\ : std_logic;
signal \N__61176\ : std_logic;
signal \N__61171\ : std_logic;
signal \N__61170\ : std_logic;
signal \N__61167\ : std_logic;
signal \N__61164\ : std_logic;
signal \N__61161\ : std_logic;
signal \N__61158\ : std_logic;
signal \N__61157\ : std_logic;
signal \N__61156\ : std_logic;
signal \N__61153\ : std_logic;
signal \N__61152\ : std_logic;
signal \N__61151\ : std_logic;
signal \N__61148\ : std_logic;
signal \N__61143\ : std_logic;
signal \N__61140\ : std_logic;
signal \N__61135\ : std_logic;
signal \N__61132\ : std_logic;
signal \N__61129\ : std_logic;
signal \N__61126\ : std_logic;
signal \N__61123\ : std_logic;
signal \N__61120\ : std_logic;
signal \N__61115\ : std_logic;
signal \N__61112\ : std_logic;
signal \N__61107\ : std_logic;
signal \N__61104\ : std_logic;
signal \N__61101\ : std_logic;
signal \N__61094\ : std_logic;
signal \N__61091\ : std_logic;
signal \N__61082\ : std_logic;
signal \N__61079\ : std_logic;
signal \N__61076\ : std_logic;
signal \N__61071\ : std_logic;
signal \N__61068\ : std_logic;
signal \N__61063\ : std_logic;
signal \N__61058\ : std_logic;
signal \N__61053\ : std_logic;
signal \N__61050\ : std_logic;
signal \N__61043\ : std_logic;
signal \N__61042\ : std_logic;
signal \N__61037\ : std_logic;
signal \N__61034\ : std_logic;
signal \N__61031\ : std_logic;
signal \N__61028\ : std_logic;
signal \N__61025\ : std_logic;
signal \N__61022\ : std_logic;
signal \N__61019\ : std_logic;
signal \N__61018\ : std_logic;
signal \N__61015\ : std_logic;
signal \N__61014\ : std_logic;
signal \N__61013\ : std_logic;
signal \N__61012\ : std_logic;
signal \N__61011\ : std_logic;
signal \N__61010\ : std_logic;
signal \N__61009\ : std_logic;
signal \N__61008\ : std_logic;
signal \N__61005\ : std_logic;
signal \N__61002\ : std_logic;
signal \N__60999\ : std_logic;
signal \N__60996\ : std_logic;
signal \N__60995\ : std_logic;
signal \N__60994\ : std_logic;
signal \N__60991\ : std_logic;
signal \N__60990\ : std_logic;
signal \N__60987\ : std_logic;
signal \N__60984\ : std_logic;
signal \N__60979\ : std_logic;
signal \N__60972\ : std_logic;
signal \N__60969\ : std_logic;
signal \N__60966\ : std_logic;
signal \N__60965\ : std_logic;
signal \N__60964\ : std_logic;
signal \N__60961\ : std_logic;
signal \N__60958\ : std_logic;
signal \N__60955\ : std_logic;
signal \N__60954\ : std_logic;
signal \N__60953\ : std_logic;
signal \N__60950\ : std_logic;
signal \N__60947\ : std_logic;
signal \N__60944\ : std_logic;
signal \N__60941\ : std_logic;
signal \N__60940\ : std_logic;
signal \N__60939\ : std_logic;
signal \N__60938\ : std_logic;
signal \N__60933\ : std_logic;
signal \N__60928\ : std_logic;
signal \N__60925\ : std_logic;
signal \N__60920\ : std_logic;
signal \N__60917\ : std_logic;
signal \N__60914\ : std_logic;
signal \N__60911\ : std_logic;
signal \N__60906\ : std_logic;
signal \N__60903\ : std_logic;
signal \N__60896\ : std_logic;
signal \N__60893\ : std_logic;
signal \N__60890\ : std_logic;
signal \N__60887\ : std_logic;
signal \N__60884\ : std_logic;
signal \N__60879\ : std_logic;
signal \N__60870\ : std_logic;
signal \N__60867\ : std_logic;
signal \N__60864\ : std_logic;
signal \N__60861\ : std_logic;
signal \N__60858\ : std_logic;
signal \N__60853\ : std_logic;
signal \N__60848\ : std_logic;
signal \N__60839\ : std_logic;
signal \N__60836\ : std_logic;
signal \N__60835\ : std_logic;
signal \N__60832\ : std_logic;
signal \N__60829\ : std_logic;
signal \N__60826\ : std_logic;
signal \N__60823\ : std_logic;
signal \N__60818\ : std_logic;
signal \N__60815\ : std_logic;
signal \N__60814\ : std_logic;
signal \N__60813\ : std_logic;
signal \N__60812\ : std_logic;
signal \N__60809\ : std_logic;
signal \N__60806\ : std_logic;
signal \N__60805\ : std_logic;
signal \N__60802\ : std_logic;
signal \N__60799\ : std_logic;
signal \N__60796\ : std_logic;
signal \N__60793\ : std_logic;
signal \N__60790\ : std_logic;
signal \N__60787\ : std_logic;
signal \N__60784\ : std_logic;
signal \N__60781\ : std_logic;
signal \N__60780\ : std_logic;
signal \N__60777\ : std_logic;
signal \N__60774\ : std_logic;
signal \N__60769\ : std_logic;
signal \N__60766\ : std_logic;
signal \N__60763\ : std_logic;
signal \N__60760\ : std_logic;
signal \N__60755\ : std_logic;
signal \N__60752\ : std_logic;
signal \N__60743\ : std_logic;
signal \N__60740\ : std_logic;
signal \N__60737\ : std_logic;
signal \N__60736\ : std_logic;
signal \N__60735\ : std_logic;
signal \N__60734\ : std_logic;
signal \N__60731\ : std_logic;
signal \N__60730\ : std_logic;
signal \N__60727\ : std_logic;
signal \N__60724\ : std_logic;
signal \N__60723\ : std_logic;
signal \N__60720\ : std_logic;
signal \N__60717\ : std_logic;
signal \N__60714\ : std_logic;
signal \N__60711\ : std_logic;
signal \N__60708\ : std_logic;
signal \N__60705\ : std_logic;
signal \N__60702\ : std_logic;
signal \N__60701\ : std_logic;
signal \N__60696\ : std_logic;
signal \N__60693\ : std_logic;
signal \N__60686\ : std_logic;
signal \N__60683\ : std_logic;
signal \N__60682\ : std_logic;
signal \N__60679\ : std_logic;
signal \N__60676\ : std_logic;
signal \N__60673\ : std_logic;
signal \N__60668\ : std_logic;
signal \N__60663\ : std_logic;
signal \N__60660\ : std_logic;
signal \N__60653\ : std_logic;
signal \N__60650\ : std_logic;
signal \N__60647\ : std_logic;
signal \N__60644\ : std_logic;
signal \N__60641\ : std_logic;
signal \N__60638\ : std_logic;
signal \N__60635\ : std_logic;
signal \N__60632\ : std_logic;
signal \N__60629\ : std_logic;
signal \N__60628\ : std_logic;
signal \N__60627\ : std_logic;
signal \N__60626\ : std_logic;
signal \N__60625\ : std_logic;
signal \N__60624\ : std_logic;
signal \N__60621\ : std_logic;
signal \N__60618\ : std_logic;
signal \N__60617\ : std_logic;
signal \N__60616\ : std_logic;
signal \N__60613\ : std_logic;
signal \N__60610\ : std_logic;
signal \N__60609\ : std_logic;
signal \N__60606\ : std_logic;
signal \N__60603\ : std_logic;
signal \N__60602\ : std_logic;
signal \N__60599\ : std_logic;
signal \N__60598\ : std_logic;
signal \N__60595\ : std_logic;
signal \N__60594\ : std_logic;
signal \N__60593\ : std_logic;
signal \N__60590\ : std_logic;
signal \N__60589\ : std_logic;
signal \N__60586\ : std_logic;
signal \N__60585\ : std_logic;
signal \N__60580\ : std_logic;
signal \N__60579\ : std_logic;
signal \N__60576\ : std_logic;
signal \N__60575\ : std_logic;
signal \N__60574\ : std_logic;
signal \N__60573\ : std_logic;
signal \N__60572\ : std_logic;
signal \N__60569\ : std_logic;
signal \N__60568\ : std_logic;
signal \N__60567\ : std_logic;
signal \N__60566\ : std_logic;
signal \N__60563\ : std_logic;
signal \N__60560\ : std_logic;
signal \N__60557\ : std_logic;
signal \N__60554\ : std_logic;
signal \N__60551\ : std_logic;
signal \N__60546\ : std_logic;
signal \N__60545\ : std_logic;
signal \N__60544\ : std_logic;
signal \N__60543\ : std_logic;
signal \N__60542\ : std_logic;
signal \N__60541\ : std_logic;
signal \N__60540\ : std_logic;
signal \N__60539\ : std_logic;
signal \N__60536\ : std_logic;
signal \N__60533\ : std_logic;
signal \N__60530\ : std_logic;
signal \N__60527\ : std_logic;
signal \N__60524\ : std_logic;
signal \N__60521\ : std_logic;
signal \N__60518\ : std_logic;
signal \N__60513\ : std_logic;
signal \N__60508\ : std_logic;
signal \N__60505\ : std_logic;
signal \N__60500\ : std_logic;
signal \N__60497\ : std_logic;
signal \N__60492\ : std_logic;
signal \N__60485\ : std_logic;
signal \N__60482\ : std_logic;
signal \N__60471\ : std_logic;
signal \N__60466\ : std_logic;
signal \N__60461\ : std_logic;
signal \N__60454\ : std_logic;
signal \N__60451\ : std_logic;
signal \N__60448\ : std_logic;
signal \N__60445\ : std_logic;
signal \N__60438\ : std_logic;
signal \N__60433\ : std_logic;
signal \N__60430\ : std_logic;
signal \N__60427\ : std_logic;
signal \N__60418\ : std_logic;
signal \N__60415\ : std_logic;
signal \N__60412\ : std_logic;
signal \N__60407\ : std_logic;
signal \N__60402\ : std_logic;
signal \N__60397\ : std_logic;
signal \N__60386\ : std_logic;
signal \N__60383\ : std_logic;
signal \N__60380\ : std_logic;
signal \N__60377\ : std_logic;
signal \N__60374\ : std_logic;
signal \N__60371\ : std_logic;
signal \N__60368\ : std_logic;
signal \N__60365\ : std_logic;
signal \N__60362\ : std_logic;
signal \N__60359\ : std_logic;
signal \N__60358\ : std_logic;
signal \N__60355\ : std_logic;
signal \N__60352\ : std_logic;
signal \N__60347\ : std_logic;
signal \N__60344\ : std_logic;
signal \N__60341\ : std_logic;
signal \N__60338\ : std_logic;
signal \N__60335\ : std_logic;
signal \N__60332\ : std_logic;
signal \N__60329\ : std_logic;
signal \N__60326\ : std_logic;
signal \N__60323\ : std_logic;
signal \N__60320\ : std_logic;
signal \N__60319\ : std_logic;
signal \N__60316\ : std_logic;
signal \N__60313\ : std_logic;
signal \N__60308\ : std_logic;
signal \N__60305\ : std_logic;
signal \N__60302\ : std_logic;
signal \N__60299\ : std_logic;
signal \N__60296\ : std_logic;
signal \N__60293\ : std_logic;
signal \N__60290\ : std_logic;
signal \N__60287\ : std_logic;
signal \N__60284\ : std_logic;
signal \N__60281\ : std_logic;
signal \N__60280\ : std_logic;
signal \N__60277\ : std_logic;
signal \N__60274\ : std_logic;
signal \N__60269\ : std_logic;
signal \N__60266\ : std_logic;
signal \N__60265\ : std_logic;
signal \N__60264\ : std_logic;
signal \N__60263\ : std_logic;
signal \N__60262\ : std_logic;
signal \N__60261\ : std_logic;
signal \N__60260\ : std_logic;
signal \N__60257\ : std_logic;
signal \N__60254\ : std_logic;
signal \N__60251\ : std_logic;
signal \N__60248\ : std_logic;
signal \N__60247\ : std_logic;
signal \N__60246\ : std_logic;
signal \N__60245\ : std_logic;
signal \N__60242\ : std_logic;
signal \N__60241\ : std_logic;
signal \N__60238\ : std_logic;
signal \N__60237\ : std_logic;
signal \N__60236\ : std_logic;
signal \N__60233\ : std_logic;
signal \N__60228\ : std_logic;
signal \N__60227\ : std_logic;
signal \N__60224\ : std_logic;
signal \N__60221\ : std_logic;
signal \N__60220\ : std_logic;
signal \N__60219\ : std_logic;
signal \N__60218\ : std_logic;
signal \N__60215\ : std_logic;
signal \N__60214\ : std_logic;
signal \N__60213\ : std_logic;
signal \N__60210\ : std_logic;
signal \N__60209\ : std_logic;
signal \N__60208\ : std_logic;
signal \N__60207\ : std_logic;
signal \N__60206\ : std_logic;
signal \N__60205\ : std_logic;
signal \N__60202\ : std_logic;
signal \N__60199\ : std_logic;
signal \N__60198\ : std_logic;
signal \N__60197\ : std_logic;
signal \N__60196\ : std_logic;
signal \N__60193\ : std_logic;
signal \N__60192\ : std_logic;
signal \N__60191\ : std_logic;
signal \N__60190\ : std_logic;
signal \N__60189\ : std_logic;
signal \N__60188\ : std_logic;
signal \N__60187\ : std_logic;
signal \N__60184\ : std_logic;
signal \N__60181\ : std_logic;
signal \N__60178\ : std_logic;
signal \N__60173\ : std_logic;
signal \N__60170\ : std_logic;
signal \N__60165\ : std_logic;
signal \N__60162\ : std_logic;
signal \N__60159\ : std_logic;
signal \N__60158\ : std_logic;
signal \N__60157\ : std_logic;
signal \N__60152\ : std_logic;
signal \N__60147\ : std_logic;
signal \N__60144\ : std_logic;
signal \N__60139\ : std_logic;
signal \N__60134\ : std_logic;
signal \N__60133\ : std_logic;
signal \N__60130\ : std_logic;
signal \N__60127\ : std_logic;
signal \N__60124\ : std_logic;
signal \N__60119\ : std_logic;
signal \N__60118\ : std_logic;
signal \N__60109\ : std_logic;
signal \N__60102\ : std_logic;
signal \N__60101\ : std_logic;
signal \N__60100\ : std_logic;
signal \N__60099\ : std_logic;
signal \N__60096\ : std_logic;
signal \N__60093\ : std_logic;
signal \N__60090\ : std_logic;
signal \N__60087\ : std_logic;
signal \N__60084\ : std_logic;
signal \N__60079\ : std_logic;
signal \N__60074\ : std_logic;
signal \N__60069\ : std_logic;
signal \N__60066\ : std_logic;
signal \N__60057\ : std_logic;
signal \N__60052\ : std_logic;
signal \N__60045\ : std_logic;
signal \N__60042\ : std_logic;
signal \N__60037\ : std_logic;
signal \N__60030\ : std_logic;
signal \N__60027\ : std_logic;
signal \N__60024\ : std_logic;
signal \N__60017\ : std_logic;
signal \N__60010\ : std_logic;
signal \N__60007\ : std_logic;
signal \N__60004\ : std_logic;
signal \N__59999\ : std_logic;
signal \N__59992\ : std_logic;
signal \N__59989\ : std_logic;
signal \N__59986\ : std_logic;
signal \N__59983\ : std_logic;
signal \N__59980\ : std_logic;
signal \N__59975\ : std_logic;
signal \N__59970\ : std_logic;
signal \N__59957\ : std_logic;
signal \N__59954\ : std_logic;
signal \N__59951\ : std_logic;
signal \N__59948\ : std_logic;
signal \N__59945\ : std_logic;
signal \N__59942\ : std_logic;
signal \N__59939\ : std_logic;
signal \N__59936\ : std_logic;
signal \N__59933\ : std_logic;
signal \N__59930\ : std_logic;
signal \N__59929\ : std_logic;
signal \N__59926\ : std_logic;
signal \N__59923\ : std_logic;
signal \N__59920\ : std_logic;
signal \N__59915\ : std_logic;
signal \N__59912\ : std_logic;
signal \N__59911\ : std_logic;
signal \N__59910\ : std_logic;
signal \N__59907\ : std_logic;
signal \N__59904\ : std_logic;
signal \N__59903\ : std_logic;
signal \N__59902\ : std_logic;
signal \N__59899\ : std_logic;
signal \N__59898\ : std_logic;
signal \N__59895\ : std_logic;
signal \N__59894\ : std_logic;
signal \N__59891\ : std_logic;
signal \N__59888\ : std_logic;
signal \N__59885\ : std_logic;
signal \N__59884\ : std_logic;
signal \N__59883\ : std_logic;
signal \N__59882\ : std_logic;
signal \N__59881\ : std_logic;
signal \N__59878\ : std_logic;
signal \N__59875\ : std_logic;
signal \N__59874\ : std_logic;
signal \N__59873\ : std_logic;
signal \N__59870\ : std_logic;
signal \N__59867\ : std_logic;
signal \N__59866\ : std_logic;
signal \N__59865\ : std_logic;
signal \N__59864\ : std_logic;
signal \N__59861\ : std_logic;
signal \N__59858\ : std_logic;
signal \N__59853\ : std_logic;
signal \N__59850\ : std_logic;
signal \N__59849\ : std_logic;
signal \N__59846\ : std_logic;
signal \N__59843\ : std_logic;
signal \N__59842\ : std_logic;
signal \N__59841\ : std_logic;
signal \N__59840\ : std_logic;
signal \N__59837\ : std_logic;
signal \N__59834\ : std_logic;
signal \N__59833\ : std_logic;
signal \N__59830\ : std_logic;
signal \N__59827\ : std_logic;
signal \N__59824\ : std_logic;
signal \N__59821\ : std_logic;
signal \N__59818\ : std_logic;
signal \N__59817\ : std_logic;
signal \N__59814\ : std_logic;
signal \N__59811\ : std_logic;
signal \N__59806\ : std_logic;
signal \N__59803\ : std_logic;
signal \N__59802\ : std_logic;
signal \N__59801\ : std_logic;
signal \N__59800\ : std_logic;
signal \N__59797\ : std_logic;
signal \N__59794\ : std_logic;
signal \N__59791\ : std_logic;
signal \N__59788\ : std_logic;
signal \N__59785\ : std_logic;
signal \N__59780\ : std_logic;
signal \N__59775\ : std_logic;
signal \N__59772\ : std_logic;
signal \N__59769\ : std_logic;
signal \N__59766\ : std_logic;
signal \N__59761\ : std_logic;
signal \N__59756\ : std_logic;
signal \N__59747\ : std_logic;
signal \N__59742\ : std_logic;
signal \N__59739\ : std_logic;
signal \N__59732\ : std_logic;
signal \N__59725\ : std_logic;
signal \N__59718\ : std_logic;
signal \N__59713\ : std_logic;
signal \N__59708\ : std_logic;
signal \N__59693\ : std_logic;
signal \N__59690\ : std_logic;
signal \N__59687\ : std_logic;
signal \N__59684\ : std_logic;
signal \N__59681\ : std_logic;
signal \N__59678\ : std_logic;
signal \N__59675\ : std_logic;
signal \N__59672\ : std_logic;
signal \N__59669\ : std_logic;
signal \N__59666\ : std_logic;
signal \N__59665\ : std_logic;
signal \N__59662\ : std_logic;
signal \N__59659\ : std_logic;
signal \N__59656\ : std_logic;
signal \N__59653\ : std_logic;
signal \N__59648\ : std_logic;
signal \N__59645\ : std_logic;
signal \N__59644\ : std_logic;
signal \N__59641\ : std_logic;
signal \N__59640\ : std_logic;
signal \N__59639\ : std_logic;
signal \N__59638\ : std_logic;
signal \N__59637\ : std_logic;
signal \N__59634\ : std_logic;
signal \N__59629\ : std_logic;
signal \N__59626\ : std_logic;
signal \N__59625\ : std_logic;
signal \N__59624\ : std_logic;
signal \N__59621\ : std_logic;
signal \N__59620\ : std_logic;
signal \N__59619\ : std_logic;
signal \N__59618\ : std_logic;
signal \N__59615\ : std_logic;
signal \N__59612\ : std_logic;
signal \N__59609\ : std_logic;
signal \N__59606\ : std_logic;
signal \N__59603\ : std_logic;
signal \N__59602\ : std_logic;
signal \N__59601\ : std_logic;
signal \N__59600\ : std_logic;
signal \N__59599\ : std_logic;
signal \N__59596\ : std_logic;
signal \N__59595\ : std_logic;
signal \N__59592\ : std_logic;
signal \N__59589\ : std_logic;
signal \N__59588\ : std_logic;
signal \N__59587\ : std_logic;
signal \N__59586\ : std_logic;
signal \N__59585\ : std_logic;
signal \N__59584\ : std_logic;
signal \N__59583\ : std_logic;
signal \N__59582\ : std_logic;
signal \N__59577\ : std_logic;
signal \N__59574\ : std_logic;
signal \N__59567\ : std_logic;
signal \N__59564\ : std_logic;
signal \N__59557\ : std_logic;
signal \N__59554\ : std_logic;
signal \N__59551\ : std_logic;
signal \N__59550\ : std_logic;
signal \N__59549\ : std_logic;
signal \N__59546\ : std_logic;
signal \N__59541\ : std_logic;
signal \N__59540\ : std_logic;
signal \N__59537\ : std_logic;
signal \N__59534\ : std_logic;
signal \N__59531\ : std_logic;
signal \N__59528\ : std_logic;
signal \N__59521\ : std_logic;
signal \N__59518\ : std_logic;
signal \N__59515\ : std_logic;
signal \N__59512\ : std_logic;
signal \N__59507\ : std_logic;
signal \N__59504\ : std_logic;
signal \N__59503\ : std_logic;
signal \N__59500\ : std_logic;
signal \N__59497\ : std_logic;
signal \N__59494\ : std_logic;
signal \N__59491\ : std_logic;
signal \N__59488\ : std_logic;
signal \N__59487\ : std_logic;
signal \N__59486\ : std_logic;
signal \N__59485\ : std_logic;
signal \N__59484\ : std_logic;
signal \N__59483\ : std_logic;
signal \N__59480\ : std_logic;
signal \N__59479\ : std_logic;
signal \N__59478\ : std_logic;
signal \N__59477\ : std_logic;
signal \N__59476\ : std_logic;
signal \N__59473\ : std_logic;
signal \N__59470\ : std_logic;
signal \N__59463\ : std_logic;
signal \N__59454\ : std_logic;
signal \N__59451\ : std_logic;
signal \N__59448\ : std_logic;
signal \N__59439\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59431\ : std_logic;
signal \N__59424\ : std_logic;
signal \N__59413\ : std_logic;
signal \N__59406\ : std_logic;
signal \N__59403\ : std_logic;
signal \N__59384\ : std_logic;
signal \N__59381\ : std_logic;
signal \N__59378\ : std_logic;
signal \N__59375\ : std_logic;
signal \N__59372\ : std_logic;
signal \N__59369\ : std_logic;
signal \N__59366\ : std_logic;
signal \N__59363\ : std_logic;
signal \N__59360\ : std_logic;
signal \N__59357\ : std_logic;
signal \N__59354\ : std_logic;
signal \N__59353\ : std_logic;
signal \N__59350\ : std_logic;
signal \N__59347\ : std_logic;
signal \N__59342\ : std_logic;
signal \N__59339\ : std_logic;
signal \N__59338\ : std_logic;
signal \N__59335\ : std_logic;
signal \N__59332\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59328\ : std_logic;
signal \N__59325\ : std_logic;
signal \N__59322\ : std_logic;
signal \N__59319\ : std_logic;
signal \N__59316\ : std_logic;
signal \N__59313\ : std_logic;
signal \N__59306\ : std_logic;
signal \N__59305\ : std_logic;
signal \N__59302\ : std_logic;
signal \N__59299\ : std_logic;
signal \N__59298\ : std_logic;
signal \N__59297\ : std_logic;
signal \N__59296\ : std_logic;
signal \N__59295\ : std_logic;
signal \N__59292\ : std_logic;
signal \N__59291\ : std_logic;
signal \N__59290\ : std_logic;
signal \N__59289\ : std_logic;
signal \N__59288\ : std_logic;
signal \N__59287\ : std_logic;
signal \N__59286\ : std_logic;
signal \N__59283\ : std_logic;
signal \N__59282\ : std_logic;
signal \N__59281\ : std_logic;
signal \N__59276\ : std_logic;
signal \N__59271\ : std_logic;
signal \N__59268\ : std_logic;
signal \N__59267\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59263\ : std_logic;
signal \N__59262\ : std_logic;
signal \N__59259\ : std_logic;
signal \N__59250\ : std_logic;
signal \N__59249\ : std_logic;
signal \N__59248\ : std_logic;
signal \N__59245\ : std_logic;
signal \N__59240\ : std_logic;
signal \N__59235\ : std_logic;
signal \N__59232\ : std_logic;
signal \N__59229\ : std_logic;
signal \N__59226\ : std_logic;
signal \N__59223\ : std_logic;
signal \N__59220\ : std_logic;
signal \N__59215\ : std_logic;
signal \N__59212\ : std_logic;
signal \N__59209\ : std_logic;
signal \N__59202\ : std_logic;
signal \N__59195\ : std_logic;
signal \N__59188\ : std_logic;
signal \N__59177\ : std_logic;
signal \N__59176\ : std_logic;
signal \N__59173\ : std_logic;
signal \N__59170\ : std_logic;
signal \N__59169\ : std_logic;
signal \N__59166\ : std_logic;
signal \N__59163\ : std_logic;
signal \N__59160\ : std_logic;
signal \N__59159\ : std_logic;
signal \N__59158\ : std_logic;
signal \N__59151\ : std_logic;
signal \N__59146\ : std_logic;
signal \N__59145\ : std_logic;
signal \N__59144\ : std_logic;
signal \N__59143\ : std_logic;
signal \N__59142\ : std_logic;
signal \N__59141\ : std_logic;
signal \N__59140\ : std_logic;
signal \N__59139\ : std_logic;
signal \N__59138\ : std_logic;
signal \N__59137\ : std_logic;
signal \N__59136\ : std_logic;
signal \N__59133\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59125\ : std_logic;
signal \N__59124\ : std_logic;
signal \N__59121\ : std_logic;
signal \N__59120\ : std_logic;
signal \N__59117\ : std_logic;
signal \N__59114\ : std_logic;
signal \N__59111\ : std_logic;
signal \N__59108\ : std_logic;
signal \N__59107\ : std_logic;
signal \N__59106\ : std_logic;
signal \N__59103\ : std_logic;
signal \N__59102\ : std_logic;
signal \N__59101\ : std_logic;
signal \N__59100\ : std_logic;
signal \N__59095\ : std_logic;
signal \N__59088\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59082\ : std_logic;
signal \N__59079\ : std_logic;
signal \N__59076\ : std_logic;
signal \N__59073\ : std_logic;
signal \N__59070\ : std_logic;
signal \N__59067\ : std_logic;
signal \N__59066\ : std_logic;
signal \N__59059\ : std_logic;
signal \N__59056\ : std_logic;
signal \N__59051\ : std_logic;
signal \N__59050\ : std_logic;
signal \N__59049\ : std_logic;
signal \N__59048\ : std_logic;
signal \N__59045\ : std_logic;
signal \N__59044\ : std_logic;
signal \N__59043\ : std_logic;
signal \N__59042\ : std_logic;
signal \N__59037\ : std_logic;
signal \N__59034\ : std_logic;
signal \N__59031\ : std_logic;
signal \N__59024\ : std_logic;
signal \N__59021\ : std_logic;
signal \N__59018\ : std_logic;
signal \N__59013\ : std_logic;
signal \N__59010\ : std_logic;
signal \N__59009\ : std_logic;
signal \N__59006\ : std_logic;
signal \N__59005\ : std_logic;
signal \N__59002\ : std_logic;
signal \N__59001\ : std_logic;
signal \N__58998\ : std_logic;
signal \N__58995\ : std_logic;
signal \N__58988\ : std_logic;
signal \N__58987\ : std_logic;
signal \N__58984\ : std_logic;
signal \N__58981\ : std_logic;
signal \N__58976\ : std_logic;
signal \N__58971\ : std_logic;
signal \N__58968\ : std_logic;
signal \N__58965\ : std_logic;
signal \N__58958\ : std_logic;
signal \N__58951\ : std_logic;
signal \N__58946\ : std_logic;
signal \N__58943\ : std_logic;
signal \N__58940\ : std_logic;
signal \N__58933\ : std_logic;
signal \N__58930\ : std_logic;
signal \N__58927\ : std_logic;
signal \N__58920\ : std_logic;
signal \N__58915\ : std_logic;
signal \N__58910\ : std_logic;
signal \N__58907\ : std_logic;
signal \N__58904\ : std_logic;
signal \N__58899\ : std_logic;
signal \N__58894\ : std_logic;
signal \N__58889\ : std_logic;
signal \N__58888\ : std_logic;
signal \N__58887\ : std_logic;
signal \N__58886\ : std_logic;
signal \N__58885\ : std_logic;
signal \N__58884\ : std_logic;
signal \N__58881\ : std_logic;
signal \N__58878\ : std_logic;
signal \N__58877\ : std_logic;
signal \N__58874\ : std_logic;
signal \N__58871\ : std_logic;
signal \N__58868\ : std_logic;
signal \N__58865\ : std_logic;
signal \N__58864\ : std_logic;
signal \N__58861\ : std_logic;
signal \N__58858\ : std_logic;
signal \N__58855\ : std_logic;
signal \N__58850\ : std_logic;
signal \N__58845\ : std_logic;
signal \N__58842\ : std_logic;
signal \N__58839\ : std_logic;
signal \N__58836\ : std_logic;
signal \N__58831\ : std_logic;
signal \N__58828\ : std_logic;
signal \N__58817\ : std_logic;
signal \N__58816\ : std_logic;
signal \N__58813\ : std_logic;
signal \N__58812\ : std_logic;
signal \N__58809\ : std_logic;
signal \N__58808\ : std_logic;
signal \N__58805\ : std_logic;
signal \N__58802\ : std_logic;
signal \N__58801\ : std_logic;
signal \N__58800\ : std_logic;
signal \N__58799\ : std_logic;
signal \N__58796\ : std_logic;
signal \N__58793\ : std_logic;
signal \N__58790\ : std_logic;
signal \N__58787\ : std_logic;
signal \N__58784\ : std_logic;
signal \N__58781\ : std_logic;
signal \N__58778\ : std_logic;
signal \N__58773\ : std_logic;
signal \N__58768\ : std_logic;
signal \N__58757\ : std_logic;
signal \N__58756\ : std_logic;
signal \N__58753\ : std_logic;
signal \N__58752\ : std_logic;
signal \N__58749\ : std_logic;
signal \N__58746\ : std_logic;
signal \N__58745\ : std_logic;
signal \N__58742\ : std_logic;
signal \N__58741\ : std_logic;
signal \N__58740\ : std_logic;
signal \N__58739\ : std_logic;
signal \N__58736\ : std_logic;
signal \N__58733\ : std_logic;
signal \N__58730\ : std_logic;
signal \N__58727\ : std_logic;
signal \N__58724\ : std_logic;
signal \N__58721\ : std_logic;
signal \N__58718\ : std_logic;
signal \N__58717\ : std_logic;
signal \N__58714\ : std_logic;
signal \N__58709\ : std_logic;
signal \N__58706\ : std_logic;
signal \N__58699\ : std_logic;
signal \N__58696\ : std_logic;
signal \N__58691\ : std_logic;
signal \N__58684\ : std_logic;
signal \N__58679\ : std_logic;
signal \N__58678\ : std_logic;
signal \N__58677\ : std_logic;
signal \N__58676\ : std_logic;
signal \N__58673\ : std_logic;
signal \N__58670\ : std_logic;
signal \N__58667\ : std_logic;
signal \N__58666\ : std_logic;
signal \N__58665\ : std_logic;
signal \N__58664\ : std_logic;
signal \N__58663\ : std_logic;
signal \N__58660\ : std_logic;
signal \N__58657\ : std_logic;
signal \N__58654\ : std_logic;
signal \N__58651\ : std_logic;
signal \N__58648\ : std_logic;
signal \N__58645\ : std_logic;
signal \N__58642\ : std_logic;
signal \N__58639\ : std_logic;
signal \N__58636\ : std_logic;
signal \N__58633\ : std_logic;
signal \N__58630\ : std_logic;
signal \N__58627\ : std_logic;
signal \N__58610\ : std_logic;
signal \N__58607\ : std_logic;
signal \N__58606\ : std_logic;
signal \N__58603\ : std_logic;
signal \N__58602\ : std_logic;
signal \N__58599\ : std_logic;
signal \N__58596\ : std_logic;
signal \N__58593\ : std_logic;
signal \N__58590\ : std_logic;
signal \N__58585\ : std_logic;
signal \N__58582\ : std_logic;
signal \N__58579\ : std_logic;
signal \N__58576\ : std_logic;
signal \N__58573\ : std_logic;
signal \N__58570\ : std_logic;
signal \N__58565\ : std_logic;
signal \N__58564\ : std_logic;
signal \N__58563\ : std_logic;
signal \N__58562\ : std_logic;
signal \N__58559\ : std_logic;
signal \N__58556\ : std_logic;
signal \N__58553\ : std_logic;
signal \N__58552\ : std_logic;
signal \N__58551\ : std_logic;
signal \N__58548\ : std_logic;
signal \N__58547\ : std_logic;
signal \N__58544\ : std_logic;
signal \N__58541\ : std_logic;
signal \N__58538\ : std_logic;
signal \N__58535\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58533\ : std_logic;
signal \N__58530\ : std_logic;
signal \N__58527\ : std_logic;
signal \N__58526\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58524\ : std_logic;
signal \N__58521\ : std_logic;
signal \N__58516\ : std_logic;
signal \N__58511\ : std_logic;
signal \N__58510\ : std_logic;
signal \N__58505\ : std_logic;
signal \N__58502\ : std_logic;
signal \N__58499\ : std_logic;
signal \N__58498\ : std_logic;
signal \N__58497\ : std_logic;
signal \N__58496\ : std_logic;
signal \N__58495\ : std_logic;
signal \N__58494\ : std_logic;
signal \N__58491\ : std_logic;
signal \N__58488\ : std_logic;
signal \N__58485\ : std_logic;
signal \N__58482\ : std_logic;
signal \N__58479\ : std_logic;
signal \N__58476\ : std_logic;
signal \N__58473\ : std_logic;
signal \N__58470\ : std_logic;
signal \N__58465\ : std_logic;
signal \N__58462\ : std_logic;
signal \N__58457\ : std_logic;
signal \N__58456\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58449\ : std_logic;
signal \N__58444\ : std_logic;
signal \N__58439\ : std_logic;
signal \N__58434\ : std_logic;
signal \N__58431\ : std_logic;
signal \N__58428\ : std_logic;
signal \N__58423\ : std_logic;
signal \N__58420\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58414\ : std_logic;
signal \N__58409\ : std_logic;
signal \N__58406\ : std_logic;
signal \N__58403\ : std_logic;
signal \N__58396\ : std_logic;
signal \N__58393\ : std_logic;
signal \N__58390\ : std_logic;
signal \N__58373\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58371\ : std_logic;
signal \N__58370\ : std_logic;
signal \N__58367\ : std_logic;
signal \N__58366\ : std_logic;
signal \N__58365\ : std_logic;
signal \N__58362\ : std_logic;
signal \N__58359\ : std_logic;
signal \N__58356\ : std_logic;
signal \N__58353\ : std_logic;
signal \N__58350\ : std_logic;
signal \N__58347\ : std_logic;
signal \N__58344\ : std_logic;
signal \N__58343\ : std_logic;
signal \N__58340\ : std_logic;
signal \N__58337\ : std_logic;
signal \N__58330\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58324\ : std_logic;
signal \N__58321\ : std_logic;
signal \N__58318\ : std_logic;
signal \N__58315\ : std_logic;
signal \N__58312\ : std_logic;
signal \N__58301\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58299\ : std_logic;
signal \N__58296\ : std_logic;
signal \N__58295\ : std_logic;
signal \N__58294\ : std_logic;
signal \N__58291\ : std_logic;
signal \N__58288\ : std_logic;
signal \N__58285\ : std_logic;
signal \N__58284\ : std_logic;
signal \N__58283\ : std_logic;
signal \N__58280\ : std_logic;
signal \N__58277\ : std_logic;
signal \N__58274\ : std_logic;
signal \N__58271\ : std_logic;
signal \N__58268\ : std_logic;
signal \N__58265\ : std_logic;
signal \N__58262\ : std_logic;
signal \N__58255\ : std_logic;
signal \N__58250\ : std_logic;
signal \N__58241\ : std_logic;
signal \N__58238\ : std_logic;
signal \N__58235\ : std_logic;
signal \N__58234\ : std_logic;
signal \N__58231\ : std_logic;
signal \N__58228\ : std_logic;
signal \N__58227\ : std_logic;
signal \N__58222\ : std_logic;
signal \N__58219\ : std_logic;
signal \N__58216\ : std_logic;
signal \N__58213\ : std_logic;
signal \N__58210\ : std_logic;
signal \N__58207\ : std_logic;
signal \N__58202\ : std_logic;
signal \N__58199\ : std_logic;
signal \N__58196\ : std_logic;
signal \N__58195\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58191\ : std_logic;
signal \N__58190\ : std_logic;
signal \N__58189\ : std_logic;
signal \N__58188\ : std_logic;
signal \N__58185\ : std_logic;
signal \N__58184\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58178\ : std_logic;
signal \N__58175\ : std_logic;
signal \N__58172\ : std_logic;
signal \N__58169\ : std_logic;
signal \N__58166\ : std_logic;
signal \N__58165\ : std_logic;
signal \N__58162\ : std_logic;
signal \N__58159\ : std_logic;
signal \N__58150\ : std_logic;
signal \N__58147\ : std_logic;
signal \N__58144\ : std_logic;
signal \N__58139\ : std_logic;
signal \N__58134\ : std_logic;
signal \N__58127\ : std_logic;
signal \N__58126\ : std_logic;
signal \N__58123\ : std_logic;
signal \N__58120\ : std_logic;
signal \N__58119\ : std_logic;
signal \N__58118\ : std_logic;
signal \N__58115\ : std_logic;
signal \N__58112\ : std_logic;
signal \N__58111\ : std_logic;
signal \N__58110\ : std_logic;
signal \N__58109\ : std_logic;
signal \N__58108\ : std_logic;
signal \N__58105\ : std_logic;
signal \N__58102\ : std_logic;
signal \N__58099\ : std_logic;
signal \N__58096\ : std_logic;
signal \N__58093\ : std_logic;
signal \N__58090\ : std_logic;
signal \N__58087\ : std_logic;
signal \N__58084\ : std_logic;
signal \N__58081\ : std_logic;
signal \N__58076\ : std_logic;
signal \N__58073\ : std_logic;
signal \N__58058\ : std_logic;
signal \N__58057\ : std_logic;
signal \N__58056\ : std_logic;
signal \N__58053\ : std_logic;
signal \N__58052\ : std_logic;
signal \N__58051\ : std_logic;
signal \N__58050\ : std_logic;
signal \N__58049\ : std_logic;
signal \N__58046\ : std_logic;
signal \N__58043\ : std_logic;
signal \N__58040\ : std_logic;
signal \N__58037\ : std_logic;
signal \N__58034\ : std_logic;
signal \N__58031\ : std_logic;
signal \N__58028\ : std_logic;
signal \N__58025\ : std_logic;
signal \N__58022\ : std_logic;
signal \N__58019\ : std_logic;
signal \N__58004\ : std_logic;
signal \N__58001\ : std_logic;
signal \N__57998\ : std_logic;
signal \N__57997\ : std_logic;
signal \N__57994\ : std_logic;
signal \N__57991\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57985\ : std_logic;
signal \N__57982\ : std_logic;
signal \N__57981\ : std_logic;
signal \N__57978\ : std_logic;
signal \N__57975\ : std_logic;
signal \N__57972\ : std_logic;
signal \N__57969\ : std_logic;
signal \N__57964\ : std_logic;
signal \N__57961\ : std_logic;
signal \N__57958\ : std_logic;
signal \N__57955\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57947\ : std_logic;
signal \N__57946\ : std_logic;
signal \N__57943\ : std_logic;
signal \N__57940\ : std_logic;
signal \N__57935\ : std_logic;
signal \N__57934\ : std_logic;
signal \N__57931\ : std_logic;
signal \N__57928\ : std_logic;
signal \N__57925\ : std_logic;
signal \N__57922\ : std_logic;
signal \N__57917\ : std_logic;
signal \N__57914\ : std_logic;
signal \N__57911\ : std_logic;
signal \N__57908\ : std_logic;
signal \N__57905\ : std_logic;
signal \N__57902\ : std_logic;
signal \N__57899\ : std_logic;
signal \N__57896\ : std_logic;
signal \N__57893\ : std_logic;
signal \N__57892\ : std_logic;
signal \N__57891\ : std_logic;
signal \N__57888\ : std_logic;
signal \N__57885\ : std_logic;
signal \N__57882\ : std_logic;
signal \N__57877\ : std_logic;
signal \N__57872\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57866\ : std_logic;
signal \N__57863\ : std_logic;
signal \N__57860\ : std_logic;
signal \N__57859\ : std_logic;
signal \N__57856\ : std_logic;
signal \N__57853\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57843\ : std_logic;
signal \N__57840\ : std_logic;
signal \N__57835\ : std_logic;
signal \N__57830\ : std_logic;
signal \N__57827\ : std_logic;
signal \N__57824\ : std_logic;
signal \N__57821\ : std_logic;
signal \N__57820\ : std_logic;
signal \N__57819\ : std_logic;
signal \N__57816\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57810\ : std_logic;
signal \N__57809\ : std_logic;
signal \N__57808\ : std_logic;
signal \N__57805\ : std_logic;
signal \N__57802\ : std_logic;
signal \N__57801\ : std_logic;
signal \N__57798\ : std_logic;
signal \N__57793\ : std_logic;
signal \N__57792\ : std_logic;
signal \N__57791\ : std_logic;
signal \N__57788\ : std_logic;
signal \N__57785\ : std_logic;
signal \N__57782\ : std_logic;
signal \N__57777\ : std_logic;
signal \N__57774\ : std_logic;
signal \N__57771\ : std_logic;
signal \N__57768\ : std_logic;
signal \N__57765\ : std_logic;
signal \N__57762\ : std_logic;
signal \N__57761\ : std_logic;
signal \N__57758\ : std_logic;
signal \N__57755\ : std_logic;
signal \N__57752\ : std_logic;
signal \N__57751\ : std_logic;
signal \N__57748\ : std_logic;
signal \N__57743\ : std_logic;
signal \N__57740\ : std_logic;
signal \N__57737\ : std_logic;
signal \N__57732\ : std_logic;
signal \N__57729\ : std_logic;
signal \N__57728\ : std_logic;
signal \N__57725\ : std_logic;
signal \N__57722\ : std_logic;
signal \N__57715\ : std_logic;
signal \N__57712\ : std_logic;
signal \N__57709\ : std_logic;
signal \N__57706\ : std_logic;
signal \N__57703\ : std_logic;
signal \N__57700\ : std_logic;
signal \N__57697\ : std_logic;
signal \N__57686\ : std_logic;
signal \N__57685\ : std_logic;
signal \N__57682\ : std_logic;
signal \N__57679\ : std_logic;
signal \N__57676\ : std_logic;
signal \N__57675\ : std_logic;
signal \N__57672\ : std_logic;
signal \N__57669\ : std_logic;
signal \N__57666\ : std_logic;
signal \N__57661\ : std_logic;
signal \N__57658\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57652\ : std_logic;
signal \N__57649\ : std_logic;
signal \N__57646\ : std_logic;
signal \N__57643\ : std_logic;
signal \N__57638\ : std_logic;
signal \N__57635\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57631\ : std_logic;
signal \N__57628\ : std_logic;
signal \N__57625\ : std_logic;
signal \N__57622\ : std_logic;
signal \N__57621\ : std_logic;
signal \N__57616\ : std_logic;
signal \N__57613\ : std_logic;
signal \N__57610\ : std_logic;
signal \N__57607\ : std_logic;
signal \N__57604\ : std_logic;
signal \N__57601\ : std_logic;
signal \N__57598\ : std_logic;
signal \N__57593\ : std_logic;
signal \N__57590\ : std_logic;
signal \N__57587\ : std_logic;
signal \N__57586\ : std_logic;
signal \N__57583\ : std_logic;
signal \N__57582\ : std_logic;
signal \N__57579\ : std_logic;
signal \N__57576\ : std_logic;
signal \N__57573\ : std_logic;
signal \N__57570\ : std_logic;
signal \N__57567\ : std_logic;
signal \N__57564\ : std_logic;
signal \N__57561\ : std_logic;
signal \N__57558\ : std_logic;
signal \N__57555\ : std_logic;
signal \N__57552\ : std_logic;
signal \N__57549\ : std_logic;
signal \N__57546\ : std_logic;
signal \N__57543\ : std_logic;
signal \N__57540\ : std_logic;
signal \N__57537\ : std_logic;
signal \N__57534\ : std_logic;
signal \N__57527\ : std_logic;
signal \N__57524\ : std_logic;
signal \N__57523\ : std_logic;
signal \N__57518\ : std_logic;
signal \N__57515\ : std_logic;
signal \N__57514\ : std_logic;
signal \N__57511\ : std_logic;
signal \N__57508\ : std_logic;
signal \N__57503\ : std_logic;
signal \N__57500\ : std_logic;
signal \N__57497\ : std_logic;
signal \N__57494\ : std_logic;
signal \N__57491\ : std_logic;
signal \N__57488\ : std_logic;
signal \N__57485\ : std_logic;
signal \N__57482\ : std_logic;
signal \N__57479\ : std_logic;
signal \N__57476\ : std_logic;
signal \N__57473\ : std_logic;
signal \N__57470\ : std_logic;
signal \N__57467\ : std_logic;
signal \N__57464\ : std_logic;
signal \N__57461\ : std_logic;
signal \N__57458\ : std_logic;
signal \N__57455\ : std_logic;
signal \N__57454\ : std_logic;
signal \N__57451\ : std_logic;
signal \N__57448\ : std_logic;
signal \N__57445\ : std_logic;
signal \N__57442\ : std_logic;
signal \N__57439\ : std_logic;
signal \N__57436\ : std_logic;
signal \N__57433\ : std_logic;
signal \N__57430\ : std_logic;
signal \N__57427\ : std_logic;
signal \N__57422\ : std_logic;
signal \N__57421\ : std_logic;
signal \N__57420\ : std_logic;
signal \N__57419\ : std_logic;
signal \N__57416\ : std_logic;
signal \N__57413\ : std_logic;
signal \N__57412\ : std_logic;
signal \N__57407\ : std_logic;
signal \N__57406\ : std_logic;
signal \N__57405\ : std_logic;
signal \N__57400\ : std_logic;
signal \N__57397\ : std_logic;
signal \N__57396\ : std_logic;
signal \N__57393\ : std_logic;
signal \N__57390\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57388\ : std_logic;
signal \N__57385\ : std_logic;
signal \N__57384\ : std_logic;
signal \N__57383\ : std_logic;
signal \N__57382\ : std_logic;
signal \N__57379\ : std_logic;
signal \N__57378\ : std_logic;
signal \N__57373\ : std_logic;
signal \N__57372\ : std_logic;
signal \N__57371\ : std_logic;
signal \N__57368\ : std_logic;
signal \N__57365\ : std_logic;
signal \N__57360\ : std_logic;
signal \N__57355\ : std_logic;
signal \N__57352\ : std_logic;
signal \N__57351\ : std_logic;
signal \N__57350\ : std_logic;
signal \N__57349\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57343\ : std_logic;
signal \N__57340\ : std_logic;
signal \N__57337\ : std_logic;
signal \N__57332\ : std_logic;
signal \N__57329\ : std_logic;
signal \N__57322\ : std_logic;
signal \N__57321\ : std_logic;
signal \N__57316\ : std_logic;
signal \N__57311\ : std_logic;
signal \N__57300\ : std_logic;
signal \N__57295\ : std_logic;
signal \N__57292\ : std_logic;
signal \N__57285\ : std_logic;
signal \N__57282\ : std_logic;
signal \N__57279\ : std_logic;
signal \N__57276\ : std_logic;
signal \N__57273\ : std_logic;
signal \N__57270\ : std_logic;
signal \N__57267\ : std_logic;
signal \N__57264\ : std_logic;
signal \N__57261\ : std_logic;
signal \N__57258\ : std_logic;
signal \N__57255\ : std_logic;
signal \N__57248\ : std_logic;
signal \N__57245\ : std_logic;
signal \N__57242\ : std_logic;
signal \N__57239\ : std_logic;
signal \N__57238\ : std_logic;
signal \N__57235\ : std_logic;
signal \N__57232\ : std_logic;
signal \N__57231\ : std_logic;
signal \N__57228\ : std_logic;
signal \N__57227\ : std_logic;
signal \N__57224\ : std_logic;
signal \N__57221\ : std_logic;
signal \N__57218\ : std_logic;
signal \N__57215\ : std_logic;
signal \N__57212\ : std_logic;
signal \N__57209\ : std_logic;
signal \N__57204\ : std_logic;
signal \N__57199\ : std_logic;
signal \N__57196\ : std_logic;
signal \N__57193\ : std_logic;
signal \N__57190\ : std_logic;
signal \N__57185\ : std_logic;
signal \N__57182\ : std_logic;
signal \N__57179\ : std_logic;
signal \N__57176\ : std_logic;
signal \N__57173\ : std_logic;
signal \N__57170\ : std_logic;
signal \N__57167\ : std_logic;
signal \N__57166\ : std_logic;
signal \N__57163\ : std_logic;
signal \N__57160\ : std_logic;
signal \N__57157\ : std_logic;
signal \N__57154\ : std_logic;
signal \N__57151\ : std_logic;
signal \N__57148\ : std_logic;
signal \N__57145\ : std_logic;
signal \N__57142\ : std_logic;
signal \N__57137\ : std_logic;
signal \N__57134\ : std_logic;
signal \N__57131\ : std_logic;
signal \N__57128\ : std_logic;
signal \N__57125\ : std_logic;
signal \N__57122\ : std_logic;
signal \N__57121\ : std_logic;
signal \N__57118\ : std_logic;
signal \N__57113\ : std_logic;
signal \N__57110\ : std_logic;
signal \N__57109\ : std_logic;
signal \N__57104\ : std_logic;
signal \N__57101\ : std_logic;
signal \N__57098\ : std_logic;
signal \N__57095\ : std_logic;
signal \N__57094\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57088\ : std_logic;
signal \N__57085\ : std_logic;
signal \N__57082\ : std_logic;
signal \N__57077\ : std_logic;
signal \N__57074\ : std_logic;
signal \N__57073\ : std_logic;
signal \N__57068\ : std_logic;
signal \N__57065\ : std_logic;
signal \N__57062\ : std_logic;
signal \N__57059\ : std_logic;
signal \N__57056\ : std_logic;
signal \N__57053\ : std_logic;
signal \N__57050\ : std_logic;
signal \N__57047\ : std_logic;
signal \N__57046\ : std_logic;
signal \N__57043\ : std_logic;
signal \N__57040\ : std_logic;
signal \N__57039\ : std_logic;
signal \N__57034\ : std_logic;
signal \N__57033\ : std_logic;
signal \N__57032\ : std_logic;
signal \N__57031\ : std_logic;
signal \N__57030\ : std_logic;
signal \N__57029\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57025\ : std_logic;
signal \N__57024\ : std_logic;
signal \N__57021\ : std_logic;
signal \N__57016\ : std_logic;
signal \N__57015\ : std_logic;
signal \N__57012\ : std_logic;
signal \N__57009\ : std_logic;
signal \N__57006\ : std_logic;
signal \N__57003\ : std_logic;
signal \N__57000\ : std_logic;
signal \N__56997\ : std_logic;
signal \N__56994\ : std_logic;
signal \N__56991\ : std_logic;
signal \N__56988\ : std_logic;
signal \N__56987\ : std_logic;
signal \N__56984\ : std_logic;
signal \N__56977\ : std_logic;
signal \N__56974\ : std_logic;
signal \N__56971\ : std_logic;
signal \N__56966\ : std_logic;
signal \N__56963\ : std_logic;
signal \N__56960\ : std_logic;
signal \N__56955\ : std_logic;
signal \N__56942\ : std_logic;
signal \N__56939\ : std_logic;
signal \N__56936\ : std_logic;
signal \N__56933\ : std_logic;
signal \N__56930\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56928\ : std_logic;
signal \N__56925\ : std_logic;
signal \N__56920\ : std_logic;
signal \N__56917\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56911\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56909\ : std_logic;
signal \N__56906\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56901\ : std_logic;
signal \N__56900\ : std_logic;
signal \N__56895\ : std_logic;
signal \N__56892\ : std_logic;
signal \N__56889\ : std_logic;
signal \N__56886\ : std_logic;
signal \N__56883\ : std_logic;
signal \N__56880\ : std_logic;
signal \N__56877\ : std_logic;
signal \N__56870\ : std_logic;
signal \N__56865\ : std_logic;
signal \N__56862\ : std_logic;
signal \N__56859\ : std_logic;
signal \N__56852\ : std_logic;
signal \N__56849\ : std_logic;
signal \N__56846\ : std_logic;
signal \N__56843\ : std_logic;
signal \N__56840\ : std_logic;
signal \N__56839\ : std_logic;
signal \N__56836\ : std_logic;
signal \N__56833\ : std_logic;
signal \N__56830\ : std_logic;
signal \N__56829\ : std_logic;
signal \N__56828\ : std_logic;
signal \N__56825\ : std_logic;
signal \N__56824\ : std_logic;
signal \N__56823\ : std_logic;
signal \N__56820\ : std_logic;
signal \N__56815\ : std_logic;
signal \N__56812\ : std_logic;
signal \N__56809\ : std_logic;
signal \N__56806\ : std_logic;
signal \N__56805\ : std_logic;
signal \N__56804\ : std_logic;
signal \N__56799\ : std_logic;
signal \N__56796\ : std_logic;
signal \N__56793\ : std_logic;
signal \N__56788\ : std_logic;
signal \N__56787\ : std_logic;
signal \N__56784\ : std_logic;
signal \N__56781\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56773\ : std_logic;
signal \N__56768\ : std_logic;
signal \N__56759\ : std_logic;
signal \N__56756\ : std_logic;
signal \N__56753\ : std_logic;
signal \N__56750\ : std_logic;
signal \N__56749\ : std_logic;
signal \N__56748\ : std_logic;
signal \N__56745\ : std_logic;
signal \N__56742\ : std_logic;
signal \N__56741\ : std_logic;
signal \N__56738\ : std_logic;
signal \N__56737\ : std_logic;
signal \N__56734\ : std_logic;
signal \N__56731\ : std_logic;
signal \N__56728\ : std_logic;
signal \N__56723\ : std_logic;
signal \N__56720\ : std_logic;
signal \N__56719\ : std_logic;
signal \N__56718\ : std_logic;
signal \N__56713\ : std_logic;
signal \N__56710\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56702\ : std_logic;
signal \N__56699\ : std_logic;
signal \N__56696\ : std_logic;
signal \N__56693\ : std_logic;
signal \N__56688\ : std_logic;
signal \N__56685\ : std_logic;
signal \N__56678\ : std_logic;
signal \N__56675\ : std_logic;
signal \N__56672\ : std_logic;
signal \N__56669\ : std_logic;
signal \N__56666\ : std_logic;
signal \N__56663\ : std_logic;
signal \N__56660\ : std_logic;
signal \N__56657\ : std_logic;
signal \N__56656\ : std_logic;
signal \N__56651\ : std_logic;
signal \N__56648\ : std_logic;
signal \N__56647\ : std_logic;
signal \N__56644\ : std_logic;
signal \N__56641\ : std_logic;
signal \N__56638\ : std_logic;
signal \N__56635\ : std_logic;
signal \N__56632\ : std_logic;
signal \N__56627\ : std_logic;
signal \N__56624\ : std_logic;
signal \N__56623\ : std_logic;
signal \N__56622\ : std_logic;
signal \N__56621\ : std_logic;
signal \N__56618\ : std_logic;
signal \N__56615\ : std_logic;
signal \N__56610\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56604\ : std_logic;
signal \N__56603\ : std_logic;
signal \N__56600\ : std_logic;
signal \N__56595\ : std_logic;
signal \N__56592\ : std_logic;
signal \N__56589\ : std_logic;
signal \N__56586\ : std_logic;
signal \N__56583\ : std_logic;
signal \N__56580\ : std_logic;
signal \N__56577\ : std_logic;
signal \N__56574\ : std_logic;
signal \N__56573\ : std_logic;
signal \N__56570\ : std_logic;
signal \N__56567\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56561\ : std_logic;
signal \N__56558\ : std_logic;
signal \N__56555\ : std_logic;
signal \N__56552\ : std_logic;
signal \N__56543\ : std_logic;
signal \N__56542\ : std_logic;
signal \N__56539\ : std_logic;
signal \N__56536\ : std_logic;
signal \N__56533\ : std_logic;
signal \N__56532\ : std_logic;
signal \N__56529\ : std_logic;
signal \N__56526\ : std_logic;
signal \N__56523\ : std_logic;
signal \N__56520\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56514\ : std_logic;
signal \N__56511\ : std_logic;
signal \N__56506\ : std_logic;
signal \N__56503\ : std_logic;
signal \N__56500\ : std_logic;
signal \N__56495\ : std_logic;
signal \N__56492\ : std_logic;
signal \N__56491\ : std_logic;
signal \N__56490\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56482\ : std_logic;
signal \N__56479\ : std_logic;
signal \N__56474\ : std_logic;
signal \N__56473\ : std_logic;
signal \N__56472\ : std_logic;
signal \N__56469\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56465\ : std_logic;
signal \N__56462\ : std_logic;
signal \N__56459\ : std_logic;
signal \N__56456\ : std_logic;
signal \N__56453\ : std_logic;
signal \N__56450\ : std_logic;
signal \N__56445\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56439\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56431\ : std_logic;
signal \N__56426\ : std_logic;
signal \N__56423\ : std_logic;
signal \N__56420\ : std_logic;
signal \N__56417\ : std_logic;
signal \N__56416\ : std_logic;
signal \N__56415\ : std_logic;
signal \N__56414\ : std_logic;
signal \N__56413\ : std_logic;
signal \N__56410\ : std_logic;
signal \N__56407\ : std_logic;
signal \N__56402\ : std_logic;
signal \N__56401\ : std_logic;
signal \N__56398\ : std_logic;
signal \N__56395\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56391\ : std_logic;
signal \N__56388\ : std_logic;
signal \N__56385\ : std_logic;
signal \N__56382\ : std_logic;
signal \N__56379\ : std_logic;
signal \N__56378\ : std_logic;
signal \N__56377\ : std_logic;
signal \N__56374\ : std_logic;
signal \N__56371\ : std_logic;
signal \N__56366\ : std_logic;
signal \N__56361\ : std_logic;
signal \N__56360\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56358\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56352\ : std_logic;
signal \N__56347\ : std_logic;
signal \N__56346\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56342\ : std_logic;
signal \N__56339\ : std_logic;
signal \N__56336\ : std_logic;
signal \N__56329\ : std_logic;
signal \N__56328\ : std_logic;
signal \N__56327\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56321\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56313\ : std_logic;
signal \N__56306\ : std_logic;
signal \N__56303\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56285\ : std_logic;
signal \N__56282\ : std_logic;
signal \N__56279\ : std_logic;
signal \N__56276\ : std_logic;
signal \N__56273\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56268\ : std_logic;
signal \N__56267\ : std_logic;
signal \N__56266\ : std_logic;
signal \N__56263\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56259\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56241\ : std_logic;
signal \N__56240\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56229\ : std_logic;
signal \N__56228\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56223\ : std_logic;
signal \N__56218\ : std_logic;
signal \N__56213\ : std_logic;
signal \N__56206\ : std_logic;
signal \N__56203\ : std_logic;
signal \N__56202\ : std_logic;
signal \N__56201\ : std_logic;
signal \N__56200\ : std_logic;
signal \N__56197\ : std_logic;
signal \N__56196\ : std_logic;
signal \N__56193\ : std_logic;
signal \N__56188\ : std_logic;
signal \N__56185\ : std_logic;
signal \N__56182\ : std_logic;
signal \N__56179\ : std_logic;
signal \N__56168\ : std_logic;
signal \N__56165\ : std_logic;
signal \N__56150\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56144\ : std_logic;
signal \N__56141\ : std_logic;
signal \N__56138\ : std_logic;
signal \N__56135\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56131\ : std_logic;
signal \N__56130\ : std_logic;
signal \N__56127\ : std_logic;
signal \N__56124\ : std_logic;
signal \N__56121\ : std_logic;
signal \N__56120\ : std_logic;
signal \N__56117\ : std_logic;
signal \N__56116\ : std_logic;
signal \N__56115\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56109\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56100\ : std_logic;
signal \N__56097\ : std_logic;
signal \N__56096\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56090\ : std_logic;
signal \N__56087\ : std_logic;
signal \N__56086\ : std_logic;
signal \N__56083\ : std_logic;
signal \N__56082\ : std_logic;
signal \N__56079\ : std_logic;
signal \N__56078\ : std_logic;
signal \N__56077\ : std_logic;
signal \N__56076\ : std_logic;
signal \N__56073\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56069\ : std_logic;
signal \N__56068\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56060\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56054\ : std_logic;
signal \N__56051\ : std_logic;
signal \N__56048\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56032\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56022\ : std_logic;
signal \N__56003\ : std_logic;
signal \N__56000\ : std_logic;
signal \N__55997\ : std_logic;
signal \N__55994\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55992\ : std_logic;
signal \N__55991\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55989\ : std_logic;
signal \N__55986\ : std_logic;
signal \N__55985\ : std_logic;
signal \N__55984\ : std_logic;
signal \N__55979\ : std_logic;
signal \N__55976\ : std_logic;
signal \N__55973\ : std_logic;
signal \N__55970\ : std_logic;
signal \N__55967\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55958\ : std_logic;
signal \N__55957\ : std_logic;
signal \N__55954\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55949\ : std_logic;
signal \N__55946\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55938\ : std_logic;
signal \N__55931\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55925\ : std_logic;
signal \N__55922\ : std_logic;
signal \N__55919\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55913\ : std_logic;
signal \N__55904\ : std_logic;
signal \N__55901\ : std_logic;
signal \N__55898\ : std_logic;
signal \N__55893\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55887\ : std_logic;
signal \N__55886\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55879\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55862\ : std_logic;
signal \N__55859\ : std_logic;
signal \N__55854\ : std_logic;
signal \N__55851\ : std_logic;
signal \N__55848\ : std_logic;
signal \N__55835\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55829\ : std_logic;
signal \N__55826\ : std_logic;
signal \N__55823\ : std_logic;
signal \N__55822\ : std_logic;
signal \N__55821\ : std_logic;
signal \N__55818\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55816\ : std_logic;
signal \N__55813\ : std_logic;
signal \N__55812\ : std_logic;
signal \N__55811\ : std_logic;
signal \N__55808\ : std_logic;
signal \N__55805\ : std_logic;
signal \N__55802\ : std_logic;
signal \N__55801\ : std_logic;
signal \N__55800\ : std_logic;
signal \N__55799\ : std_logic;
signal \N__55796\ : std_logic;
signal \N__55793\ : std_logic;
signal \N__55788\ : std_logic;
signal \N__55783\ : std_logic;
signal \N__55780\ : std_logic;
signal \N__55777\ : std_logic;
signal \N__55772\ : std_logic;
signal \N__55769\ : std_logic;
signal \N__55768\ : std_logic;
signal \N__55767\ : std_logic;
signal \N__55764\ : std_logic;
signal \N__55761\ : std_logic;
signal \N__55752\ : std_logic;
signal \N__55749\ : std_logic;
signal \N__55746\ : std_logic;
signal \N__55743\ : std_logic;
signal \N__55740\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55734\ : std_logic;
signal \N__55727\ : std_logic;
signal \N__55726\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55721\ : std_logic;
signal \N__55716\ : std_logic;
signal \N__55713\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55691\ : std_logic;
signal \N__55688\ : std_logic;
signal \N__55687\ : std_logic;
signal \N__55686\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55682\ : std_logic;
signal \N__55681\ : std_logic;
signal \N__55678\ : std_logic;
signal \N__55675\ : std_logic;
signal \N__55674\ : std_logic;
signal \N__55671\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55665\ : std_logic;
signal \N__55662\ : std_logic;
signal \N__55661\ : std_logic;
signal \N__55660\ : std_logic;
signal \N__55657\ : std_logic;
signal \N__55654\ : std_logic;
signal \N__55651\ : std_logic;
signal \N__55648\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55644\ : std_logic;
signal \N__55641\ : std_logic;
signal \N__55638\ : std_logic;
signal \N__55635\ : std_logic;
signal \N__55628\ : std_logic;
signal \N__55625\ : std_logic;
signal \N__55622\ : std_logic;
signal \N__55619\ : std_logic;
signal \N__55612\ : std_logic;
signal \N__55609\ : std_logic;
signal \N__55598\ : std_logic;
signal \N__55595\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55589\ : std_logic;
signal \N__55586\ : std_logic;
signal \N__55585\ : std_logic;
signal \N__55582\ : std_logic;
signal \N__55579\ : std_logic;
signal \N__55578\ : std_logic;
signal \N__55577\ : std_logic;
signal \N__55576\ : std_logic;
signal \N__55573\ : std_logic;
signal \N__55570\ : std_logic;
signal \N__55565\ : std_logic;
signal \N__55562\ : std_logic;
signal \N__55559\ : std_logic;
signal \N__55558\ : std_logic;
signal \N__55555\ : std_logic;
signal \N__55550\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55547\ : std_logic;
signal \N__55546\ : std_logic;
signal \N__55543\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55535\ : std_logic;
signal \N__55526\ : std_logic;
signal \N__55517\ : std_logic;
signal \N__55514\ : std_logic;
signal \N__55511\ : std_logic;
signal \N__55508\ : std_logic;
signal \N__55505\ : std_logic;
signal \N__55502\ : std_logic;
signal \N__55499\ : std_logic;
signal \N__55496\ : std_logic;
signal \N__55493\ : std_logic;
signal \N__55490\ : std_logic;
signal \N__55487\ : std_logic;
signal \N__55484\ : std_logic;
signal \N__55481\ : std_logic;
signal \N__55478\ : std_logic;
signal \N__55475\ : std_logic;
signal \N__55474\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55472\ : std_logic;
signal \N__55471\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55467\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55462\ : std_logic;
signal \N__55457\ : std_logic;
signal \N__55456\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55453\ : std_logic;
signal \N__55452\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55436\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55424\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55422\ : std_logic;
signal \N__55421\ : std_logic;
signal \N__55418\ : std_logic;
signal \N__55413\ : std_logic;
signal \N__55408\ : std_logic;
signal \N__55405\ : std_logic;
signal \N__55400\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55393\ : std_logic;
signal \N__55386\ : std_logic;
signal \N__55381\ : std_logic;
signal \N__55376\ : std_logic;
signal \N__55373\ : std_logic;
signal \N__55370\ : std_logic;
signal \N__55365\ : std_logic;
signal \N__55360\ : std_logic;
signal \N__55357\ : std_logic;
signal \N__55354\ : std_logic;
signal \N__55351\ : std_logic;
signal \N__55346\ : std_logic;
signal \N__55343\ : std_logic;
signal \N__55334\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55330\ : std_logic;
signal \N__55327\ : std_logic;
signal \N__55324\ : std_logic;
signal \N__55321\ : std_logic;
signal \N__55318\ : std_logic;
signal \N__55315\ : std_logic;
signal \N__55312\ : std_logic;
signal \N__55309\ : std_logic;
signal \N__55306\ : std_logic;
signal \N__55301\ : std_logic;
signal \N__55298\ : std_logic;
signal \N__55295\ : std_logic;
signal \N__55294\ : std_logic;
signal \N__55291\ : std_logic;
signal \N__55288\ : std_logic;
signal \N__55283\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55277\ : std_logic;
signal \N__55274\ : std_logic;
signal \N__55271\ : std_logic;
signal \N__55268\ : std_logic;
signal \N__55265\ : std_logic;
signal \N__55262\ : std_logic;
signal \N__55259\ : std_logic;
signal \N__55256\ : std_logic;
signal \N__55253\ : std_logic;
signal \N__55250\ : std_logic;
signal \N__55247\ : std_logic;
signal \N__55244\ : std_logic;
signal \N__55241\ : std_logic;
signal \N__55238\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55232\ : std_logic;
signal \N__55229\ : std_logic;
signal \N__55226\ : std_logic;
signal \N__55223\ : std_logic;
signal \N__55222\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55215\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55205\ : std_logic;
signal \N__55202\ : std_logic;
signal \N__55199\ : std_logic;
signal \N__55196\ : std_logic;
signal \N__55193\ : std_logic;
signal \N__55190\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55184\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55177\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55168\ : std_logic;
signal \N__55167\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55159\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55155\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55146\ : std_logic;
signal \N__55139\ : std_logic;
signal \N__55138\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55134\ : std_logic;
signal \N__55131\ : std_logic;
signal \N__55128\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55122\ : std_logic;
signal \N__55121\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55119\ : std_logic;
signal \N__55118\ : std_logic;
signal \N__55115\ : std_logic;
signal \N__55112\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55104\ : std_logic;
signal \N__55099\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55078\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55074\ : std_logic;
signal \N__55071\ : std_logic;
signal \N__55068\ : std_logic;
signal \N__55065\ : std_logic;
signal \N__55064\ : std_logic;
signal \N__55059\ : std_logic;
signal \N__55058\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55056\ : std_logic;
signal \N__55055\ : std_logic;
signal \N__55054\ : std_logic;
signal \N__55053\ : std_logic;
signal \N__55050\ : std_logic;
signal \N__55047\ : std_logic;
signal \N__55044\ : std_logic;
signal \N__55041\ : std_logic;
signal \N__55036\ : std_logic;
signal \N__55033\ : std_logic;
signal \N__55028\ : std_logic;
signal \N__55013\ : std_logic;
signal \N__55010\ : std_logic;
signal \N__55007\ : std_logic;
signal \N__55004\ : std_logic;
signal \N__55001\ : std_logic;
signal \N__54998\ : std_logic;
signal \N__54995\ : std_logic;
signal \N__54992\ : std_logic;
signal \N__54989\ : std_logic;
signal \N__54986\ : std_logic;
signal \N__54983\ : std_logic;
signal \N__54980\ : std_logic;
signal \N__54977\ : std_logic;
signal \N__54974\ : std_logic;
signal \N__54971\ : std_logic;
signal \N__54968\ : std_logic;
signal \N__54965\ : std_logic;
signal \N__54962\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54956\ : std_logic;
signal \N__54953\ : std_logic;
signal \N__54950\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54944\ : std_logic;
signal \N__54941\ : std_logic;
signal \N__54938\ : std_logic;
signal \N__54935\ : std_logic;
signal \N__54932\ : std_logic;
signal \N__54929\ : std_logic;
signal \N__54926\ : std_logic;
signal \N__54923\ : std_logic;
signal \N__54922\ : std_logic;
signal \N__54919\ : std_logic;
signal \N__54916\ : std_logic;
signal \N__54913\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54905\ : std_logic;
signal \N__54902\ : std_logic;
signal \N__54901\ : std_logic;
signal \N__54898\ : std_logic;
signal \N__54895\ : std_logic;
signal \N__54890\ : std_logic;
signal \N__54889\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54878\ : std_logic;
signal \N__54875\ : std_logic;
signal \N__54872\ : std_logic;
signal \N__54869\ : std_logic;
signal \N__54866\ : std_logic;
signal \N__54863\ : std_logic;
signal \N__54860\ : std_logic;
signal \N__54857\ : std_logic;
signal \N__54854\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54848\ : std_logic;
signal \N__54845\ : std_logic;
signal \N__54842\ : std_logic;
signal \N__54839\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54833\ : std_logic;
signal \N__54830\ : std_logic;
signal \N__54827\ : std_logic;
signal \N__54824\ : std_logic;
signal \N__54821\ : std_logic;
signal \N__54818\ : std_logic;
signal \N__54815\ : std_logic;
signal \N__54814\ : std_logic;
signal \N__54811\ : std_logic;
signal \N__54808\ : std_logic;
signal \N__54803\ : std_logic;
signal \N__54802\ : std_logic;
signal \N__54799\ : std_logic;
signal \N__54796\ : std_logic;
signal \N__54791\ : std_logic;
signal \N__54788\ : std_logic;
signal \N__54785\ : std_logic;
signal \N__54782\ : std_logic;
signal \N__54779\ : std_logic;
signal \N__54776\ : std_logic;
signal \N__54773\ : std_logic;
signal \N__54770\ : std_logic;
signal \N__54767\ : std_logic;
signal \N__54766\ : std_logic;
signal \N__54763\ : std_logic;
signal \N__54760\ : std_logic;
signal \N__54757\ : std_logic;
signal \N__54752\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54746\ : std_logic;
signal \N__54741\ : std_logic;
signal \N__54738\ : std_logic;
signal \N__54735\ : std_logic;
signal \N__54732\ : std_logic;
signal \N__54729\ : std_logic;
signal \N__54726\ : std_logic;
signal \N__54723\ : std_logic;
signal \N__54720\ : std_logic;
signal \N__54719\ : std_logic;
signal \N__54716\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54708\ : std_logic;
signal \N__54707\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54699\ : std_logic;
signal \N__54696\ : std_logic;
signal \N__54689\ : std_logic;
signal \N__54688\ : std_logic;
signal \N__54687\ : std_logic;
signal \N__54686\ : std_logic;
signal \N__54685\ : std_logic;
signal \N__54682\ : std_logic;
signal \N__54681\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54679\ : std_logic;
signal \N__54678\ : std_logic;
signal \N__54677\ : std_logic;
signal \N__54674\ : std_logic;
signal \N__54671\ : std_logic;
signal \N__54670\ : std_logic;
signal \N__54669\ : std_logic;
signal \N__54668\ : std_logic;
signal \N__54665\ : std_logic;
signal \N__54662\ : std_logic;
signal \N__54661\ : std_logic;
signal \N__54660\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54658\ : std_logic;
signal \N__54657\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54655\ : std_logic;
signal \N__54654\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54652\ : std_logic;
signal \N__54651\ : std_logic;
signal \N__54648\ : std_logic;
signal \N__54641\ : std_logic;
signal \N__54636\ : std_logic;
signal \N__54635\ : std_logic;
signal \N__54634\ : std_logic;
signal \N__54633\ : std_logic;
signal \N__54632\ : std_logic;
signal \N__54627\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54615\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54602\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54587\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54584\ : std_logic;
signal \N__54583\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54579\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54575\ : std_logic;
signal \N__54574\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54572\ : std_logic;
signal \N__54571\ : std_logic;
signal \N__54570\ : std_logic;
signal \N__54569\ : std_logic;
signal \N__54568\ : std_logic;
signal \N__54563\ : std_logic;
signal \N__54560\ : std_logic;
signal \N__54553\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54545\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54543\ : std_logic;
signal \N__54542\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54540\ : std_logic;
signal \N__54539\ : std_logic;
signal \N__54536\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54514\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54506\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54494\ : std_logic;
signal \N__54491\ : std_logic;
signal \N__54486\ : std_logic;
signal \N__54477\ : std_logic;
signal \N__54474\ : std_logic;
signal \N__54469\ : std_logic;
signal \N__54466\ : std_logic;
signal \N__54461\ : std_logic;
signal \N__54458\ : std_logic;
signal \N__54453\ : std_logic;
signal \N__54446\ : std_logic;
signal \N__54435\ : std_logic;
signal \N__54426\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54398\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54392\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54386\ : std_logic;
signal \N__54383\ : std_logic;
signal \N__54380\ : std_logic;
signal \N__54377\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54371\ : std_logic;
signal \N__54368\ : std_logic;
signal \N__54365\ : std_logic;
signal \N__54362\ : std_logic;
signal \N__54359\ : std_logic;
signal \N__54358\ : std_logic;
signal \N__54357\ : std_logic;
signal \N__54356\ : std_logic;
signal \N__54355\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54335\ : std_logic;
signal \N__54332\ : std_logic;
signal \N__54329\ : std_logic;
signal \N__54328\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54320\ : std_logic;
signal \N__54317\ : std_logic;
signal \N__54314\ : std_logic;
signal \N__54311\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54305\ : std_logic;
signal \N__54304\ : std_logic;
signal \N__54303\ : std_logic;
signal \N__54300\ : std_logic;
signal \N__54299\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54296\ : std_logic;
signal \N__54295\ : std_logic;
signal \N__54294\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54292\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54286\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54284\ : std_logic;
signal \N__54281\ : std_logic;
signal \N__54276\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54266\ : std_logic;
signal \N__54261\ : std_logic;
signal \N__54258\ : std_logic;
signal \N__54255\ : std_logic;
signal \N__54250\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54244\ : std_logic;
signal \N__54237\ : std_logic;
signal \N__54236\ : std_logic;
signal \N__54235\ : std_logic;
signal \N__54234\ : std_logic;
signal \N__54231\ : std_logic;
signal \N__54228\ : std_logic;
signal \N__54225\ : std_logic;
signal \N__54222\ : std_logic;
signal \N__54217\ : std_logic;
signal \N__54212\ : std_logic;
signal \N__54209\ : std_logic;
signal \N__54194\ : std_logic;
signal \N__54191\ : std_logic;
signal \N__54188\ : std_logic;
signal \N__54187\ : std_logic;
signal \N__54186\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54175\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54169\ : std_logic;
signal \N__54166\ : std_logic;
signal \N__54161\ : std_logic;
signal \N__54158\ : std_logic;
signal \N__54155\ : std_logic;
signal \N__54152\ : std_logic;
signal \N__54149\ : std_logic;
signal \N__54146\ : std_logic;
signal \N__54143\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54141\ : std_logic;
signal \N__54140\ : std_logic;
signal \N__54139\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54135\ : std_logic;
signal \N__54134\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54129\ : std_logic;
signal \N__54128\ : std_logic;
signal \N__54125\ : std_logic;
signal \N__54122\ : std_logic;
signal \N__54119\ : std_logic;
signal \N__54118\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54114\ : std_logic;
signal \N__54113\ : std_logic;
signal \N__54112\ : std_logic;
signal \N__54111\ : std_logic;
signal \N__54110\ : std_logic;
signal \N__54107\ : std_logic;
signal \N__54104\ : std_logic;
signal \N__54101\ : std_logic;
signal \N__54098\ : std_logic;
signal \N__54093\ : std_logic;
signal \N__54090\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54082\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54074\ : std_logic;
signal \N__54069\ : std_logic;
signal \N__54066\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54062\ : std_logic;
signal \N__54061\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54059\ : std_logic;
signal \N__54056\ : std_logic;
signal \N__54047\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54041\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54029\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54019\ : std_logic;
signal \N__54012\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__53990\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53984\ : std_logic;
signal \N__53981\ : std_logic;
signal \N__53978\ : std_logic;
signal \N__53975\ : std_logic;
signal \N__53972\ : std_logic;
signal \N__53969\ : std_logic;
signal \N__53968\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53966\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53964\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53962\ : std_logic;
signal \N__53961\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53953\ : std_logic;
signal \N__53952\ : std_logic;
signal \N__53951\ : std_logic;
signal \N__53946\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53942\ : std_logic;
signal \N__53941\ : std_logic;
signal \N__53940\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53938\ : std_logic;
signal \N__53937\ : std_logic;
signal \N__53936\ : std_logic;
signal \N__53931\ : std_logic;
signal \N__53924\ : std_logic;
signal \N__53919\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53910\ : std_logic;
signal \N__53909\ : std_logic;
signal \N__53904\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53890\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53888\ : std_logic;
signal \N__53887\ : std_logic;
signal \N__53882\ : std_logic;
signal \N__53879\ : std_logic;
signal \N__53876\ : std_logic;
signal \N__53873\ : std_logic;
signal \N__53870\ : std_logic;
signal \N__53867\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53861\ : std_logic;
signal \N__53860\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53837\ : std_logic;
signal \N__53828\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53820\ : std_logic;
signal \N__53817\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53796\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53774\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53768\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53762\ : std_logic;
signal \N__53759\ : std_logic;
signal \N__53758\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53749\ : std_logic;
signal \N__53744\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53738\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53732\ : std_logic;
signal \N__53729\ : std_logic;
signal \N__53726\ : std_logic;
signal \N__53723\ : std_logic;
signal \N__53720\ : std_logic;
signal \N__53719\ : std_logic;
signal \N__53718\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53714\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53706\ : std_logic;
signal \N__53705\ : std_logic;
signal \N__53704\ : std_logic;
signal \N__53701\ : std_logic;
signal \N__53698\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53677\ : std_logic;
signal \N__53674\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53668\ : std_logic;
signal \N__53667\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53663\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53661\ : std_logic;
signal \N__53658\ : std_logic;
signal \N__53653\ : std_logic;
signal \N__53650\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53642\ : std_logic;
signal \N__53639\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53627\ : std_logic;
signal \N__53624\ : std_logic;
signal \N__53621\ : std_logic;
signal \N__53618\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53611\ : std_logic;
signal \N__53608\ : std_logic;
signal \N__53605\ : std_logic;
signal \N__53602\ : std_logic;
signal \N__53599\ : std_logic;
signal \N__53596\ : std_logic;
signal \N__53593\ : std_logic;
signal \N__53588\ : std_logic;
signal \N__53585\ : std_logic;
signal \N__53584\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53580\ : std_logic;
signal \N__53575\ : std_logic;
signal \N__53574\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53572\ : std_logic;
signal \N__53571\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53567\ : std_logic;
signal \N__53564\ : std_logic;
signal \N__53561\ : std_logic;
signal \N__53558\ : std_logic;
signal \N__53555\ : std_logic;
signal \N__53550\ : std_logic;
signal \N__53545\ : std_logic;
signal \N__53534\ : std_logic;
signal \N__53531\ : std_logic;
signal \N__53530\ : std_logic;
signal \N__53527\ : std_logic;
signal \N__53524\ : std_logic;
signal \N__53521\ : std_logic;
signal \N__53518\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53514\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53508\ : std_logic;
signal \N__53505\ : std_logic;
signal \N__53502\ : std_logic;
signal \N__53499\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53480\ : std_logic;
signal \N__53479\ : std_logic;
signal \N__53478\ : std_logic;
signal \N__53477\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53471\ : std_logic;
signal \N__53468\ : std_logic;
signal \N__53467\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53463\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53455\ : std_logic;
signal \N__53450\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53434\ : std_logic;
signal \N__53431\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53429\ : std_logic;
signal \N__53426\ : std_logic;
signal \N__53425\ : std_logic;
signal \N__53422\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53407\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53402\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53400\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53389\ : std_logic;
signal \N__53384\ : std_logic;
signal \N__53381\ : std_logic;
signal \N__53376\ : std_logic;
signal \N__53363\ : std_logic;
signal \N__53360\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53354\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53348\ : std_logic;
signal \N__53345\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53336\ : std_logic;
signal \N__53333\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53323\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53317\ : std_logic;
signal \N__53314\ : std_logic;
signal \N__53309\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53305\ : std_logic;
signal \N__53304\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53301\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53299\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53297\ : std_logic;
signal \N__53296\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53294\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53292\ : std_logic;
signal \N__53291\ : std_logic;
signal \N__53290\ : std_logic;
signal \N__53289\ : std_logic;
signal \N__53288\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53267\ : std_logic;
signal \N__53264\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53249\ : std_logic;
signal \N__53246\ : std_logic;
signal \N__53245\ : std_logic;
signal \N__53242\ : std_logic;
signal \N__53239\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53234\ : std_logic;
signal \N__53233\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53231\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53216\ : std_logic;
signal \N__53209\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53205\ : std_logic;
signal \N__53204\ : std_logic;
signal \N__53201\ : std_logic;
signal \N__53198\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53178\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53174\ : std_logic;
signal \N__53171\ : std_logic;
signal \N__53166\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53162\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53158\ : std_logic;
signal \N__53155\ : std_logic;
signal \N__53152\ : std_logic;
signal \N__53147\ : std_logic;
signal \N__53146\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53138\ : std_logic;
signal \N__53133\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53122\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53112\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53106\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53094\ : std_logic;
signal \N__53089\ : std_logic;
signal \N__53086\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53072\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53045\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53039\ : std_logic;
signal \N__53036\ : std_logic;
signal \N__53033\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53027\ : std_logic;
signal \N__53024\ : std_logic;
signal \N__53021\ : std_logic;
signal \N__53018\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52994\ : std_logic;
signal \N__52991\ : std_logic;
signal \N__52988\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52974\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52968\ : std_logic;
signal \N__52965\ : std_logic;
signal \N__52958\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52950\ : std_logic;
signal \N__52947\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52937\ : std_logic;
signal \N__52936\ : std_logic;
signal \N__52935\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52932\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52913\ : std_logic;
signal \N__52910\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52902\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52878\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52870\ : std_logic;
signal \N__52867\ : std_logic;
signal \N__52866\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52856\ : std_logic;
signal \N__52853\ : std_logic;
signal \N__52850\ : std_logic;
signal \N__52847\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52839\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52825\ : std_logic;
signal \N__52822\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52808\ : std_logic;
signal \N__52807\ : std_logic;
signal \N__52806\ : std_logic;
signal \N__52805\ : std_logic;
signal \N__52802\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52798\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52792\ : std_logic;
signal \N__52789\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52787\ : std_logic;
signal \N__52786\ : std_logic;
signal \N__52783\ : std_logic;
signal \N__52780\ : std_logic;
signal \N__52777\ : std_logic;
signal \N__52772\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52766\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52744\ : std_logic;
signal \N__52741\ : std_logic;
signal \N__52738\ : std_logic;
signal \N__52735\ : std_logic;
signal \N__52732\ : std_logic;
signal \N__52729\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52720\ : std_logic;
signal \N__52717\ : std_logic;
signal \N__52714\ : std_logic;
signal \N__52709\ : std_logic;
signal \N__52706\ : std_logic;
signal \N__52705\ : std_logic;
signal \N__52702\ : std_logic;
signal \N__52699\ : std_logic;
signal \N__52696\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52688\ : std_logic;
signal \N__52685\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52680\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52666\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52657\ : std_logic;
signal \N__52654\ : std_logic;
signal \N__52645\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52637\ : std_logic;
signal \N__52636\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52627\ : std_logic;
signal \N__52624\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52612\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52597\ : std_logic;
signal \N__52592\ : std_logic;
signal \N__52589\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52572\ : std_logic;
signal \N__52565\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52538\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52528\ : std_logic;
signal \N__52527\ : std_logic;
signal \N__52524\ : std_logic;
signal \N__52521\ : std_logic;
signal \N__52518\ : std_logic;
signal \N__52515\ : std_logic;
signal \N__52510\ : std_logic;
signal \N__52507\ : std_logic;
signal \N__52504\ : std_logic;
signal \N__52499\ : std_logic;
signal \N__52496\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52412\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52389\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52366\ : std_logic;
signal \N__52363\ : std_logic;
signal \N__52358\ : std_logic;
signal \N__52357\ : std_logic;
signal \N__52354\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52341\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52329\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52315\ : std_logic;
signal \N__52312\ : std_logic;
signal \N__52307\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52298\ : std_logic;
signal \N__52295\ : std_logic;
signal \N__52292\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52270\ : std_logic;
signal \N__52267\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52252\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52242\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52196\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52178\ : std_logic;
signal \N__52175\ : std_logic;
signal \N__52166\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52138\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52129\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52123\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52117\ : std_logic;
signal \N__52114\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52097\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52080\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52067\ : std_logic;
signal \N__52064\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52053\ : std_logic;
signal \N__52052\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52049\ : std_logic;
signal \N__52046\ : std_logic;
signal \N__52043\ : std_logic;
signal \N__52040\ : std_logic;
signal \N__52037\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52011\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51989\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51981\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51968\ : std_logic;
signal \N__51967\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51961\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51952\ : std_logic;
signal \N__51949\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51941\ : std_logic;
signal \N__51938\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51933\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51930\ : std_logic;
signal \N__51929\ : std_logic;
signal \N__51926\ : std_logic;
signal \N__51923\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51911\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51898\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51883\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51872\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51862\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51848\ : std_logic;
signal \N__51845\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51839\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51806\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51799\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51788\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51780\ : std_logic;
signal \N__51779\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51777\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51757\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51692\ : std_logic;
signal \N__51689\ : std_logic;
signal \N__51686\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51680\ : std_logic;
signal \N__51677\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51635\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51632\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51611\ : std_logic;
signal \N__51608\ : std_logic;
signal \N__51605\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51584\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51580\ : std_logic;
signal \N__51577\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51565\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51554\ : std_logic;
signal \N__51551\ : std_logic;
signal \N__51548\ : std_logic;
signal \N__51545\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51529\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51512\ : std_logic;
signal \N__51509\ : std_logic;
signal \N__51506\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51461\ : std_logic;
signal \N__51458\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51385\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51350\ : std_logic;
signal \N__51347\ : std_logic;
signal \N__51344\ : std_logic;
signal \N__51341\ : std_logic;
signal \N__51338\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51334\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51304\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51292\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51263\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51253\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51214\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51173\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51155\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51149\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51125\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51121\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51107\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51098\ : std_logic;
signal \N__51095\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51083\ : std_logic;
signal \N__51080\ : std_logic;
signal \N__51077\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51068\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51064\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51053\ : std_logic;
signal \N__51050\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51035\ : std_logic;
signal \N__51032\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51023\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51017\ : std_logic;
signal \N__51014\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51008\ : std_logic;
signal \N__51005\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50996\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50987\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50959\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50947\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50935\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50918\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50890\ : std_logic;
signal \N__50887\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50863\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50843\ : std_logic;
signal \N__50842\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50838\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50827\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50738\ : std_logic;
signal \N__50735\ : std_logic;
signal \N__50732\ : std_logic;
signal \N__50729\ : std_logic;
signal \N__50726\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50720\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50690\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50684\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50639\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50630\ : std_logic;
signal \N__50627\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50591\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50569\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50474\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50441\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50383\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50222\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50190\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50133\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50102\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50029\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50021\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49969\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49622\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49601\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49595\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49584\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49006\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48083\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43214\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42665\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \INVCONTROL.addrstack_addrstack_0_0RCLKN_net\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_3RCLKN_net\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_2RCLKN_net\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_1RCLKN_net\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_0RCLKN_net\ : std_logic;
signal \GNDG0\ : std_logic;
signal \clkdivZ0Z_0\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \clkdivZ0Z_1\ : std_logic;
signal clkdiv_cry_0 : std_logic;
signal \clkdivZ0Z_2\ : std_logic;
signal clkdiv_cry_1 : std_logic;
signal \clkdivZ0Z_3\ : std_logic;
signal clkdiv_cry_2 : std_logic;
signal \clkdivZ0Z_4\ : std_logic;
signal clkdiv_cry_3 : std_logic;
signal \clkdivZ0Z_5\ : std_logic;
signal clkdiv_cry_4 : std_logic;
signal \clkdivZ0Z_6\ : std_logic;
signal clkdiv_cry_5 : std_logic;
signal \clkdivZ0Z_7\ : std_logic;
signal clkdiv_cry_6 : std_logic;
signal clkdiv_cry_7 : std_logic;
signal \clkdivZ0Z_8\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \clkdivZ0Z_9\ : std_logic;
signal clkdiv_cry_8 : std_logic;
signal \clkdivZ0Z_10\ : std_logic;
signal clkdiv_cry_9 : std_logic;
signal \clkdivZ0Z_11\ : std_logic;
signal clkdiv_cry_10 : std_logic;
signal \clkdivZ0Z_12\ : std_logic;
signal clkdiv_cry_11 : std_logic;
signal \clkdivZ0Z_13\ : std_logic;
signal clkdiv_cry_12 : std_logic;
signal \clkdivZ0Z_14\ : std_logic;
signal clkdiv_cry_13 : std_logic;
signal \clkdivZ0Z_15\ : std_logic;
signal clkdiv_cry_14 : std_logic;
signal clkdiv_cry_15 : std_logic;
signal \clkdivZ0Z_16\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \clkdivZ0Z_17\ : std_logic;
signal clkdiv_cry_16 : std_logic;
signal \clkdivZ0Z_18\ : std_logic;
signal clkdiv_cry_17 : std_logic;
signal \clkdivZ0Z_19\ : std_logic;
signal clkdiv_cry_18 : std_logic;
signal \clkdivZ0Z_20\ : std_logic;
signal clkdiv_cry_19 : std_logic;
signal \clkdivZ0Z_21\ : std_logic;
signal clkdiv_cry_20 : std_logic;
signal \clkdivZ0Z_22\ : std_logic;
signal clkdiv_cry_21 : std_logic;
signal clkdiv_cry_22 : std_logic;
signal \GPIO3_c\ : std_logic;
signal \B_OE_c_i\ : std_logic;
signal \B_OE_c\ : std_logic;
signal \gpuAddress_11\ : std_logic;
signal \INVCONTROL.gpuAddReg_11C_net\ : std_logic;
signal \gpuAddress_14\ : std_logic;
signal \INVCONTROL.gpuAddReg_14C_net\ : std_logic;
signal \gpuAddress_9\ : std_logic;
signal \INVCONTROL.gpuAddReg_9C_net\ : std_logic;
signal \N_6_0\ : std_logic;
signal \RAM_un1_WR_i\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \ALU.status_17_data_tmp_0\ : std_logic;
signal \ALU.status_17_data_tmp_1\ : std_logic;
signal \ALU.status_17_data_tmp_2\ : std_logic;
signal \ALU.status_17_data_tmp_3\ : std_logic;
signal \ALU.status_17_data_tmp_4\ : std_logic;
signal \ALU.status_17_data_tmp_5\ : std_logic;
signal \ALU.status_17_data_tmp_6\ : std_logic;
signal \ALU.status_17_data_tmp_7\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \ALU.status_17_I_45_c_RNOZ0\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \ALU.combOperand2_i_1\ : std_logic;
signal \ALU.status_18_cry_0\ : std_logic;
signal \ALU.status_18_cry_1\ : std_logic;
signal \ALU.status_18_cry_2\ : std_logic;
signal \ALU.status_18_cry_3\ : std_logic;
signal \ALU.status_18_cry_4\ : std_logic;
signal \ALU.status_17_I_27_c_RNOZ0\ : std_logic;
signal \ALU.status_18_cry_5\ : std_logic;
signal \ALU.combOperand2_i_7\ : std_logic;
signal \ALU.status_18_cry_6\ : std_logic;
signal \ALU.status_18_cry_7\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \ALU.status_18_cry_8\ : std_logic;
signal \ALU.status_18_cry_9\ : std_logic;
signal \ALU.combOperand2_i_11\ : std_logic;
signal \ALU.status_18_cry_10\ : std_logic;
signal \ALU.status_18_cry_11\ : std_logic;
signal \ALU.status_18_cry_12\ : std_logic;
signal \ALU.combOperand2_i_14\ : std_logic;
signal \ALU.status_18_cry_13\ : std_logic;
signal \ALU.combOperand2_i_15\ : std_logic;
signal \ALU.status_18_cry_14\ : std_logic;
signal \ALU.status_18_4\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \ALU.status_18_cry_10_c_RNOZ0\ : std_logic;
signal \ALU.status_18_cry_13_c_RNOZ0\ : std_logic;
signal \CONTROL.busState_1_RNIG7366Z0Z_2_cascade_\ : std_logic;
signal \CONTROL.busState_1_RNI1JVK1_0Z0Z_2\ : std_logic;
signal \gpuOut_c_5\ : std_logic;
signal \CONTROL.N_166\ : std_logic;
signal \D5_in_c\ : std_logic;
signal \CONTROL.N_166_cascade_\ : std_logic;
signal \romOut_5\ : std_logic;
signal \INVCONTROL.dout_5C_net\ : std_logic;
signal \ALU.operand2_12_cascade_\ : std_logic;
signal \ALU.N_126_cascade_\ : std_logic;
signal \ALU.c_RNI670LZ0Z_12_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_12\ : std_logic;
signal \ALU.d_RNI8FCTZ0Z_12\ : std_logic;
signal \ALU.operand2_12\ : std_logic;
signal \ALU.status_18_cry_12_c_RNOZ0\ : std_logic;
signal \ALU.log_1_3cf0_1_10\ : std_logic;
signal \ALU.log_1_3cf0_10_cascade_\ : std_logic;
signal \ALU.log_1_3cf1_10\ : std_logic;
signal \ALU.log_1_3cf1_1_10\ : std_logic;
signal \CONTROL.bus_7_a0_2_8_cascade_\ : std_logic;
signal \ALU.status_18_cry_8_c_RNOZ0\ : std_logic;
signal \DROM_ROMDATA_dintern_8ro_cascade_\ : std_logic;
signal \DROM_ROMDATA_dintern_8ro\ : std_logic;
signal bus_8 : std_logic;
signal \DROM.ROMDATA.dintern_0_0_NEW_1\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_OLDZ0Z_1\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C_net\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_NEW_0\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_OLDZ0Z_0\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net\ : std_logic;
signal \DROM_ROMDATA_dintern_12ro_cascade_\ : std_logic;
signal \INVCONTROL.aluOperation_3C_net\ : std_logic;
signal \DROM_ROMDATA_dintern_12ro\ : std_logic;
signal bus_12 : std_logic;
signal \DROM.ROMDATA.dintern_0_3_OLDZ0Z_2\ : std_logic;
signal \DROM.ROMDATA.dintern_0_3_NEW_2\ : std_logic;
signal \DROM.ROMDATA.dintern_0_3_OLDZ0Z_3\ : std_logic;
signal \DROM.ROMDATA.dintern_0_3_NEW_3\ : std_logic;
signal bus_10 : std_logic;
signal \gpuAddress_0\ : std_logic;
signal \gpuAddress_1\ : std_logic;
signal \gpuAddress_10\ : std_logic;
signal \gpuAddress_12\ : std_logic;
signal \gpuAddress_13\ : std_logic;
signal \gpuAddress_15\ : std_logic;
signal \INVCONTROL.gpuAddReg_0C_net\ : std_logic;
signal \CONTROL_romAddReg_7_2\ : std_logic;
signal \CONTROL_romAddReg_7_3\ : std_logic;
signal \INVCONTROL.dout_3C_net\ : std_logic;
signal \CONTROL_romAddReg_7_5\ : std_logic;
signal \PROM_ROMDATA_dintern_23ro_cascade_\ : std_logic;
signal \CONTROL_romAddReg_7_7\ : std_logic;
signal \CONTROL_romAddReg_7_6\ : std_logic;
signal \PROM.ROMDATA.m465_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m471_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m471_ns_cascade_\ : std_logic;
signal \controlWord_24_cascade_\ : std_logic;
signal \CONTROL_romAddReg_7_8\ : std_logic;
signal \CONTROL_romAddReg_7_4\ : std_logic;
signal \CONTROL.g0_3_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_N_10_mux_0_0_0_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_N_7_0_i\ : std_logic;
signal \CONTROL.N_6_1_cascade_\ : std_logic;
signal \CONTROL.N_4_2\ : std_logic;
signal \CONTROL.N_4_2_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_N_10_mux_0_0_0\ : std_logic;
signal \INVCONTROL.addrstackptr_6C_net\ : std_logic;
signal \CONTROL.tempCounterZ0Z_13\ : std_logic;
signal \CONTROL.tempCounterZ0Z_6\ : std_logic;
signal \INVCONTROL.tempCounter_13C_net\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \CONTROL.addrstack_1_cry_0\ : std_logic;
signal \CONTROL.addrstack_1_cry_1\ : std_logic;
signal \CONTROL.addrstack_1_cry_2\ : std_logic;
signal \CONTROL.addrstack_1_cry_3\ : std_logic;
signal \CONTROL.addrstack_1_cry_4\ : std_logic;
signal \CONTROL.addrstackptrZ0Z_6\ : std_logic;
signal \CONTROL.addrstack_1_6\ : std_logic;
signal \CONTROL.addrstack_1_cry_5\ : std_logic;
signal \CONTROL.addrstack_1_cry_6\ : std_logic;
signal \ALU.dout_3_ns_1_5_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_5_cascade_\ : std_logic;
signal \ALU.N_1138_cascade_\ : std_logic;
signal \ALU.N_1090\ : std_logic;
signal \aluOut_5_cascade_\ : std_logic;
signal \ALU.status_19_4_cascade_\ : std_logic;
signal \ALU.status_17_I_15_c_RNOZ0\ : std_logic;
signal \ALU.combOperand2_0_6\ : std_logic;
signal \ALU.combOperand2_0_6_cascade_\ : std_logic;
signal \ALU.status_19_5_cascade_\ : std_logic;
signal \ALU.combOperand2_0_4_cascade_\ : std_logic;
signal \N_181_cascade_\ : std_logic;
signal \ALU.d_RNIVKK66Z0Z_4\ : std_logic;
signal \ALU.d_RNIVKK66Z0Z_4_cascade_\ : std_logic;
signal \ALU.combOperand2_0_4\ : std_logic;
signal \ALU.status_17_I_33_c_RNOZ0\ : std_logic;
signal \N_182\ : std_logic;
signal \ALU.combOperand2_0_0_6\ : std_logic;
signal \ALU.b_RNI4VJC1Z0Z_12\ : std_logic;
signal \ALU.d_RNI4BCTZ0Z_10\ : std_logic;
signal \ALU.b_RNI0RJC1Z0Z_10_cascade_\ : std_logic;
signal \ALU.operand2_10\ : std_logic;
signal \ALU.operand2_10_cascade_\ : std_logic;
signal \ALU.status_19_9_cascade_\ : std_logic;
signal \ALU.e_RNIBHMNZ0Z_8_cascade_\ : std_logic;
signal \ALU.d_RNIIINJZ0Z_8\ : std_logic;
signal \ALU.operand2_7_ns_1_8\ : std_logic;
signal \ALU.b_RNIE6BVZ0Z_8_cascade_\ : std_logic;
signal \ALU.operand2_8\ : std_logic;
signal \busState_1_RNI05PC2_0\ : std_logic;
signal \ALU.operand2_8_cascade_\ : std_logic;
signal \ALU.status_18_cry_3_c_RNOZ0\ : std_logic;
signal \N_228_0_cascade_\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C_net\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_OLDZ0Z_3\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_NEW_3\ : std_logic;
signal \DROM_ROMDATA_dintern_3ro_cascade_\ : std_logic;
signal \DROM_ROMDATA_dintern_1ro\ : std_logic;
signal \DROM_ROMDATA_dintern_adflt_cascade_\ : std_logic;
signal \DROM.ROMDATA.dintern_adfltZ0Z_3\ : std_logic;
signal \DROM.ROMDATA.dintern_adfltZ0Z_3_cascade_\ : std_logic;
signal \DROM.ROMDATA.dintern_adflt_sxZ0\ : std_logic;
signal \dataRomAddress_13\ : std_logic;
signal \dataRomAddress_14\ : std_logic;
signal \dataRomAddress_15\ : std_logic;
signal \INVCONTROL.romAddReg_13C_net\ : std_logic;
signal \INVCONTROL.aluOperation_ne_0C_net\ : std_logic;
signal \DROM.ROMDATA.dintern_0_3_OLDZ0Z_1\ : std_logic;
signal \DROM.ROMDATA.dintern_0_3_NEW_1\ : std_logic;
signal \DROM_ROMDATA_dintern_13ro_cascade_\ : std_logic;
signal \CONTROL.bus_7_a0_2_8\ : std_logic;
signal \DROM_ROMDATA_dintern_13ro\ : std_logic;
signal bus_13 : std_logic;
signal \DROM_ROMDATA_dintern_10ro\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_NEW_1\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_OLDZ0Z_1\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_NEW_2\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_OLDZ0Z_2\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_NEW_1\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_OLDZ0Z_1\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_NEW_2\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_OLDZ0Z_2\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_NEW_3\ : std_logic;
signal \DROM.ROMDATA.dintern_0_2_OLDZ0Z_3\ : std_logic;
signal \DROM.ROMDATA.dintern_0_3_NEW_0\ : std_logic;
signal \DROM.ROMDATA.dintern_0_3_OLDZ0Z_0\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\ : std_logic;
signal \DROM_ROMDATA_dintern_6ro\ : std_logic;
signal \CONTROL.N_199_cascade_\ : std_logic;
signal \gpuOut_c_6\ : std_logic;
signal \D6_in_c\ : std_logic;
signal \CONTROL.N_167_cascade_\ : std_logic;
signal \N_183\ : std_logic;
signal \INVCONTROL.dout_6C_net\ : std_logic;
signal \CONTROL.addrstackptr_N_8_mux_1_0_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_N_6_0_1_i\ : std_logic;
signal \CONTROL.g0_3_i_2_cascade_\ : std_logic;
signal \CONTROL.N_4_0\ : std_logic;
signal \CONTROL.addrstack_1_5\ : std_logic;
signal \CONTROL.N_4_0_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_N_8_mux_1_0\ : std_logic;
signal \CONTROL.addrstackptrZ0Z_5\ : std_logic;
signal \INVCONTROL.addrstackptr_5C_net\ : std_logic;
signal \CONTROL.g0_3_iZ0Z_1\ : std_logic;
signal \CONTROL.g0_3_i_a7Z0Z_2\ : std_logic;
signal \CONTROL.g0_0_2\ : std_logic;
signal \CONTROL.addrstack_12\ : std_logic;
signal \CONTROL.addrstack_11\ : std_logic;
signal \CONTROL.addrstack_7\ : std_logic;
signal \CONTROL.addrstack_14\ : std_logic;
signal \CONTROL.tempCounterZ0Z_11\ : std_logic;
signal \CONTROL.tempCounterZ0Z_15\ : std_logic;
signal \CONTROL.tempCounterZ0Z_14\ : std_logic;
signal \INVCONTROL.tempCounter_11C_net\ : std_logic;
signal \CONTROL.addrstack_8\ : std_logic;
signal \CONTROL.addrstack_9\ : std_logic;
signal \ALU.status_17_I_9_c_RNOZ0\ : std_logic;
signal \ALU.addsub_cry_3_c_RNIGCKVJZ0Z5_cascade_\ : std_logic;
signal \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9_cascade_\ : std_logic;
signal \ALU.e_RNI26JMZ0Z_4_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_4_cascade_\ : std_logic;
signal \ALU.operand2_4\ : std_logic;
signal \ALU.c_RNI6IVQZ0Z_4\ : std_logic;
signal \ALU.dout_6_ns_1_4_cascade_\ : std_logic;
signal \ALU.aZ0Z_4\ : std_logic;
signal \ALU.dout_3_ns_1_4_cascade_\ : std_logic;
signal \ALU.N_1089_cascade_\ : std_logic;
signal \ALU.N_1137\ : std_logic;
signal \aluOut_4_cascade_\ : std_logic;
signal \ALU.d_RNIBJM75Z0Z_4\ : std_logic;
signal \ALU.status_19_8_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_6_cascade_\ : std_logic;
signal \ALU.operand2_6\ : std_logic;
signal \ALU.b_RNI9JSPZ0Z_6\ : std_logic;
signal \ALU.e_RNI6AJMZ0Z_6\ : std_logic;
signal \ALU.c_RNIAMVQZ0Z_6\ : std_logic;
signal \ALU.d_RNIDV8EZ0Z_6\ : std_logic;
signal \ALU.c_RNI230LZ0Z_10\ : std_logic;
signal \ALU.a_RNIUI741Z0Z_10_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_10\ : std_logic;
signal \ALU.dout_6_ns_1_8_cascade_\ : std_logic;
signal \ALU_N_1141_cascade_\ : std_logic;
signal \CONTROL.bus_0_sx_8_cascade_\ : std_logic;
signal \CONTROL_bus_0_8\ : std_logic;
signal \ALU.dout_3_ns_1_8_cascade_\ : std_logic;
signal \ALU.c_RNIFT2SZ0Z_8\ : std_logic;
signal \dataRomAddress_10\ : std_logic;
signal \dataRomAddress_12\ : std_logic;
signal \PROM.ROMDATA.dintern_adfltZ0Z_4_cascade_\ : std_logic;
signal \PROM.ROMDATA.dintern_12dflt_0Z0Z_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.dintern_adfltZ0Z_4\ : std_logic;
signal \dataRomAddress_11\ : std_logic;
signal \INVCONTROL.romAddReg_10C_net\ : std_logic;
signal \CONTROL.busState_1_e_1_0_cascade_\ : std_logic;
signal \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0_cascade_\ : std_logic;
signal \N_29\ : std_logic;
signal \CONTROL.N_352\ : std_logic;
signal \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0\ : std_logic;
signal \INVCONTROL.busState_1_0C_net\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_OLDZ0Z_3\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_NEW_3\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_OLDZ0Z_0\ : std_logic;
signal \DROM.ROMDATA.dintern_0_1_NEW_0\ : std_logic;
signal \DROM_ROMDATA_dintern_4ro\ : std_logic;
signal \controlWord_29\ : std_logic;
signal \controlWord_29_cascade_\ : std_logic;
signal \controlWord_28\ : std_logic;
signal \controlWord_28_cascade_\ : std_logic;
signal \INVCONTROL.ramAddReg_13C_net\ : std_logic;
signal \A12_c\ : std_logic;
signal \A13_c\ : std_logic;
signal \RAM.un1_WR_105_0Z0Z_10\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \CONTROL.programCounter_1_cry_0\ : std_logic;
signal \CONTROL.programCounter_1_cry_1\ : std_logic;
signal \CONTROL.programCounter_1_axb_3\ : std_logic;
signal \CONTROL.programCounter_1_cry_2\ : std_logic;
signal \CONTROL.programCounter_1_cry_3\ : std_logic;
signal \CONTROL.programCounter_1_cry_4\ : std_logic;
signal \CONTROL.programCounter_1_cry_5\ : std_logic;
signal \CONTROL.programCounter_1_cry_6\ : std_logic;
signal \CONTROL.programCounter_1_cry_7\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \CONTROL.programCounter_1_cry_8\ : std_logic;
signal \CONTROL.programCounter_1_cry_9\ : std_logic;
signal \CONTROL.programCounter_1_cry_10\ : std_logic;
signal \CONTROL.programCounter_1_cry_11\ : std_logic;
signal \CONTROL.programCounter_1_cry_12\ : std_logic;
signal \CONTROL.programCounter_1_cry_13\ : std_logic;
signal \CONTROL.programCounter_1_cry_14\ : std_logic;
signal \CONTROL.programCounter_1_13\ : std_logic;
signal \CONTROL.programCounter_1_reto_13\ : std_logic;
signal \CONTROL.dout_reto_13\ : std_logic;
signal \CONTROL.N_428_cascade_\ : std_logic;
signal \progRomAddress_13\ : std_logic;
signal \CONTROL.addrstack_reto_14\ : std_logic;
signal \progRomAddress_14\ : std_logic;
signal \CONTROL.addrstack_13\ : std_logic;
signal \CONTROL.addrstack_reto_13\ : std_logic;
signal \progRomAddress_10\ : std_logic;
signal \CONTROL.addrstack_reto_12\ : std_logic;
signal \progRomAddress_12\ : std_logic;
signal \CONTROL.addrstack_10\ : std_logic;
signal \CONTROL.addrstack_reto_10\ : std_logic;
signal \CONTROL.programCounter_1_reto_8\ : std_logic;
signal \N_423_cascade_\ : std_logic;
signal \CONTROL.programCounter_1_axb_8\ : std_logic;
signal \CONTROL.programCounter10\ : std_logic;
signal \CONTROL.programCounter_1_reto_9\ : std_logic;
signal \CONTROL.addrstack_reto_9\ : std_logic;
signal \CONTROL.N_424_cascade_\ : std_logic;
signal \progRomAddress_9\ : std_logic;
signal \CONTROL_addrstack_reto_8\ : std_logic;
signal \N_423\ : std_logic;
signal \progRomAddress_9_cascade_\ : std_logic;
signal \PROM.ROMDATA.dintern_adfltZ0Z_3\ : std_logic;
signal \CONTROL.tempCounterZ0Z_10\ : std_logic;
signal \CONTROL.programCounter_1_9\ : std_logic;
signal \CONTROL.tempCounterZ0Z_9\ : std_logic;
signal \INVCONTROL.tempCounter_10C_net\ : std_logic;
signal \INVCONTROL.addrstackptr_0C_net\ : std_logic;
signal \ALU.rshift_3_ns_1_2\ : std_logic;
signal \ALU.status_17_I_1_c_RNOZ0\ : std_logic;
signal \ALU.N_834_cascade_\ : std_logic;
signal \busState_1_RNIDU0U1_2\ : std_logic;
signal \ALU.status_19_2_cascade_\ : std_logic;
signal \romOut_4\ : std_logic;
signal \CONTROL.busState_1_RNI7U266Z0Z_2\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \ALU.mult_3_c3\ : std_logic;
signal \ALU.d_RNITK2D51Z0Z_2\ : std_logic;
signal \ALU.mult_3_c4\ : std_logic;
signal \ALU.d_RNIJBM6GZ0Z_3\ : std_logic;
signal \ALU.d_RNIKG0L11Z0Z_2\ : std_logic;
signal \ALU.mult_3_c5\ : std_logic;
signal \ALU.d_RNI9DAEHZ0Z_3\ : std_logic;
signal \ALU.d_RNI07V431Z0Z_2\ : std_logic;
signal \ALU.mult_3_c6\ : std_logic;
signal \ALU.d_RNIJ0U031Z0Z_2\ : std_logic;
signal \ALU.d_RNIV1LMHZ0Z_3\ : std_logic;
signal \ALU.mult_3_c7\ : std_logic;
signal \ALU.d_RNIS69AHZ0Z_3\ : std_logic;
signal \ALU.d_RNI12A911Z0Z_2\ : std_logic;
signal \ALU.mult_3_c8\ : std_logic;
signal \ALU.d_RNINIF011Z0Z_2\ : std_logic;
signal \ALU.mult_3_c9\ : std_logic;
signal \ALU.mult_3_c10\ : std_logic;
signal \ALU.d_RNIINE1HZ0Z_3\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \ALU.d_RNIMCVI41Z0Z_2\ : std_logic;
signal \ALU.d_RNITCCHHZ0Z_3\ : std_logic;
signal \ALU.mult_3_c11\ : std_logic;
signal \ALU.d_RNI18J1JZ0Z_3\ : std_logic;
signal \ALU.mult_3_c12\ : std_logic;
signal \ALU.mult_3_c13\ : std_logic;
signal \ALU.mult_3_c14\ : std_logic;
signal \ALU.d_RNI2IA441Z0Z_2\ : std_logic;
signal \ALU.d_RNI7SQI21Z0Z_2\ : std_logic;
signal \ALU.d_RNID31VFZ0Z_3\ : std_logic;
signal \ALU.d_RNIBRFE41Z0Z_2\ : std_logic;
signal \ALU.d_RNI9IN2HZ0Z_3\ : std_logic;
signal \ALU.a_RNI2N741Z0Z_12\ : std_logic;
signal \ALU.d_RNIJRM75Z0Z_5\ : std_logic;
signal \DROM_ROMDATA_dintern_5ro\ : std_logic;
signal \ALU.d_RNIC0VE6Z0Z_5\ : std_logic;
signal \ALU.d_RNI693UNZ0Z_3\ : std_logic;
signal \ALU.mult_95_c_RNOZ0Z_0\ : std_logic;
signal \ALU.dout_6_ns_1_11_cascade_\ : std_logic;
signal \ALU.N_1144\ : std_logic;
signal \ALU.N_1096_cascade_\ : std_logic;
signal \DROM_ROMDATA_dintern_11ro\ : std_logic;
signal \aluOut_11_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_11_cascade_\ : std_logic;
signal \ALU.b_RNI2TJC1Z0Z_11\ : std_logic;
signal \ALU.operand2_11_cascade_\ : std_logic;
signal \ALU.d_RNIMR627Z0Z_11_cascade_\ : std_logic;
signal \ALU.a_RNIV5PUZ0Z_11\ : std_logic;
signal \ALU.c_RNI3MHFZ0Z_11\ : std_logic;
signal \ALU.dout_3_ns_1_11\ : std_logic;
signal \ALU.dout_3_ns_1_10_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_10_cascade_\ : std_logic;
signal \ALU.N_1143_cascade_\ : std_logic;
signal \ALU.N_1095\ : std_logic;
signal \aluOut_10_cascade_\ : std_logic;
signal \CONTROL.bus_0_10\ : std_logic;
signal \ALU_N_1141\ : std_logic;
signal \ALU_N_1093\ : std_logic;
signal \INVCONTROL.dout_7C_net\ : std_logic;
signal \gpuOut_c_7\ : std_logic;
signal \N_168\ : std_logic;
signal \N_168_cascade_\ : std_logic;
signal \D7_in_c\ : std_logic;
signal \CONTROL.bus_7_ns_1_7_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_23ro\ : std_logic;
signal \CONTROL.bus_7_a1_1_8_cascade_\ : std_logic;
signal \CONTROL.bus_sx_8\ : std_logic;
signal \gpuAddress_2\ : std_logic;
signal \gpuAddress_3\ : std_logic;
signal \gpuAddress_4\ : std_logic;
signal \gpuAddress_5\ : std_logic;
signal \gpuAddress_6\ : std_logic;
signal \gpuAddress_7\ : std_logic;
signal \gpuAddress_8\ : std_logic;
signal \INVCONTROL.gpuAddReg_2C_net\ : std_logic;
signal \CONTROL.un1_busState119_1_i_0_1_cascade_\ : std_logic;
signal \CONTROL.gpuWrite_RNOZ0Z_2_cascade_\ : std_logic;
signal \CONTROL.busState96_cascade_\ : std_logic;
signal \CONTROL.busState96\ : std_logic;
signal \CONTROL.N_66_0\ : std_logic;
signal \CONTROL.gpuWrite_RNOZ0Z_0\ : std_logic;
signal \gpuWrite\ : std_logic;
signal \INVCONTROL.gpuWriteC_net\ : std_logic;
signal \controlWord_21\ : std_logic;
signal \RAM.un1_WR_105_0Z0Z_3_cascade_\ : std_logic;
signal \A5_c\ : std_logic;
signal \RAM.un1_WR_105_0Z0Z_11\ : std_logic;
signal \controlWord_23\ : std_logic;
signal \A7_c\ : std_logic;
signal \controlWord_18\ : std_logic;
signal \controlWord_18_cascade_\ : std_logic;
signal \A2_c\ : std_logic;
signal \INVCONTROL.ramAddReg_5C_net\ : std_logic;
signal \CONTROL.g0_3_i_1_0_cascade_\ : std_logic;
signal \CONTROL.N_4_1_cascade_\ : std_logic;
signal \INVCONTROL.addrstackptr_4C_net\ : std_logic;
signal \CONTROL.N_81_0\ : std_logic;
signal \CONTROL.g0_3_i_a7_2_0\ : std_logic;
signal \CONTROL.N_429\ : std_logic;
signal \CONTROL.dout_reto_8\ : std_logic;
signal \progRomAddress_15\ : std_logic;
signal \CONTROL.programCounter_1_11\ : std_logic;
signal \CONTROL.addrstack_1_4\ : std_logic;
signal \CONTROL.N_4_1\ : std_logic;
signal \CONTROL.un1_addrstackptr_c4_0\ : std_logic;
signal \CONTROL.addrstackptr_8_4\ : std_logic;
signal \CONTROL.programCounter_1_14\ : std_logic;
signal \CONTROL.programCounter_1_reto_14\ : std_logic;
signal \CONTROL.programCounter_1_reto_11\ : std_logic;
signal \CONTROL.dout_reto_11\ : std_logic;
signal \PROM.ROMDATA.m470_am\ : std_logic;
signal \CONTROL.dout_reto_14\ : std_logic;
signal \CONTROL.programCounter_1_10\ : std_logic;
signal \CONTROL.programCounter11_reto_rep1\ : std_logic;
signal \CONTROL.programCounter_1_reto_10\ : std_logic;
signal \CONTROL.N_425\ : std_logic;
signal \CONTROL.programCounter_1_axb_1\ : std_logic;
signal \CONTROL.addrstackptr_8_1\ : std_logic;
signal \CONTROL.addrstackptr_RNI19JNL91Z0Z_0\ : std_logic;
signal \CONTROL.dout_reto_9\ : std_logic;
signal \ALU.d_RNILJMRC1Z0Z_8_cascade_\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \ALU.mult_7_c7\ : std_logic;
signal \ALU.d_RNITLGILZ0Z_7\ : std_logic;
signal \ALU.mult_7_c8\ : std_logic;
signal \ALU.d_RNIUFQIGZ0Z_7\ : std_logic;
signal \ALU.d_RNI8JFO21Z0Z_6\ : std_logic;
signal \ALU.mult_7_c9\ : std_logic;
signal \ALU.d_RNIKHEQHZ0Z_7\ : std_logic;
signal \ALU.d_RNIK9E841Z0Z_6\ : std_logic;
signal \ALU.mult_7_c10\ : std_logic;
signal \ALU.d_RNI73D441Z0Z_6\ : std_logic;
signal \ALU.mult_7_c11\ : std_logic;
signal \ALU.d_RNI7BDMHZ0Z_7\ : std_logic;
signal \ALU.mult_7_c12\ : std_logic;
signal \ALU.d_RNIBLU321Z0Z_6\ : std_logic;
signal \ALU.mult_7_c13\ : std_logic;
signal \ALU.mult_7_c14\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \ALU.d_RNIHNHG61Z0Z_6\ : std_logic;
signal \ALU.d_RNI4LU7E1Z0Z_6\ : std_logic;
signal \ALU.d_RNIA6P2IZ0Z_7\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \ALU.mult_1_c1\ : std_logic;
signal \ALU.d_RNIFBJI61Z0Z_0\ : std_logic;
signal \ALU.mult_1_c2\ : std_logic;
signal \ALU.d_RNIIOGRGZ0Z_1\ : std_logic;
signal \ALU.d_RNI67HQ21Z0Z_0\ : std_logic;
signal \ALU.mult_1_c3\ : std_logic;
signal \ALU.d_RNI8Q43IZ0Z_1\ : std_logic;
signal \ALU.d_RNIITFA41Z0Z_0\ : std_logic;
signal \ALU.mult_1_c4\ : std_logic;
signal \ALU.d_RNI5NE641Z0Z_0\ : std_logic;
signal \ALU.d_RNIUEFBIZ0Z_1\ : std_logic;
signal \ALU.mult_1_c5\ : std_logic;
signal \ALU.d_RNIRJ3VHZ0Z_1\ : std_logic;
signal \ALU.mult_1_c6\ : std_logic;
signal \ALU.d_RNI990621Z0Z_0\ : std_logic;
signal \ALU.mult_1_c7\ : std_logic;
signal \ALU.mult_1_c8\ : std_logic;
signal \ALU.d_RNIH49MHZ0Z_1\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \ALU.d_RNISP66IZ0Z_1\ : std_logic;
signal \ALU.mult_1_c9\ : std_logic;
signal \ALU.d_RNI0LDMJZ0Z_1\ : std_logic;
signal \ALU.d_RNIK8R951Z0Z_0\ : std_logic;
signal \ALU.mult_1_c10\ : std_logic;
signal \ALU.mult_1_c11\ : std_logic;
signal \ALU.d_RNI9UI0KZ0Z_1\ : std_logic;
signal \ALU.mult_1_c12\ : std_logic;
signal \ALU.mult_1_c13\ : std_logic;
signal \ALU.mult_3_c14_THRU_CO\ : std_logic;
signal \ALU.d_RNI3D2O61Z0Z_2\ : std_logic;
signal \ALU.mult_1_c14\ : std_logic;
signal \ALU.d_RNI83GO51Z0Z_0\ : std_logic;
signal \ALU.d_RNIPIBO31Z0Z_0\ : std_logic;
signal \ALU.d_RNIIHC6LZ0Z_3\ : std_logic;
signal \ALU.d_RNITH0K51Z0Z_0\ : std_logic;
signal \ALU.d_RNI0H41KZ0Z_1\ : std_logic;
signal \ALU.d_RNIETL861Z0Z_0\ : std_logic;
signal \ALU.d_RNI8FM541Z0Z_0\ : std_logic;
signal \ALU.d_RNIGIF4D1Z0Z_2\ : std_logic;
signal \CONTROL_addrstack_reto_11\ : std_logic;
signal \N_426\ : std_logic;
signal \progRomAddress_11\ : std_logic;
signal \ALU.d_RNILJMRC1_0Z0Z_8\ : std_logic;
signal \ALU.combOperand2_1Z0Z_0_cascade_\ : std_logic;
signal dintern_adflt_3_x : std_logic;
signal \DROM_ROMDATA_dintern_0ro_cascade_\ : std_logic;
signal \CONTROL.bus_6_a0_sx_0\ : std_logic;
signal \ALU.mult_5_c_RNOZ0Z_0\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_NEW_0\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_OLDZ0Z_0\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C_net\ : std_logic;
signal \INVCONTROL.dout_14C_net\ : std_logic;
signal \gpuOut_c_14\ : std_logic;
signal \CONTROL.ctrlOut_14\ : std_logic;
signal \D14_in_c\ : std_logic;
signal \CONTROL.N_175_cascade_\ : std_logic;
signal \N_191_cascade_\ : std_logic;
signal \CONTROL.busState_1_RNIRA1I6Z0Z_2_cascade_\ : std_logic;
signal \ALU.d_RNI8VHNHZ0Z_1\ : std_logic;
signal \ALU.dout_3_ns_1_12_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_12_cascade_\ : std_logic;
signal \ALU.N_1097\ : std_logic;
signal \ALU.N_1145_cascade_\ : std_logic;
signal \aluOut_12_cascade_\ : std_logic;
signal \CONTROL.bus_0_12\ : std_logic;
signal \gpuOut_c_11\ : std_logic;
signal \D11_in_c\ : std_logic;
signal \CONTROL.N_172_cascade_\ : std_logic;
signal \N_188\ : std_logic;
signal \N_204\ : std_logic;
signal \N_188_cascade_\ : std_logic;
signal \CONTROL.ctrlOut_11\ : std_logic;
signal \INVCONTROL.dout_11C_net\ : std_logic;
signal \gpuOut_c_12\ : std_logic;
signal \D12_in_c\ : std_logic;
signal \CONTROL.N_173_cascade_\ : std_logic;
signal \CONTROL.N_189\ : std_logic;
signal \CONTROL.un1_busState14_1_i_o2_0_cascade_\ : std_logic;
signal \CONTROL.un1_busState12_2_i_a2_0_1_tz_0_cascade_\ : std_logic;
signal \CONTROL.N_244_cascade_\ : std_logic;
signal \INVCONTROL.aluReadBusC_net\ : std_logic;
signal \CONTROL.un1_busState14_1_i_o2_0\ : std_logic;
signal \CONTROL.aluReadBus_r_1\ : std_logic;
signal \CONTROL.un1_busState14_1_i_a2_1_iZ0Z_1\ : std_logic;
signal \CONTROL.N_244\ : std_logic;
signal \CONTROL.N_58\ : std_logic;
signal \CONTROL.N_89\ : std_logic;
signal \CONTROL.N_89_cascade_\ : std_logic;
signal \CONTROL.aluReadBus_1_sqmuxa_0_a2_0Z0Z_0_cascade_\ : std_logic;
signal \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_0\ : std_logic;
signal \gpuOut_c_10\ : std_logic;
signal \D10_in_c\ : std_logic;
signal \CONTROL.N_171_cascade_\ : std_logic;
signal \CONTROL.N_187\ : std_logic;
signal \INVCONTROL.dout_10C_net\ : std_logic;
signal \gpuOut_c_0\ : std_logic;
signal \D0_in_c\ : std_logic;
signal \CONTROL.N_161_cascade_\ : std_logic;
signal \PROM.ROMDATA.m520\ : std_logic;
signal \gpuOut_c_15\ : std_logic;
signal \N_176\ : std_logic;
signal \D15_in_c\ : std_logic;
signal \N_176_cascade_\ : std_logic;
signal \PROM.ROMDATA.m471_ns\ : std_logic;
signal \INVCONTROL.dout_15C_net\ : std_logic;
signal \gpuOut_c_8\ : std_logic;
signal \CONTROL.ctrlOut_8\ : std_logic;
signal \A0_c\ : std_logic;
signal \A1_c\ : std_logic;
signal \controlWord_26\ : std_logic;
signal \controlWord_27\ : std_logic;
signal \A10_c\ : std_logic;
signal \A11_c\ : std_logic;
signal \RAM.un1_WR_105_0Z0Z_9\ : std_logic;
signal \controlWord_25\ : std_logic;
signal \A9_c\ : std_logic;
signal \controlWord_24\ : std_logic;
signal \A8_c\ : std_logic;
signal \INVCONTROL.ramAddReg_0C_net\ : std_logic;
signal \CONTROL.g1_0\ : std_logic;
signal \CONTROL.addrstack_1_1\ : std_logic;
signal \CONTROL.g1_0_cascade_\ : std_logic;
signal \INVCONTROL.addrstackptr_1C_net\ : std_logic;
signal \CONTROL.g0_1_i_a6Z0Z_4_cascade_\ : std_logic;
signal \CONTROL.N_9\ : std_logic;
signal \CONTROL.g0_0_1\ : std_logic;
signal \CONTROL.N_366\ : std_logic;
signal \CONTROL.g0_1_i_3\ : std_logic;
signal \CONTROL.addrstack_15\ : std_logic;
signal \CONTROL.addrstack_reto_15\ : std_logic;
signal \controlWord_30\ : std_logic;
signal \INVCONTROL.ramAddReg_14C_net\ : std_logic;
signal \ALU.mult_173_c_RNOZ0Z_0\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \ALU.mult_5_c5\ : std_logic;
signal \ALU.d_RNIFGNR61Z0Z_4\ : std_logic;
signal \ALU.mult_5_c6\ : std_logic;
signal \ALU.d_RNICP0UGZ0Z_5\ : std_logic;
signal \ALU.d_RNI6CL331Z0Z_4\ : std_logic;
signal \ALU.mult_5_c7\ : std_logic;
signal \ALU.d_RNI2RK5IZ0Z_5\ : std_logic;
signal \ALU.mult_5_c8\ : std_logic;
signal \ALU.d_RNIOFVDIZ0Z_5\ : std_logic;
signal \ALU.d_RNI5SIF41Z0Z_4\ : std_logic;
signal \ALU.mult_5_c9\ : std_logic;
signal \ALU.d_RNILKJ1IZ0Z_5\ : std_logic;
signal \ALU.d_RNIJTUN21Z0Z_4\ : std_logic;
signal \ALU.mult_5_c10\ : std_logic;
signal \ALU.d_RNI6HBMGZ0Z_5\ : std_logic;
signal \ALU.d_RNI9E4F21Z0Z_4\ : std_logic;
signal \ALU.mult_5_c11\ : std_logic;
signal \ALU.mult_5_c12\ : std_logic;
signal \ALU.d_RNIB5POHZ0Z_5\ : std_logic;
signal \ALU.d_RNIPNF141Z0Z_4\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \ALU.d_RNI88K161Z0Z_4\ : std_logic;
signal \ALU.d_RNIMQM8IZ0Z_5\ : std_logic;
signal \ALU.mult_5_c13\ : std_logic;
signal \ALU.mult_7_c14_THRU_CO\ : std_logic;
signal \ALU.d_RNIKDVI51Z0Z_4\ : std_logic;
signal \ALU.d_RNIRU9M31Z0Z_6\ : std_logic;
signal \ALU.mult_5_c14\ : std_logic;
signal bus_0_12 : std_logic;
signal \ALU.mult_239_c_RNOZ0Z_0\ : std_logic;
signal \ALU.mult_239_c_RNOZ0\ : std_logic;
signal \ALU.mult_1_2\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \ALU.mult_1_3\ : std_logic;
signal \ALU.mult_17_c2\ : std_logic;
signal \ALU.mult_3_4\ : std_logic;
signal \ALU.mult_1_4\ : std_logic;
signal \ALU.mult_17_c3\ : std_logic;
signal \ALU.mult_1_5\ : std_logic;
signal \ALU.mult_3_5\ : std_logic;
signal \ALU.mult_17_c4\ : std_logic;
signal \ALU.mult_1_6\ : std_logic;
signal \ALU.mult_3_6\ : std_logic;
signal \ALU.mult_17_c5\ : std_logic;
signal \ALU.mult_1_7\ : std_logic;
signal \ALU.mult_3_7\ : std_logic;
signal \ALU.mult_17_c6\ : std_logic;
signal \ALU.mult_1_8\ : std_logic;
signal \ALU.mult_3_8\ : std_logic;
signal \ALU.mult_17_c7\ : std_logic;
signal \ALU.mult_1_9\ : std_logic;
signal \ALU.mult_3_9\ : std_logic;
signal \ALU.mult_17_c8\ : std_logic;
signal \ALU.mult_17_c9\ : std_logic;
signal \ALU.mult_3_10\ : std_logic;
signal \ALU.mult_1_10\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \ALU.mult_1_11\ : std_logic;
signal \ALU.mult_3_11\ : std_logic;
signal \ALU.mult_17_c10\ : std_logic;
signal \ALU.mult_1_12\ : std_logic;
signal \ALU.mult_3_12\ : std_logic;
signal \ALU.mult_17_c11\ : std_logic;
signal \ALU.mult_1_13\ : std_logic;
signal \ALU.mult_3_13\ : std_logic;
signal \ALU.mult_17_c12\ : std_logic;
signal \ALU.mult_1_14\ : std_logic;
signal \ALU.mult_3_14\ : std_logic;
signal \ALU.mult_17_c13\ : std_logic;
signal \ALU.mult_227_c_RNIBPRVZ0Z92\ : std_logic;
signal \ALU.mult_83_c_RNIKEU6BZ0Z2\ : std_logic;
signal \ALU.mult_17_c14\ : std_logic;
signal \ALU.d_RNIHU6RLZ0Z_1\ : std_logic;
signal \ALU.d_RNI2E4JE1Z0Z_4\ : std_logic;
signal \ALU.N_860\ : std_logic;
signal \ALU.mult_5_c_RNOZ0\ : std_logic;
signal \ALU.d_RNI290AE1Z0Z_0\ : std_logic;
signal \ALU.d_RNI5MTIOZ0Z_1\ : std_logic;
signal \busState_1_RNICT0U1_2_cascade_\ : std_logic;
signal \busState_1_RNICT0U1_2\ : std_logic;
signal \N_227_0_cascade_\ : std_logic;
signal \ALU.status_18_cry_2_c_RNOZ0\ : std_logic;
signal \DROM_ROMDATA_dintern_2ro\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_NEW_2\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_OLDZ0Z_2\ : std_logic;
signal \INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C_net\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_sr_enZ0\ : std_logic;
signal \ALU.eZ0Z_4\ : std_logic;
signal \ALU.eZ0Z_10\ : std_logic;
signal \ALU.eZ0Z_11\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ALU.dout_6_ns_1_6_cascade_\ : std_logic;
signal \ALU.eZ0Z_6\ : std_logic;
signal \ALU.dout_3_ns_1_6_cascade_\ : std_logic;
signal \ALU.N_1091_cascade_\ : std_logic;
signal \ALU.N_1139\ : std_logic;
signal \aluOut_6_cascade_\ : std_logic;
signal \ALU.d_RNIR3N75Z0Z_6\ : std_logic;
signal \ALU.dout_6_ns_1_1_cascade_\ : std_logic;
signal \ALU_N_1134_cascade_\ : std_logic;
signal \CONTROL.operand1_ne_RNIBQE03Z0Z_0\ : std_logic;
signal \busState_1_RNI9P5V3_2\ : std_logic;
signal \ALU.dout_3_ns_1_1_cascade_\ : std_logic;
signal \ALU_N_1086_cascade_\ : std_logic;
signal \ALU_N_1134\ : std_logic;
signal \INVCONTROL.operand1_ne_1C_net\ : std_logic;
signal \ALU.d_RNIHD7AOZ0Z_7\ : std_logic;
signal \CONTROL.operand1_ne_RNIHKCU2Z0Z_0_cascade_\ : std_logic;
signal \operand1_ne_RNIDN8E7_0\ : std_logic;
signal \ALU.dout_6_ns_1_0\ : std_logic;
signal \aluOperand1_2_rep1\ : std_logic;
signal \ALU.dout_3_ns_1_0_cascade_\ : std_logic;
signal \ALU_N_1085_cascade_\ : std_logic;
signal \CONTROL.operand1_ne_RNIHKCU2_0Z0Z_0\ : std_logic;
signal \ALU_N_1133\ : std_logic;
signal \ALU_N_1085\ : std_logic;
signal \ALU.operand2_3_ns_1_2_cascade_\ : std_logic;
signal \ALU.N_1199_cascade_\ : std_logic;
signal \ALU.N_1199\ : std_logic;
signal \ALU.c_RNIJ1JO4_0Z0Z_2_cascade_\ : std_logic;
signal \ALU.c_RNIJ1JO4Z0Z_2\ : std_logic;
signal \ALU.d_RNIARKGBZ0Z_2\ : std_logic;
signal \ALU.operand2_6_ns_1_2\ : std_logic;
signal \ALU.N_1247\ : std_logic;
signal \gpuOut_c_13\ : std_logic;
signal \D13_in_c\ : std_logic;
signal \CONTROL.N_174_cascade_\ : std_logic;
signal \CONTROL.N_169\ : std_logic;
signal \D8_in_c\ : std_logic;
signal \CONTROL.N_185\ : std_logic;
signal \INVCONTROL.busState_1_2C_net\ : std_logic;
signal \D4_in_c\ : std_logic;
signal \CONTROL.busState_1_RNIU83C1_0Z0Z_2\ : std_logic;
signal \D2_in_c\ : std_logic;
signal \N_228_0\ : std_logic;
signal \CONTROL.busState_1_RNILAEH1Z0Z_2\ : std_logic;
signal \gpuOut_c_1\ : std_logic;
signal \N_162\ : std_logic;
signal \D1_in_c\ : std_logic;
signal \N_162_cascade_\ : std_logic;
signal \INVCONTROL.busState_1_1C_net\ : std_logic;
signal \CONTROL.N_180\ : std_logic;
signal \gpuOut_c_3\ : std_logic;
signal \N_164\ : std_logic;
signal \D3_in_c\ : std_logic;
signal \N_164_cascade_\ : std_logic;
signal \controlWord_16\ : std_logic;
signal \CONTROL_romAddReg_7_0\ : std_logic;
signal \controlWord_17\ : std_logic;
signal \controlWord_17_cascade_\ : std_logic;
signal \CONTROL_romAddReg_7_1\ : std_logic;
signal \INVCONTROL.dout_1C_net\ : std_logic;
signal \CONTROL.N_430\ : std_logic;
signal \CONTROL.un1_busState98_1_1_0Z0Z_0\ : std_logic;
signal \CONTROL.programCounter_1_15\ : std_logic;
signal \CONTROL.programCounter_1_reto_15\ : std_logic;
signal \CONTROL.ctrlOut_15\ : std_logic;
signal \CONTROL.dout_reto_15\ : std_logic;
signal \PROM.ROMDATA.m465_am\ : std_logic;
signal \CONTROL.ctrlOut_7\ : std_logic;
signal \CONTROL.tempCounterZ0Z_0\ : std_logic;
signal \CONTROL.tempCounterZ0Z_5\ : std_logic;
signal \CONTROL.tempCounterZ0Z_3\ : std_logic;
signal \CONTROL.programCounter_1_8\ : std_logic;
signal \CONTROL.tempCounterZ0Z_8\ : std_logic;
signal \INVCONTROL.tempCounter_0C_net\ : std_logic;
signal \CONTROL.tempCounterZ0Z_4\ : std_logic;
signal \CONTROL.tempCounterZ0Z_1\ : std_logic;
signal \CONTROL.tempCounterZ0Z_7\ : std_logic;
signal \CONTROL.tempCounterZ0Z_12\ : std_logic;
signal \CONTROL.tempCounterZ0Z_2\ : std_logic;
signal \INVCONTROL.tempCounter_4C_net\ : std_logic;
signal \CONTROL.addrstack_1_i\ : std_logic;
signal \ALU.d_RNII2KJ41Z0Z_4\ : std_logic;
signal bus_4 : std_logic;
signal \ALU.mult_173_c_RNOZ0\ : std_logic;
signal \ALU.mult_5_6\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \ALU.mult_7_7\ : std_logic;
signal \ALU.mult_5_7\ : std_logic;
signal \ALU.mult_19_c6\ : std_logic;
signal \ALU.mult_7_8\ : std_logic;
signal \ALU.mult_5_8\ : std_logic;
signal \ALU.mult_19_c7\ : std_logic;
signal \ALU.mult_7_9\ : std_logic;
signal \ALU.mult_5_9\ : std_logic;
signal \ALU.mult_19_c8\ : std_logic;
signal \ALU.mult_7_10\ : std_logic;
signal \ALU.mult_5_10\ : std_logic;
signal \ALU.mult_19_c9\ : std_logic;
signal \ALU.mult_7_11\ : std_logic;
signal \ALU.mult_5_11\ : std_logic;
signal \ALU.mult_19_c10\ : std_logic;
signal \ALU.mult_5_12\ : std_logic;
signal \ALU.mult_7_12\ : std_logic;
signal \ALU.mult_19_c11\ : std_logic;
signal \ALU.mult_5_13\ : std_logic;
signal \ALU.mult_7_13\ : std_logic;
signal \ALU.mult_19_c12\ : std_logic;
signal \ALU.mult_19_c13\ : std_logic;
signal \ALU.mult_5_14\ : std_logic;
signal \ALU.mult_7_14\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \ALU.mult_19_c14\ : std_logic;
signal \ALU.mult_19_c14_THRU_CO\ : std_logic;
signal \ALU.mult_3_2\ : std_logic;
signal \ALU.mult_486_c_RNIPJD0IZ0Z5_cascade_\ : std_logic;
signal \ALU.combOperand2_0_5\ : std_logic;
signal \ALU.d_RNICGRJGZ0Z_1\ : std_logic;
signal \ALU.addsub_cry_4_c_RNI2RZ0Z6596\ : std_logic;
signal \ALU.d_RNIBVMTLZ0Z_5\ : std_logic;
signal \ALU.d_RNIVMDLOZ0Z_5\ : std_logic;
signal \ALU.mult_3_3\ : std_logic;
signal \busState_1_RNIBS0U1_2\ : std_logic;
signal \operand1_ne_RNIR8FK7_0\ : std_logic;
signal \ALU.status_19_0_cascade_\ : std_logic;
signal \ALU.mult_95_c_RNOZ0\ : std_logic;
signal \ALU.mult_3\ : std_logic;
signal \ALU.addsub_cry_2_c_RNIUFTGNZ0Z3_cascade_\ : std_logic;
signal \ALU.mult_388_c_RNIBULDPZ0Z3\ : std_logic;
signal \ALU.mult_388_c_RNIEAAJHZ0Z7_cascade_\ : std_logic;
signal bus_3 : std_logic;
signal \ALU.mult_388_c_RNIEAAJHZ0Z7\ : std_logic;
signal \ALU.mult_388_c_RNIPGN6QZ0Z7_cascade_\ : std_logic;
signal \ALU.a_15_d_sZ0Z_5\ : std_logic;
signal \ALU.mult_2\ : std_logic;
signal \ALU.log_1_2\ : std_logic;
signal \ALU.a_15_d_sZ0Z_3\ : std_logic;
signal \ALU.addsub_cry_1_c_RNI8FKPLZ0Z3_cascade_\ : std_logic;
signal \ALU.mult_5_c_RNI6ET5DZ0Z3\ : std_logic;
signal \ALU.addsub_cry_1_c_RNIJP8KZ0Z37_cascade_\ : std_logic;
signal \ALU.addsub_cry_1_c_RNIJP8KZ0Z37\ : std_logic;
signal \ALU.addsub_cry_1_c_RNIICPECZ0Z7_cascade_\ : std_logic;
signal \ALU.dout_3_ns_1_9_cascade_\ : std_logic;
signal \ALU.dout_6_ns_1_9_cascade_\ : std_logic;
signal \ALU.N_1094\ : std_logic;
signal \ALU.N_1142_cascade_\ : std_logic;
signal \aluOut_9_cascade_\ : std_logic;
signal h_2 : std_logic;
signal \ALU.dout_6_ns_1_2_cascade_\ : std_logic;
signal \ALU.aZ0Z_2\ : std_logic;
signal \ALU.eZ0Z_2\ : std_logic;
signal \ALU.dout_3_ns_1_2_cascade_\ : std_logic;
signal \ALU.N_1087_cascade_\ : std_logic;
signal \ALU.N_1135\ : std_logic;
signal \ALU_N_1086\ : std_logic;
signal \CONTROL.operand1_ne_RNIBQE03_0Z0Z_0\ : std_logic;
signal \PROM.ROMDATA.m238_am_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m238_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m244_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m244_ns_1\ : std_logic;
signal \INVCONTROL.operand1_fast_ne_1C_net\ : std_logic;
signal \ALU.dout_6_ns_1_3_cascade_\ : std_logic;
signal \ALU.dout_3_ns_1_3_cascade_\ : std_logic;
signal \ALU.N_1136\ : std_logic;
signal \ALU.N_1088_cascade_\ : std_logic;
signal \aluOut_3_cascade_\ : std_logic;
signal \busState_1_RNIH16V3_2\ : std_logic;
signal \ALU.dout_3_ns_1_13_cascade_\ : std_logic;
signal \aluOperand1_2_rep2\ : std_logic;
signal \ALU.dout_6_ns_1_13_cascade_\ : std_logic;
signal \ALU.N_1098\ : std_logic;
signal \ALU.N_1146_cascade_\ : std_logic;
signal \CONTROL.N_190\ : std_logic;
signal \CONTROL.bus_7_a1_1_8\ : std_logic;
signal \aluOut_13_cascade_\ : std_logic;
signal \CONTROL.bus_0_13\ : std_logic;
signal \ALU.c_RNIJMOB4_0Z0Z_1_cascade_\ : std_logic;
signal \ALU.d_RNID42JAZ0Z_1\ : std_logic;
signal \ALU.operand2_6_ns_1_1\ : std_logic;
signal \ALU.N_1246\ : std_logic;
signal \ALU.operand2_3_ns_1_1_cascade_\ : std_logic;
signal \ALU.N_1198\ : std_logic;
signal \ALU.combOperand2_d_bmZ0Z_1\ : std_logic;
signal \ALU.N_1198_cascade_\ : std_logic;
signal \ALU.c_RNIJMOB4Z0Z_1\ : std_logic;
signal \CONTROL.g0_3_i_a7_2_1\ : std_logic;
signal \CONTROL.N_5_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_8_3\ : std_logic;
signal \gpuOut_c_2\ : std_logic;
signal \CONTROL.N_163\ : std_logic;
signal \CONTROL.g0_3_i_2_1\ : std_logic;
signal \CONTROL.un1_addrstackptr_c3_0\ : std_logic;
signal \CONTROL.addrstack_1_3\ : std_logic;
signal \CONTROL.N_5\ : std_logic;
signal \CONTROL.addrstackptrZ0Z_3\ : std_logic;
signal \INVCONTROL.addrstackptr_3C_net\ : std_logic;
signal \INVCONTROL.aluOperation_ne_1C_net\ : std_logic;
signal \CONTROL.N_83_0_cascade_\ : std_logic;
signal \CONTROL.m28_0_120_i_i_4\ : std_logic;
signal \CONTROL.N_75_0\ : std_logic;
signal \CONTROL.N_75_0_cascade_\ : std_logic;
signal \CONTROL.m38_i_2\ : std_logic;
signal \CONTROL.N_339\ : std_logic;
signal \CONTROL.N_219_cascade_\ : std_logic;
signal \CONTROL.m28_0_120_i_i_a2_0_0_cascade_\ : std_logic;
signal \CONTROL.busState_1_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \CONTROL.busState_1_RNO_0Z0Z_1\ : std_logic;
signal \CONTROL.g0_3_i_1_1\ : std_logic;
signal \CONTROL.N_350_1\ : std_logic;
signal \CONTROL.N_345\ : std_logic;
signal \CONTROL.N_346\ : std_logic;
signal \CONTROL.N_255\ : std_logic;
signal \CONTROL.N_345_cascade_\ : std_logic;
signal \ramWrite\ : std_logic;
signal \INVCONTROL.ramWriteC_net\ : std_logic;
signal \CONTROL.un1_busState114_1_0Z0Z_0\ : std_logic;
signal \CONTROL.ctrlOut_10\ : std_logic;
signal \CONTROL.dout_reto_10\ : std_logic;
signal \PROM.ROMDATA.m1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m2_cascade_\ : std_logic;
signal \ALU.mult_7_6\ : std_logic;
signal \ALU.status_18_cry_0_c_RNOZ0\ : std_logic;
signal \ALU.mult_5_4\ : std_logic;
signal \ALU.mult_17_4\ : std_logic;
signal \ALU.mult_391_c_RNIEC73TZ0Z4\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \ALU.mult_17_5\ : std_logic;
signal \ALU.mult_5\ : std_logic;
signal \ALU.mult_25_c4\ : std_logic;
signal \ALU.mult_173_c_RNIO8AOZ0Z16\ : std_logic;
signal \ALU.mult_17_6\ : std_logic;
signal \ALU.mult_25_c5\ : std_logic;
signal \ALU.mult_19_7\ : std_logic;
signal \ALU.mult_17_7\ : std_logic;
signal \ALU.mult_25_c6\ : std_logic;
signal \ALU.mult_17_8\ : std_logic;
signal \ALU.mult_19_8\ : std_logic;
signal \ALU.mult_25_c7\ : std_logic;
signal \ALU.mult_17_9\ : std_logic;
signal \ALU.mult_19_9\ : std_logic;
signal \ALU.mult_25_c8\ : std_logic;
signal \ALU.mult_19_10\ : std_logic;
signal \ALU.mult_17_10\ : std_logic;
signal \ALU.mult_25_c9\ : std_logic;
signal \ALU.mult_17_11\ : std_logic;
signal \ALU.mult_19_11\ : std_logic;
signal \ALU.mult_25_c10\ : std_logic;
signal \ALU.mult_25_c11\ : std_logic;
signal \ALU.mult_17_12\ : std_logic;
signal \ALU.mult_19_12\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \ALU.mult_17_13\ : std_logic;
signal \ALU.mult_19_13\ : std_logic;
signal \ALU.mult_25_c12\ : std_logic;
signal \ALU.mult_17_14\ : std_logic;
signal \ALU.mult_19_14\ : std_logic;
signal \ALU.mult_25_c13\ : std_logic;
signal \ALU.mult_424_c_RNIUVTALZ0Z4\ : std_logic;
signal \ALU.mult_25_c14\ : std_logic;
signal \ALU.d_RNIUT8OG4Z0Z_0\ : std_logic;
signal \ALU.lshift_3_ns_1_14\ : std_logic;
signal \ALU.N_646_cascade_\ : std_logic;
signal \ALU.lshift_15_ns_1_14_cascade_\ : std_logic;
signal g_2 : std_logic;
signal g_4 : std_logic;
signal g_6 : std_logic;
signal g_10 : std_logic;
signal g_11 : std_logic;
signal f_2 : std_logic;
signal f_10 : std_logic;
signal f_11 : std_logic;
signal \CONSTANT_ZERO_NET\ : std_logic;
signal \ALU.cZ0Z_2\ : std_logic;
signal \ALU.cZ0Z_4\ : std_logic;
signal \ALU.cZ0Z_6\ : std_logic;
signal \ALU.cZ0Z_10\ : std_logic;
signal \ALU.cZ0Z_11\ : std_logic;
signal \ALU.dZ0Z_2\ : std_logic;
signal \ALU.dZ0Z_6\ : std_logic;
signal \ALU.dZ0Z_10\ : std_logic;
signal \ALU.dZ0Z_11\ : std_logic;
signal \ALU.d_RNI6DCTZ0Z_11\ : std_logic;
signal \INVCONTROL.operand2_fast_ne_2C_net\ : std_logic;
signal \ALU.N_920\ : std_logic;
signal \ALU.operand2_3_ns_1_15\ : std_logic;
signal \ALU.dout_3_ns_1_15_cascade_\ : std_logic;
signal \aluOperand1_fast_2\ : std_logic;
signal \aluOperand1_fast_1\ : std_logic;
signal \CONTROL.increment28lto5_1_1_3\ : std_logic;
signal \CONTROL.increment28lto5_1_1_1_cascade_\ : std_logic;
signal \CONTROL.g0_3_i_a7Z0Z_3\ : std_logic;
signal \PROM.ROMDATA.m221cf1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m221cf1\ : std_logic;
signal \INVCONTROL.operand1_ne_0C_net\ : std_logic;
signal \CONTROL.un1_busState98_1_0_0_0\ : std_logic;
signal \PROM.ROMDATA.m217\ : std_logic;
signal \PROM.ROMDATA.m221cf0\ : std_logic;
signal \CONTROL.increment28lto5_1_1_0\ : std_logic;
signal \CONTROL.N_101_0\ : std_logic;
signal \CONTROL.N_320_cascade_\ : std_logic;
signal \CONTROL.un1_busState103_0_0_cascade_\ : std_logic;
signal \INVCONTROL.aluParams_1_0C_net\ : std_logic;
signal \CONTROL.N_95_0\ : std_logic;
signal \CONTROL.N_318\ : std_logic;
signal \CONTROL.N_340_cascade_\ : std_logic;
signal \INVCONTROL.aluParams_1_ne_1C_net\ : std_logic;
signal \CONTROL.un1_busState103_0_0\ : std_logic;
signal \CONTROL.un1_busState114_2_0_0_xZ0Z0_cascade_\ : std_logic;
signal \CONTROL.un1_busState114_2_0_0_xZ0Z1\ : std_logic;
signal \CONTROL.un1_busState114_2_0_0_0_cascade_\ : std_logic;
signal \CONTROL.aluReadBus_1_sqmuxa_0_a2_2Z0Z_0\ : std_logic;
signal \CONTROL.N_83_0\ : std_logic;
signal \CONTROL.N_48_0_cascade_\ : std_logic;
signal \INVCONTROL.aluOperation_4C_net\ : std_logic;
signal \CONTROL.un1_controlWord_14_i_0\ : std_logic;
signal \CONTROL.N_87_0\ : std_logic;
signal \CONTROL.un1_busState97_1_0_1_0\ : std_logic;
signal \CONTROL.dout_reto_7\ : std_logic;
signal \CONTROL.addrstack_reto_7\ : std_logic;
signal \CONTROL.N_422_cascade_\ : std_logic;
signal \progRomAddress_7_cascade_\ : std_logic;
signal \INVCONTROL.dout_2C_net\ : std_logic;
signal \CONTROL.N_420_cascade_\ : std_logic;
signal \CONTROL.programCounter_1_axb_5\ : std_logic;
signal \CONTROL.programCounter_1_axb_0\ : std_logic;
signal \CONTROL.N_105_i\ : std_logic;
signal \CONTROL.N_427\ : std_logic;
signal \PROM_ROMDATA_dintern_5ro_cascade_\ : std_logic;
signal \CONTROL.N_80_0\ : std_logic;
signal \CONTROL.g0_1_i_3Z0Z_1\ : std_logic;
signal \CONTROL.N_384_0\ : std_logic;
signal \CONTROL.N_209_cascade_\ : std_logic;
signal \CONTROL.un1_busState114_1_0_0_0\ : std_logic;
signal \CONTROL.N_349_cascade_\ : std_logic;
signal \CONTROL.N_246\ : std_logic;
signal \CONTROL.m38_i_1\ : std_logic;
signal \CONTROL.N_348\ : std_logic;
signal \CONTROL.programCounter_1_12\ : std_logic;
signal \CONTROL.programCounter_1_reto_12\ : std_logic;
signal \controlWord_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m506_cascade_\ : std_logic;
signal \PROM.ROMDATA.N_571_mux\ : std_logic;
signal \N_177\ : std_logic;
signal \ALU.d_RNI64MA6Z0Z_0_cascade_\ : std_logic;
signal \ALU.log_1_3_ns_1_1_0_cascade_\ : std_logic;
signal \ALU.log_1_3_ns_1_0_cascade_\ : std_logic;
signal \ALU.log_1_0_cascade_\ : std_logic;
signal \ALU.status_8_5_0_cascade_\ : std_logic;
signal \ALU.mult_365_c_RNOZ0\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \ALU.c_RNIF6GEF1Z0Z_12\ : std_logic;
signal \ALU.c_RNINUT6PZ0Z_13\ : std_logic;
signal \ALU.mult_13_c13\ : std_logic;
signal \ALU.c_RNIS83N71Z0Z_12\ : std_logic;
signal \ALU.mult_13_c14\ : std_logic;
signal \ALU.d_RNIL4PC21Z0Z_6\ : std_logic;
signal \ALU.mult_5_5\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \ALU.mult_9_9\ : std_logic;
signal \ALU.mult_25_9\ : std_logic;
signal \ALU.mult_29_c8\ : std_logic;
signal \ALU.mult_29_c9\ : std_logic;
signal \ALU.mult_25_11\ : std_logic;
signal \ALU.mult_29_c10\ : std_logic;
signal \ALU.mult_29_c11\ : std_logic;
signal \ALU.mult_25_13\ : std_logic;
signal \ALU.mult_29_c12\ : std_logic;
signal \ALU.mult_25_14\ : std_logic;
signal \ALU.mult_29_c13\ : std_logic;
signal \ALU.mult_516_c_RNI98SKDCZ0\ : std_logic;
signal \ALU.mult_29_c14\ : std_logic;
signal bus_0_10 : std_logic;
signal \ALU.mult_10\ : std_logic;
signal \ALU.mult_549_c_RNIB6TIDGZ0_cascade_\ : std_logic;
signal \ALU.a_15_am_1_10\ : std_logic;
signal \ALU.mult_549_c_RNIE7260OZ0_cascade_\ : std_logic;
signal \ALU.aZ0Z_10\ : std_logic;
signal \ALU.a_15_m3_sZ0Z_13_cascade_\ : std_logic;
signal \ALU.a32Z0Z_0_cascade_\ : std_logic;
signal \ALU.aZ0Z_1\ : std_logic;
signal \ALU.d_RNICUA7B5Z0Z_0_cascade_\ : std_logic;
signal \ALU.d_RNIL3JT71Z0Z_0\ : std_logic;
signal \ALU.N_556\ : std_logic;
signal \ALU.N_556_cascade_\ : std_logic;
signal \ALU.d_RNI3MGBH1Z0Z_1\ : std_logic;
signal \ALU.status_17_I_39_c_RNOZ0\ : std_logic;
signal \ALU.mult_365_c_RNOZ0Z_0\ : std_logic;
signal \ALU.N_572\ : std_logic;
signal bus_11 : std_logic;
signal \ALU.mult_11\ : std_logic;
signal \ALU.mult_552_c_RNI70R9DAZ0_cascade_\ : std_logic;
signal \ALU.rshift_11\ : std_logic;
signal \ALU.a_15_am_rn_0_11\ : std_logic;
signal \ALU.mult_552_c_RNI70R9DAZ0\ : std_logic;
signal \ALU.mult_552_c_RNIOT7VLFZ0_cascade_\ : std_logic;
signal \ALU.aZ0Z_11\ : std_logic;
signal \ALU.a_15_am_snZ0Z_11\ : std_logic;
signal h_1 : std_logic;
signal \ALU.mult_6\ : std_logic;
signal \ALU.mult_489_c_RNIGEUL1AZ0_cascade_\ : std_logic;
signal \ALU.mult_489_c_RNIGEUL1AZ0\ : std_logic;
signal \ALU.mult_489_c_RNIPGBQMCZ0Z_0_cascade_\ : std_logic;
signal \ALU.mult_489_c_RNIPGBQMCZ0\ : std_logic;
signal \ALU.mult_489_c_RNI1J3GCUZ0_cascade_\ : std_logic;
signal h_6 : std_logic;
signal \ALU.a_15_m2_d_d_ns_1_0_0_cascade_\ : std_logic;
signal bus_0 : std_logic;
signal \ALU.lshift62\ : std_logic;
signal \ALU.d_RNI4D6E01Z0Z_0_cascade_\ : std_logic;
signal \ALU.d_RNIQQ9O83Z0Z_0_cascade_\ : std_logic;
signal \ALU.d_RNI4HL061Z0Z_0\ : std_logic;
signal \ALU.d_RNINUGCF4Z0Z_0_cascade_\ : std_logic;
signal \ALU.aZ0Z_0\ : std_logic;
signal h_0 : std_logic;
signal \ALU.e_RNI933SZ0Z_0\ : std_logic;
signal \ALU.c_RNIDFF01Z0Z_0_cascade_\ : std_logic;
signal \ALU.d_RNI0G5DZ0Z_0\ : std_logic;
signal \ALU.b_RNIS3POZ0Z_0_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_0\ : std_logic;
signal \ALU.operand2_0\ : std_logic;
signal \ALU.dZ0Z_3\ : std_logic;
signal \ALU.operand2_6_ns_1_3_cascade_\ : std_logic;
signal \ALU.aZ0Z_3\ : std_logic;
signal \ALU.eZ0Z_3\ : std_logic;
signal \ALU.cZ0Z_3\ : std_logic;
signal g_3 : std_logic;
signal \ALU.operand2_3_ns_1_3_cascade_\ : std_logic;
signal \ALU.N_1200_cascade_\ : std_logic;
signal \ALU.N_1248\ : std_logic;
signal \ALU.d_RNIGMEO4Z0Z_3_cascade_\ : std_logic;
signal \ALU.combOperand2_d_bmZ0Z_3\ : std_logic;
signal \ALU.d_RNI2CUG6Z0Z_3\ : std_logic;
signal \gpuOut_c_4\ : std_logic;
signal \CONTROL.N_165\ : std_logic;
signal h_9 : std_logic;
signal \ALU.e_RNICGJMZ0Z_9\ : std_logic;
signal \ALU.d_RNIKKNJZ0Z_9\ : std_logic;
signal \ALU.operand2_7_ns_1_9_cascade_\ : std_logic;
signal \ALU.b_RNIG8BVZ0Z_9\ : std_logic;
signal \ALU.operand2_9_cascade_\ : std_logic;
signal \ALU.status_RNO_2Z0Z_0\ : std_logic;
signal \ALU.status_e_1_0\ : std_logic;
signal \CONTROL.increment28lto5_1Z0Z_1_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_8ro\ : std_logic;
signal \CONTROL.increment28lto5_1_1_2_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_7ro\ : std_logic;
signal \CONTROL.increment28lto5_1Z0Z_2\ : std_logic;
signal \INVCONTROL.aluOperation_ne_5C_net\ : std_logic;
signal \CONTROL.N_48_0\ : std_logic;
signal \controlWord_6_cascade_\ : std_logic;
signal \CONTROL.N_140_0\ : std_logic;
signal \CONTROL.un1_busState96_1_i_i_a2_1Z0Z_1_cascade_\ : std_logic;
signal \CONTROL.un1_busState96_1_i_i_a2_0Z0Z_1\ : std_logic;
signal \CONTROL.un1_busState96_1_i_iZ0Z_0_cascade_\ : std_logic;
signal \controlWord_5_cascade_\ : std_logic;
signal \CONTROL.N_134_0\ : std_logic;
signal \CONTROL.N_327\ : std_logic;
signal \CONTROL.N_133_0_1\ : std_logic;
signal \PROM_ROMDATA_dintern_3ro_cascade_\ : std_logic;
signal \CONTROL.g0_3_i_2_0\ : std_logic;
signal \CONTROL.g0_2_i_a7Z0Z_3\ : std_logic;
signal \CONTROL.g0_2_i_a7Z0Z_2\ : std_logic;
signal \CONTROL.g0_2_i_2_cascade_\ : std_logic;
signal \CONTROL.addrstack_1_2\ : std_logic;
signal \CONTROL.addrstackptrZ0Z_1\ : std_logic;
signal \CONTROL.N_5_0_cascade_\ : std_logic;
signal \CONTROL.g0_12_1_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_8_2\ : std_logic;
signal \controlWord_4_cascade_\ : std_logic;
signal \CONTROL.N_5_0\ : std_logic;
signal \CONTROL.g0_12_1\ : std_logic;
signal \INVCONTROL.addrstackptr_2C_net\ : std_logic;
signal \CONTROL.N_360\ : std_logic;
signal \CONTROL.N_362\ : std_logic;
signal \CONTROL.m28_0_120_i_i_0\ : std_logic;
signal \CONTROL.N_321\ : std_logic;
signal \CONTROL.N_338\ : std_logic;
signal \PROM_ROMDATA_dintern_0ro\ : std_logic;
signal \PROM_ROMDATA_dintern_0ro_cascade_\ : std_logic;
signal \CONTROL.un1_busState_0_sqmuxa_i_a2_0\ : std_logic;
signal \CONTROL.N_304_0\ : std_logic;
signal \PROM.ROMDATA.m433_ns\ : std_logic;
signal \PROM.ROMDATA.m294_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m31_cascade_\ : std_logic;
signal \CONTROL.ctrlOut_12\ : std_logic;
signal \CONTROL.dout_reto_12\ : std_logic;
signal \PROM.ROMDATA.m391_cascade_\ : std_logic;
signal \PROM.ROMDATA.m433_bm\ : std_logic;
signal \PROM.ROMDATA.m382_ns\ : std_logic;
signal \busState_1_RNIAR0U1_2\ : std_logic;
signal \N_225_0_cascade_\ : std_logic;
signal \ALU.mult_13_15\ : std_logic;
signal \ALU.mult_15_14_cascade_\ : std_logic;
signal \ALU.mult_13_14\ : std_logic;
signal \ALU.lshift_3_ns_1_15_cascade_\ : std_logic;
signal \ALU.d_RNI64MA6Z0Z_0\ : std_logic;
signal \N_225_0\ : std_logic;
signal \ALU.mult_25_12\ : std_logic;
signal \ALU.mult_13_12_cascade_\ : std_logic;
signal \ALU.mult_467_c_RNICRDK6BZ0\ : std_logic;
signal \ALU.mult_13_12\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \ALU.mult_13_13\ : std_logic;
signal \ALU.mult_27_13\ : std_logic;
signal \ALU.mult_27_c12\ : std_logic;
signal \ALU.mult_365_c_RNI8ALOZ0Z96\ : std_logic;
signal \ALU.mult_27_14\ : std_logic;
signal \ALU.mult_27_c13\ : std_logic;
signal \ALU.mult_27_c14\ : std_logic;
signal \ALU.mult_27_c14_THRU_CO\ : std_logic;
signal \ALU.mult_9\ : std_logic;
signal \ALU.mult_13\ : std_logic;
signal \ALU.N_642\ : std_logic;
signal \ALU.d_RNIULN025Z0Z_2_cascade_\ : std_logic;
signal \ALU.d_RNIULN025_0Z0Z_2\ : std_logic;
signal \ALU.lshift_10_cascade_\ : std_logic;
signal \ALU.c_RNIO0KOKEZ0Z_10_cascade_\ : std_logic;
signal \ALU.bZ0Z_10\ : std_logic;
signal \ALU.N_1025\ : std_logic;
signal \ALU.N_864\ : std_logic;
signal \ALU.N_965_cascade_\ : std_logic;
signal \ALU.d_RNIFHCRU4Z0Z_2\ : std_logic;
signal \ALU.mult_15_15\ : std_logic;
signal \ALU.c_RNINT9PO2Z0Z_10\ : std_logic;
signal \ALU.c_RNI890LZ0Z_13\ : std_logic;
signal \ALU.a_RNI4P741Z0Z_13_cascade_\ : std_logic;
signal \ALU.d_RNIAHCTZ0Z_13\ : std_logic;
signal \ALU.operand2_7_ns_1_13_cascade_\ : std_logic;
signal \ALU.b_RNI61KC1Z0Z_13\ : std_logic;
signal \ALU.operand2_13\ : std_logic;
signal bus_0_13 : std_logic;
signal \ALU.operand2_13_cascade_\ : std_logic;
signal \ALU.d_RNI02EVNBZ0Z_4\ : std_logic;
signal \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\ : std_logic;
signal \ALU.addsub_cry_1_c_RNIICPECZ0Z7\ : std_logic;
signal \ALU.bZ0Z_2\ : std_logic;
signal \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9\ : std_logic;
signal \ALU.addsub_cry_4_c_RNI5L6IQAZ0\ : std_logic;
signal \ALU.bZ0Z_6\ : std_logic;
signal \ALU.bZ0Z_3\ : std_logic;
signal \ALU.bZ0Z_11\ : std_logic;
signal \ALU.bZ0Z_12\ : std_logic;
signal \CONTROL.gZ0Z3\ : std_logic;
signal \ALU.lshift_15_0_sx_1\ : std_logic;
signal bus_14 : std_logic;
signal \ALU.lshift_15_0_1_cascade_\ : std_logic;
signal \ALU.a_15_m0_sx_14\ : std_logic;
signal \ALU.lshift_15_0_1\ : std_logic;
signal \ALU.mult_1_cascade_\ : std_logic;
signal \ALU.a_15_m3_d_ns_1_1\ : std_logic;
signal \ALU.d_RNIJOQE21Z0Z_0\ : std_logic;
signal g_5 : std_logic;
signal \ALU.cZ0Z_5\ : std_logic;
signal \ALU.eZ0Z_5\ : std_logic;
signal \ALU.aZ0Z_5\ : std_logic;
signal \ALU.c_RNI8KVQZ0Z_5\ : std_logic;
signal \ALU.e_RNI48JMZ0Z_5_cascade_\ : std_logic;
signal \ALU.operand2_7_ns_1_5_cascade_\ : std_logic;
signal \ALU.operand2_5\ : std_logic;
signal f_5 : std_logic;
signal \ALU.bZ0Z_5\ : std_logic;
signal \ALU.b_RNI7HSPZ0Z_5\ : std_logic;
signal h_5 : std_logic;
signal \ALU.dZ0Z_5\ : std_logic;
signal \ALU.d_RNIBT8EZ0Z_5\ : std_logic;
signal \INVCONTROL.operand2_2_rep1_neC_net\ : std_logic;
signal \PROM.ROMDATA.m407_cascade_\ : std_logic;
signal \PROM.ROMDATA.m488_ns_cascade_\ : std_logic;
signal \INVCONTROL.operand2_fast_ne_1C_net\ : std_logic;
signal \CONTROL.aluReadBus_1_sqmuxa\ : std_logic;
signal \ALU.un14_log_a0_2Z0Z_15\ : std_logic;
signal \ALU.d_RNIN8NU4Z0Z_9\ : std_logic;
signal \ALU.combOperand2_0_0_9\ : std_logic;
signal \DROM_ROMDATA_dintern_9ro\ : std_logic;
signal \gpuOut_c_9\ : std_logic;
signal \D9_in_c\ : std_logic;
signal \CONTROL.N_170_cascade_\ : std_logic;
signal \N_186\ : std_logic;
signal \CONTROL.N_202\ : std_logic;
signal \N_186_cascade_\ : std_logic;
signal bus_9 : std_logic;
signal \CONTROL.ctrlOut_9\ : std_logic;
signal \INVCONTROL.dout_9C_net\ : std_logic;
signal \PROM.ROMDATA.m284\ : std_logic;
signal \PROM.ROMDATA.dintern_12dfltZ0Z_0\ : std_logic;
signal \PROM.ROMDATA.m284_cascade_\ : std_logic;
signal \controlWord_12_cascade_\ : std_logic;
signal \CONTROL.increment28lto5_0\ : std_logic;
signal \PROM.ROMDATA.m273\ : std_logic;
signal \PROM.ROMDATA.m273_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_11ro_cascade_\ : std_logic;
signal \CONTROL.increment28lto5_0_xZ0Z1\ : std_logic;
signal \CONTROL.increment28lto5_0_xZ0Z0\ : std_logic;
signal \PROM_ROMDATA_dintern_11ro\ : std_logic;
signal \aluStatus_4\ : std_logic;
signal \controlWord_12\ : std_logic;
signal \CONTROL.g0_1_i_a6Z0Z_0\ : std_logic;
signal \CONTROL.g0_1_i_a6Z0Z_1\ : std_logic;
signal \CONTROL.g0_3_i_a7Z0Z_0\ : std_logic;
signal \PROM.ROMDATA.m271_1\ : std_logic;
signal \PROM.ROMDATA.m271_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m258_ns\ : std_logic;
signal \PROM.ROMDATA.m258_ns_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_9ro_cascade_\ : std_logic;
signal \CONTROL.increment28lto5_1Z0Z_0\ : std_logic;
signal \PROM.ROMDATA.N_566_mux\ : std_logic;
signal \PROM.ROMDATA.m470_bm\ : std_logic;
signal \CONTROL.N_215\ : std_logic;
signal \CONTROL.N_86_0_cascade_\ : std_logic;
signal \controlWord_1\ : std_logic;
signal \CONTROL.N_135\ : std_logic;
signal \CONTROL.N_74_0\ : std_logic;
signal \CONTROL.N_249\ : std_logic;
signal \controlWord_5\ : std_logic;
signal \CONTROL.N_74_0_cascade_\ : std_logic;
signal \controlWord_6\ : std_logic;
signal \CONTROL.un1_busState96_1_i_i_232_1_cascade_\ : std_logic;
signal \CONTROL.programCounter_ret_36_RNINU4NARZ0Z_7\ : std_logic;
signal \PROM.ROMDATA.m23_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_31_0__N_556_mux\ : std_logic;
signal \PROM.ROMDATA.m294_am\ : std_logic;
signal \PROM.ROMDATA.m31\ : std_logic;
signal \m125_e_cascade_\ : std_logic;
signal \PROM.ROMDATA.N_557_mux\ : std_logic;
signal \PROM.ROMDATA.m77\ : std_logic;
signal m93_ns : std_logic;
signal \m93_ns_cascade_\ : std_logic;
signal \CONTROL.addrstack_5\ : std_logic;
signal \CONTROL.addrstack_reto_5\ : std_logic;
signal \CONTROL.programCounter_1_5\ : std_logic;
signal \CONTROL.programCounter_1_reto_5\ : std_logic;
signal \CONTROL.un1_programCounter9_reto_rep1\ : std_logic;
signal \CONTROL.g0_2Z0Z_1\ : std_logic;
signal \CONTROL.N_133_0_0\ : std_logic;
signal \CONTROL.N_114_i\ : std_logic;
signal \CONTROL.g1_1_4\ : std_logic;
signal \CONTROL.un1_busState114_2_0_0\ : std_logic;
signal \CONTROL.g1_1_cascade_\ : std_logic;
signal \CONTROL.addrstackptr_N_7_i\ : std_logic;
signal \CONTROL.g1_0_0\ : std_logic;
signal \CONTROL.g0_i_m2_1\ : std_logic;
signal \CONTROL.addrstack_1_7\ : std_logic;
signal \CONTROL.g0_4Z0Z_2\ : std_logic;
signal \CONTROL.g0_i_m2_1_cascade_\ : std_logic;
signal \CONTROL.g1_1\ : std_logic;
signal \CONTROL.addrstackptrZ0Z_7\ : std_logic;
signal \INVCONTROL.increment_0C_net\ : std_logic;
signal \PROM_ROMDATA_dintern_5ro\ : std_logic;
signal \CONTROL.g0_2_iZ0Z_1\ : std_logic;
signal \PROM.ROMDATA.m381_am\ : std_logic;
signal \PROM.ROMDATA.m375_am\ : std_logic;
signal \PROM.ROMDATA.m382_ns_1\ : std_logic;
signal \ALU.rshift_3_ns_1_0\ : std_logic;
signal \ALU.N_858_cascade_\ : std_logic;
signal \ALU.rshift_15_ns_1_0_cascade_\ : std_logic;
signal \ALU.rshift_3_ns_1_4_cascade_\ : std_logic;
signal \ALU.N_862\ : std_logic;
signal \ALU.N_862_cascade_\ : std_logic;
signal \ALU.N_922_cascade_\ : std_logic;
signal \ALU.d_RNIR6J013Z0Z_2\ : std_logic;
signal \ALU.d_RNI1AHUF8Z0Z_2\ : std_logic;
signal \ALU.mult_25_10\ : std_logic;
signal \ALU.mult_11_10\ : std_logic;
signal \ALU.mult_293_c_RNIOCJMDZ0Z9\ : std_logic;
signal \bfn_19_9_0_\ : std_logic;
signal \ALU.mult_11_11\ : std_logic;
signal \ALU.mult_21_11\ : std_logic;
signal \ALU.mult_21_c10\ : std_logic;
signal \ALU.mult_21_12\ : std_logic;
signal \ALU.mult_21_c11\ : std_logic;
signal \ALU.mult_21_13\ : std_logic;
signal \ALU.mult_21_c12\ : std_logic;
signal \ALU.mult_21_14\ : std_logic;
signal \ALU.mult_21_c13\ : std_logic;
signal \ALU.mult_23_15\ : std_logic;
signal \ALU.mult_21_c14\ : std_logic;
signal \ALU.mult_476_c_RNIFLP0OZ0Z7\ : std_logic;
signal \ALU.N_836\ : std_logic;
signal \ALU.mult_293_c_RNOZ0\ : std_logic;
signal \bfn_19_10_0_\ : std_logic;
signal \ALU.d_RNI34ECOZ0Z_9\ : std_logic;
signal \ALU.d_RNI0PI3E1Z0Z_8\ : std_logic;
signal \ALU.mult_9_10\ : std_logic;
signal \ALU.mult_9_c9\ : std_logic;
signal \ALU.d_RNIFCNKLZ0Z_9\ : std_logic;
signal \ALU.d_RNIDR5C61Z0Z_8\ : std_logic;
signal \ALU.mult_9_11\ : std_logic;
signal \ALU.mult_9_c10\ : std_logic;
signal \ALU.d_RNIG61LGZ0Z_9\ : std_logic;
signal \ALU.mult_9_12\ : std_logic;
signal \ALU.mult_9_c11\ : std_logic;
signal \ALU.d_RNI68LSHZ0Z_9\ : std_logic;
signal \ALU.mult_9_13\ : std_logic;
signal \ALU.mult_9_c12\ : std_logic;
signal \ALU.d_RNISSV4IZ0Z_9\ : std_logic;
signal \ALU.d_RNI371041Z0Z_8\ : std_logic;
signal \ALU.mult_9_14\ : std_logic;
signal \ALU.mult_9_c13\ : std_logic;
signal \ALU.c_RNI0QV651Z0Z_10\ : std_logic;
signal \ALU.mult_9_c14\ : std_logic;
signal \ALU.mult_323_c_RNIAA0BZ0Z82\ : std_logic;
signal \ALU.d_RNIGD2441Z0Z_8\ : std_logic;
signal \ALU.N_639_cascade_\ : std_logic;
signal \ALU.d_RNIC6EBM2Z0Z_2\ : std_logic;
signal \ALU.d_RNIFVCT15Z0Z_8_cascade_\ : std_logic;
signal \ALU.lshift_11\ : std_logic;
signal \ALU.N_851\ : std_logic;
signal \ALU.N_851_cascade_\ : std_logic;
signal \ALU.c_RNINT9PO2_0Z0Z_10\ : std_logic;
signal \ALU.N_978\ : std_logic;
signal \ALU.N_978_cascade_\ : std_logic;
signal \ALU.addsub_axb_1_1\ : std_logic;
signal \ALU.N_1026\ : std_logic;
signal \ALU.mult_293_c_RNOZ0Z_0\ : std_logic;
signal \ALU.N_1011\ : std_logic;
signal \ALU.N_852_cascade_\ : std_logic;
signal \ALU.N_966\ : std_logic;
signal \ALU.N_766_cascade_\ : std_logic;
signal \ALU.N_634\ : std_logic;
signal \ALU.N_634_cascade_\ : std_logic;
signal \ALU.N_811_cascade_\ : std_logic;
signal \ALU.d_RNIK8M6K5Z0Z_6\ : std_logic;
signal \ALU.a_15_sZ0Z_11\ : std_logic;
signal \ALU.d_RNIK8M6K5Z0Z_6_cascade_\ : std_logic;
signal \ALU.mult_489_c_RNI1J3GCUZ0\ : std_logic;
signal \ALU.aZ0Z_6\ : std_logic;
signal \ALU.N_766\ : std_logic;
signal \ALU.N_606_cascade_\ : std_logic;
signal \ALU.N_606\ : std_logic;
signal \ALU.N_638\ : std_logic;
signal \ALU.a_15_m0_amZ0Z_2\ : std_logic;
signal \ALU.a_15_m1_9_cascade_\ : std_logic;
signal \ALU.aZ0Z_9\ : std_logic;
signal \N_227_0\ : std_logic;
signal \N_179\ : std_logic;
signal bus_2 : std_logic;
signal \ALU.bZ0Z_4\ : std_logic;
signal \ALU.b_RNI5FSPZ0Z_4\ : std_logic;
signal \ALU.c_RNIHV2SZ0Z_9\ : std_logic;
signal h_4 : std_logic;
signal \ALU.dZ0Z_4\ : std_logic;
signal \ALU.d_RNI9R8EZ0Z_4\ : std_logic;
signal \aluOperand2_2\ : std_logic;
signal \ALU.N_1252_cascade_\ : std_logic;
signal \ALU.N_1204\ : std_logic;
signal \ALU.d_RNIO5IF4Z0Z_7_cascade_\ : std_logic;
signal \ALU.combOperand2_d_bmZ0Z_7\ : std_logic;
signal \ALU.d_RNIM3JB6Z0Z_7_cascade_\ : std_logic;
signal \ALU.dout_3_ns_1_7_cascade_\ : std_logic;
signal \ALU.operand2_6_ns_1_7\ : std_logic;
signal \aluOperand2_2_rep1\ : std_logic;
signal \ALU.operand2_3_ns_1_7\ : std_logic;
signal \aluOperand1_1_rep1\ : std_logic;
signal h_7 : std_logic;
signal \ALU.dout_6_ns_1_7_cascade_\ : std_logic;
signal \ALU.N_1140_cascade_\ : std_logic;
signal \ALU.N_1092\ : std_logic;
signal \DROM_ROMDATA_dintern_7ro\ : std_logic;
signal \aluOut_7_cascade_\ : std_logic;
signal \N_200\ : std_logic;
signal \PROM.ROMDATA.m267_cascade_\ : std_logic;
signal \PROM.ROMDATA.m442\ : std_logic;
signal \PROM.ROMDATA.m282\ : std_logic;
signal \PROM.ROMDATA.dintern_29dfltZ0Z_1\ : std_logic;
signal \PROM.ROMDATA.m282_cascade_\ : std_logic;
signal \CONTROL.ctrlOut_13\ : std_logic;
signal \INVCONTROL.dout_13C_net\ : std_logic;
signal \CONTROL.N_35\ : std_logic;
signal \PROM.ROMDATA.m444_am\ : std_logic;
signal \PROM.ROMDATA.m444_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m289\ : std_logic;
signal \PROM.ROMDATA.m418_ns_1\ : std_logic;
signal \PROM_ROMDATA_dintern_19ro\ : std_logic;
signal \PROM_ROMDATA_dintern_19ro_cascade_\ : std_logic;
signal \controlWord_19\ : std_logic;
signal f_3 : std_logic;
signal \controlWord_19_cascade_\ : std_logic;
signal \controlWord_20\ : std_logic;
signal f_4 : std_logic;
signal \A14_c\ : std_logic;
signal \A4_c\ : std_logic;
signal \A3_c\ : std_logic;
signal \RAM.un1_WR_105_0Z0Z_7\ : std_logic;
signal \controlWord_31\ : std_logic;
signal \A15_c\ : std_logic;
signal \INVCONTROL.ramAddReg_3C_net\ : std_logic;
signal \PROM.ROMDATA.m266\ : std_logic;
signal \PROM.ROMDATA.m157_cascade_\ : std_logic;
signal \PROM.ROMDATA.m265_cascade_\ : std_logic;
signal \PROM.ROMDATA.m268\ : std_logic;
signal \PROM.ROMDATA.m270_bm\ : std_logic;
signal \CONTROL.aluOperation_12_i_0_6\ : std_logic;
signal \controlWord_3\ : std_logic;
signal \CONTROL.N_219\ : std_logic;
signal \controlWord_2\ : std_logic;
signal \INVCONTROL.aluOperation_6C_net\ : std_logic;
signal \PROM.ROMDATA.N_544_mux\ : std_logic;
signal \PROM.ROMDATA.m258_bm\ : std_logic;
signal \CONTROL.programCounter_1_1\ : std_logic;
signal \CONTROL.programCounter_ret_19_RNIT3IGZ0Z_5\ : std_logic;
signal \CONTROL.programCounter_ret_1_RNI4MHFZ0Z_5\ : std_logic;
signal \CONTROL.un1_programCounter9_reto\ : std_logic;
signal \progRomAddress_5_cascade_\ : std_logic;
signal \PROM.ROMDATA.m243_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m244_ns_1_1\ : std_logic;
signal \CONTROL.ctrlOut_0\ : std_logic;
signal \PROM.ROMDATA.m243_1\ : std_logic;
signal \PROM.ROMDATA.m260_1\ : std_logic;
signal \N_417_cascade_\ : std_logic;
signal \CONTROL.programCounter_1_2\ : std_logic;
signal \CONTROL.programCounter_ret_1_RNI6OHFZ0Z_6\ : std_logic;
signal \CONTROL.ctrlOut_3\ : std_logic;
signal \CONTROL.programCounter_1_4\ : std_logic;
signal \PROM.ROMDATA.m215_ns_1_N_2L1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m215_ns_1\ : std_logic;
signal \CONTROL.g0_3_i_a7_0_0\ : std_logic;
signal \CONTROL.addrstack_2\ : std_logic;
signal \PROM.ROMDATA.m36\ : std_logic;
signal \PROM.ROMDATA.N_526_mux_cascade_\ : std_logic;
signal \PROM.ROMDATA.m238_bm\ : std_logic;
signal \aluStatus_i_3\ : std_logic;
signal \PROM_ROMDATA_dintern_10ro\ : std_logic;
signal \CONTROL.g0_5Z0Z_0\ : std_logic;
signal \PROM.ROMDATA.m258_am\ : std_logic;
signal \PROM_ROMDATA_dintern_31_0__N_555_mux\ : std_logic;
signal \CONTROL.ctrlOut_5\ : std_logic;
signal \CONTROL.dout_reto_5\ : std_logic;
signal \CONTROL.programCounter_ret_19_RNIV5IGZ0Z_6\ : std_logic;
signal \CONTROL.addrstack_6\ : std_logic;
signal \CONTROL.addrstack_reto_6\ : std_logic;
signal \PROM.ROMDATA.m48\ : std_logic;
signal \CONTROL.ctrlOut_6\ : std_logic;
signal \CONTROL.dout_reto_6\ : std_logic;
signal \PROM.ROMDATA.m7\ : std_logic;
signal \PROM.ROMDATA.m392_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m392_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m134\ : std_logic;
signal \PROM.ROMDATA.m396_bm\ : std_logic;
signal \PROM.ROMDATA.m396_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m396_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m401_ns_1\ : std_logic;
signal \PROM.ROMDATA.m401_ns\ : std_logic;
signal \ALU.N_607\ : std_logic;
signal \ALU.N_767\ : std_logic;
signal \ALU.N_607_cascade_\ : std_logic;
signal \ALU.lshift_3_ns_1_11\ : std_logic;
signal \ALU.d_RNI4N3K21Z0Z_8\ : std_logic;
signal \ALU.d_RNIH8D821Z0Z_8\ : std_logic;
signal \ALU.mult_335_c_RNOZ0\ : std_logic;
signal \bfn_20_10_0_\ : std_logic;
signal \ALU.c_RNIBQSTOZ0Z_11\ : std_logic;
signal \ALU.c_RNIG5G6F1Z0Z_10\ : std_logic;
signal \ALU.mult_11_12\ : std_logic;
signal \ALU.mult_11_c11\ : std_logic;
signal \ALU.c_RNIN266MZ0Z_11\ : std_logic;
signal \ALU.c_RNIT73F71Z0Z_10\ : std_logic;
signal \ALU.mult_11_13\ : std_logic;
signal \ALU.mult_11_c12\ : std_logic;
signal \ALU.c_RNIK31N31Z0Z_10\ : std_logic;
signal \ALU.mult_11_14\ : std_logic;
signal \ALU.mult_11_c13\ : std_logic;
signal \ALU.mult_11_c14\ : std_logic;
signal \ALU.mult_11_c14_THRU_CO\ : std_logic;
signal \ALU.c_RNIOSF6HZ0Z_11\ : std_logic;
signal \ALU.mult_335_c_RNOZ0Z_0\ : std_logic;
signal \ALU.N_835_cascade_\ : std_logic;
signal \ALU.N_852\ : std_logic;
signal \ALU.rshift_7_ns_1_7_cascade_\ : std_logic;
signal \ALU.N_925_cascade_\ : std_logic;
signal \ALU.N_833\ : std_logic;
signal \ALU.N_837\ : std_logic;
signal \ALU.rshift_7_ns_1_3_cascade_\ : std_logic;
signal \ALU.N_921\ : std_logic;
signal bus_7 : std_logic;
signal \ALU.N_1030\ : std_logic;
signal \ALU.c_RNI08R632Z0Z_15\ : std_logic;
signal \ALU.eZ0Z_1\ : std_logic;
signal \ALU.eZ0Z_0\ : std_logic;
signal \ALU.eZ0Z_7\ : std_logic;
signal \ALU.eZ0Z_8\ : std_logic;
signal \ALU.eZ0Z_15\ : std_logic;
signal \ALU.eZ0Z_9\ : std_logic;
signal \ALU.N_647\ : std_logic;
signal \ALU.N_643\ : std_logic;
signal \ALU.N_707\ : std_logic;
signal \ALU.addsub_cry_14_c_RNI134CV5Z0Z_0_cascade_\ : std_logic;
signal \ALU.addsub_cry_14_c_RNIKS9S5HZ0_cascade_\ : std_logic;
signal \ALU.c_RNIE4B6N4Z0Z_15\ : std_logic;
signal \ALU.a_15_1_15_cascade_\ : std_logic;
signal \ALU.aZ0Z_15\ : std_logic;
signal \ALU.N_812\ : std_logic;
signal \ALU.N_812_cascade_\ : std_logic;
signal \ALU.addsub_cry_14_c_RNI134CVZ0Z5\ : std_logic;
signal \ALU.N_635\ : std_logic;
signal \ALU.N_639\ : std_logic;
signal \ALU.cZ0Z_1\ : std_logic;
signal \ALU.cZ0Z_0\ : std_logic;
signal \ALU.cZ0Z_7\ : std_logic;
signal \ALU.cZ0Z_8\ : std_logic;
signal \ALU.cZ0Z_15\ : std_logic;
signal \ALU.cZ0Z_9\ : std_logic;
signal \ALU.log_1_7_cascade_\ : std_logic;
signal \ALU.mult_7\ : std_logic;
signal \ALU.mult_492_c_RNIQ5BZ0Z457_cascade_\ : std_logic;
signal \ALU.lshift_7\ : std_logic;
signal \ALU.mult_492_c_RNIGN2JECZ0_cascade_\ : std_logic;
signal \ALU.aZ0Z_7\ : std_logic;
signal \ALU.d_RNIO75BGZ0Z_7\ : std_logic;
signal \aluOperand2_2_rep2\ : std_logic;
signal \ALU.c_RNI9SHFZ0Z_14\ : std_logic;
signal \ALU.a_RNI5CPUZ0Z_14_cascade_\ : std_logic;
signal \aluOperand2_1\ : std_logic;
signal \ALU.d_RNICJCTZ0Z_14\ : std_logic;
signal \ALU.operand2_7_ns_1_14_cascade_\ : std_logic;
signal \ALU.b_RNI83KC1Z0Z_14\ : std_logic;
signal \N_191\ : std_logic;
signal \ALU.operand2_14_cascade_\ : std_logic;
signal \ALU.d_RNINISC7Z0Z_14\ : std_logic;
signal \ALU.dout_3_ns_1_14_cascade_\ : std_logic;
signal \aluOperand1_2\ : std_logic;
signal \ALU.dout_6_ns_1_14_cascade_\ : std_logic;
signal \aluOperand1_1\ : std_logic;
signal \ALU.N_1099\ : std_logic;
signal \ALU.N_1147_cascade_\ : std_logic;
signal \DROM_ROMDATA_dintern_14ro\ : std_logic;
signal \aluOut_14_cascade_\ : std_logic;
signal \N_207\ : std_logic;
signal \CONTROL.un1_busState114_2_0_o2_0_0\ : std_logic;
signal \CONTROL.N_361_1\ : std_logic;
signal \CONTROL.un1_busState114_2_0_0_0\ : std_logic;
signal \INVCONTROL.increment_1C_net\ : std_logic;
signal \PROM.ROMDATA.m422_am\ : std_logic;
signal \PROM.ROMDATA.m422_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m381_bm\ : std_logic;
signal \PROM.ROMDATA.m298_am\ : std_logic;
signal \CONTROL.programCounter_1_axb_4\ : std_logic;
signal \PROM.ROMDATA.N_543_mux_2_cascade_\ : std_logic;
signal \PROM.ROMDATA.N_559_mux\ : std_logic;
signal \PROM.ROMDATA.m392_am\ : std_logic;
signal \PROM.ROMDATA.m163_cascade_\ : std_logic;
signal \PROM.ROMDATA.m176_x\ : std_logic;
signal \PROM.ROMDATA.N_543_mux_2\ : std_logic;
signal \PROM.ROMDATA.N_569_mux\ : std_logic;
signal \PROM.ROMDATA.m109_am_1_cascade_\ : std_logic;
signal \CONTROL.addrstack_0\ : std_logic;
signal \N_415\ : std_logic;
signal \N_419\ : std_logic;
signal \CONTROL.addrstackZ0Z_1\ : std_logic;
signal \CONTROL.dout_reto_3\ : std_logic;
signal \CONTROL.programCounter_ret_1_RNILA8IZ0Z_3_cascade_\ : std_logic;
signal \CONTROL.programCounter_ret_19_RNIEO8JZ0Z_3\ : std_logic;
signal \CONTROL.programCounter_1_reto_0\ : std_logic;
signal \CONTROL.addrstack_3\ : std_logic;
signal \PROM.ROMDATA.m30\ : std_logic;
signal \PROM.ROMDATA.m35_1\ : std_logic;
signal \PROM.ROMDATA.m35\ : std_logic;
signal \CONTROL.programCounter_1_reto_2\ : std_logic;
signal \PROM.ROMDATA.m215_ns_1_1_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m215_ns_1_1\ : std_logic;
signal \PROM.ROMDATA.m256\ : std_logic;
signal \PROM.ROMDATA.m38\ : std_logic;
signal \PROM.ROMDATA.m251\ : std_logic;
signal \PROM.ROMDATA.m253\ : std_logic;
signal \CONTROL.programCounter_1_6\ : std_logic;
signal \CONTROL.programCounter_1_reto_6\ : std_logic;
signal \PROM.ROMDATA.m51\ : std_logic;
signal \PROM.ROMDATA.m433_am\ : std_logic;
signal \PROM.ROMDATA.m399_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m399_bm\ : std_logic;
signal \PROM.ROMDATA.m399_ns\ : std_logic;
signal \PROM.ROMDATA.m461_ns_1\ : std_logic;
signal \CONTROL.addrstack_4\ : std_logic;
signal \PROM.ROMDATA.m22\ : std_logic;
signal \PROM.ROMDATA.m451_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m451_am\ : std_logic;
signal \PROM.ROMDATA.m451_ns\ : std_logic;
signal \PROM.ROMDATA.m375_bm\ : std_logic;
signal \PROM.ROMDATA.m376\ : std_logic;
signal \PROM.ROMDATA.N_256_i\ : std_logic;
signal \PROM.ROMDATA.m389_bm\ : std_logic;
signal \PROM.ROMDATA.m389_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m389_ns\ : std_logic;
signal \ALU.lshift_3_ns_1_13_cascade_\ : std_logic;
signal \ALU.N_645_cascade_\ : std_logic;
signal \ALU.N_806_1\ : std_logic;
signal \ALU.a_15_m1_am_1_13_cascade_\ : std_logic;
signal \ALU.N_611_cascade_\ : std_logic;
signal \ALU.N_609\ : std_logic;
signal \ALU.N_641\ : std_logic;
signal \ALU.N_641_cascade_\ : std_logic;
signal \ALU.N_637\ : std_logic;
signal \ALU.d_RNITG2137Z0Z_0\ : std_logic;
signal \ALU.N_765\ : std_logic;
signal \ALU.a_15_m1_am_1_9\ : std_logic;
signal \ALU.a_15_m3_d_d_0_ns_1_3\ : std_logic;
signal \ALU.d_RNILTVJG3Z0Z_3\ : std_logic;
signal \ALU.mult_555_c_RNIJF56AMZ0_cascade_\ : std_logic;
signal \ALU.aZ0Z_12\ : std_logic;
signal \ALU.N_612\ : std_logic;
signal \ALU.N_614\ : std_logic;
signal \ALU.lshift_7_ns_1_12_cascade_\ : std_logic;
signal \ALU.N_704_cascade_\ : std_logic;
signal \ALU.d_RNIGNBT49Z0Z_8\ : std_logic;
signal \ALU.d_RNIGNBT49Z0Z_8_cascade_\ : std_logic;
signal \ALU.N_18_0\ : std_logic;
signal h_8 : std_logic;
signal \ALU.mult_12\ : std_logic;
signal \ALU.mult_555_c_RNI5VJUOIZ0\ : std_logic;
signal \ALU.mult_546_c_RNIG1E6IZ0Z8\ : std_logic;
signal \aluStatus_0\ : std_logic;
signal \ALU.status_14_12_0_cascade_\ : std_logic;
signal \ALU.status_RNO_1Z0Z_0\ : std_logic;
signal \ALU.bZ0Z_1\ : std_logic;
signal \ALU.bZ0Z_0\ : std_logic;
signal \ALU.bZ0Z_7\ : std_logic;
signal \ALU.bZ0Z_8\ : std_logic;
signal \ALU.bZ0Z_9\ : std_logic;
signal \ALU.mult_9_8\ : std_logic;
signal \ALU.mult_25_8\ : std_logic;
signal \ALU.mult_495_c_RNIKOB51JZ0_cascade_\ : std_logic;
signal \ALU.aZ0Z_8\ : std_logic;
signal \ALU.lshift_15_ns_1_8\ : std_logic;
signal \ALU.N_610\ : std_logic;
signal \ALU.N_608\ : std_logic;
signal \ALU.N_640\ : std_logic;
signal \ALU.addsub_cry_7_c_RNIDLTNZ0Z71_cascade_\ : std_logic;
signal \ALU.lshift_8\ : std_logic;
signal \ALU.N_636\ : std_logic;
signal \ALU.N_794_1\ : std_logic;
signal \ALU.N_809\ : std_logic;
signal f_1 : std_logic;
signal f_0 : std_logic;
signal f_7 : std_logic;
signal f_8 : std_logic;
signal f_9 : std_logic;
signal g_1 : std_logic;
signal g_0 : std_logic;
signal g_7 : std_logic;
signal g_8 : std_logic;
signal g_15 : std_logic;
signal \ALU.c_RNID85GQ_0Z0Z_15_cascade_\ : std_logic;
signal \ALU.c_RNI9DCRE2Z0Z_15\ : std_logic;
signal \DROM_ROMDATA_dintern_adflt\ : std_logic;
signal \DROM_ROMDATA_dintern_15ro\ : std_logic;
signal \busState_1\ : std_logic;
signal \N_208_cascade_\ : std_logic;
signal \ALU.status_19_14_cascade_\ : std_logic;
signal \N_208\ : std_logic;
signal \busState_0\ : std_logic;
signal \CONTROL.bus_7_ns_1_15\ : std_logic;
signal \busState_2\ : std_logic;
signal bus_15 : std_logic;
signal \ALU.a_15_m2_d_d_sZ0Z_0\ : std_logic;
signal \bus_15_cascade_\ : std_logic;
signal \ALU.c_RNIJI6SHZ0Z_15\ : std_logic;
signal \ALU.c_RNID85GQZ0Z_15\ : std_logic;
signal \PROM.ROMDATA.m248_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m249\ : std_logic;
signal \PROM.ROMDATA.m359\ : std_logic;
signal \PROM.ROMDATA.m150_cascade_\ : std_logic;
signal \PROM.ROMDATA.m228_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m25\ : std_logic;
signal \PROM.ROMDATA.m280\ : std_logic;
signal \PROM.ROMDATA.m438\ : std_logic;
signal \PROM.ROMDATA.m173\ : std_logic;
signal \PROM.ROMDATA.m23\ : std_logic;
signal \PROM_ROMDATA_dintern_31_0__g1\ : std_logic;
signal \PROM.ROMDATA.m169_cascade_\ : std_logic;
signal \PROM.ROMDATA.m270_am\ : std_logic;
signal \PROM.ROMDATA.m13_cascade_\ : std_logic;
signal \PROM.ROMDATA.m188\ : std_logic;
signal \PROM.ROMDATA.m13\ : std_logic;
signal \PROM.ROMDATA.m263\ : std_logic;
signal \CONTROL.ctrlOut_1\ : std_logic;
signal \CONTROL.dout_reto_0\ : std_logic;
signal \CONTROL_addrstack_reto_0\ : std_logic;
signal \PROM.ROMDATA.m248_ns_1\ : std_logic;
signal \CONTROL.incrementZ0Z_0\ : std_logic;
signal \CONTROL.incrementZ0Z_1\ : std_logic;
signal \PROM.ROMDATA.m284_1\ : std_logic;
signal \CONTROL.programCounter_ret_19_RNI8I8JZ0Z_0\ : std_logic;
signal \CONTROL.programCounter_ret_1_RNIF48IZ0Z_0\ : std_logic;
signal \progRomAddress_0_cascade_\ : std_logic;
signal \PROM.ROMDATA.m72_cascade_\ : std_logic;
signal \PROM.ROMDATA.m74\ : std_logic;
signal \PROM.ROMDATA.m80_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m93_ns_1\ : std_logic;
signal \CONTROL.programCounter_ret_1_RNIJ88IZ0Z_2\ : std_logic;
signal \CONTROL.programCounter_ret_19_RNICM8JZ0Z_2\ : std_logic;
signal \progRomAddress_2_cascade_\ : std_logic;
signal \PROM.ROMDATA.m195_am\ : std_logic;
signal \PROM.ROMDATA.m196_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m179\ : std_logic;
signal \PROM.ROMDATA.m185_am\ : std_logic;
signal \PROM.ROMDATA.m191_cascade_\ : std_logic;
signal \PROM.ROMDATA.m193\ : std_logic;
signal \PROM.ROMDATA.m195_bm\ : std_logic;
signal \CONTROL.programCounter_1_3\ : std_logic;
signal \CONTROL.programCounter_1_reto_3\ : std_logic;
signal \PROM.ROMDATA.m92_am\ : std_logic;
signal \PROM.ROMDATA.m62_cascade_\ : std_logic;
signal \PROM.ROMDATA.m53_am\ : std_logic;
signal \PROM.ROMDATA.m53_bm\ : std_logic;
signal \PROM.ROMDATA.m64_bm\ : std_logic;
signal \PROM.ROMDATA.m65_ns_1_cascade_\ : std_logic;
signal m65_ns : std_logic;
signal \PROM.ROMDATA.m58_cascade_\ : std_logic;
signal \PROM.ROMDATA.m64_am\ : std_logic;
signal \PROM.ROMDATA.m45\ : std_logic;
signal \ALU.log_1_7\ : std_logic;
signal \ALU.log_1_5\ : std_logic;
signal \ALU.log_1_11\ : std_logic;
signal \ALU.log_1_10\ : std_logic;
signal \ALU.N_22_0\ : std_logic;
signal \ALU.N_20_0\ : std_logic;
signal \ALU.status_8_10_0_cascade_\ : std_logic;
signal \ALU.status_8_13_0\ : std_logic;
signal \ALU.status_8_3_1_0\ : std_logic;
signal \ALU.log_1_15_cascade_\ : std_logic;
signal \ALU.status_8_13_1_0\ : std_logic;
signal \ALU.c_RNIV5AOKZ0Z_13_cascade_\ : std_logic;
signal \ALU.c_RNIO5N04A_0Z0Z_13_cascade_\ : std_logic;
signal \ALU.bZ0Z_13\ : std_logic;
signal \ALU.c_RNIV5AOKZ0Z_13\ : std_logic;
signal \ALU.d_RNIRFBHE9Z0Z_0\ : std_logic;
signal \ALU.log_1_4\ : std_logic;
signal \ALU.N_16_0_cascade_\ : std_logic;
signal \ALU.status_8_8_0\ : std_logic;
signal \ALU.log_1_9\ : std_logic;
signal \ALU.d_RNI7KS2IZ0Z_9\ : std_logic;
signal \ALU.eZ0Z_12\ : std_logic;
signal \ALU.eZ0Z_13\ : std_logic;
signal \ALU.eZ0Z_14\ : std_logic;
signal g_12 : std_logic;
signal g_13 : std_logic;
signal g_14 : std_logic;
signal \ALU.a_15_ns_1_1\ : std_logic;
signal \ALU.dZ0Z_1\ : std_logic;
signal \ALU.d_RNINUGCF4Z0Z_0\ : std_logic;
signal \ALU.rshift_0\ : std_logic;
signal \ALU.dZ0Z_0\ : std_logic;
signal \ALU.a_15_m0_7\ : std_logic;
signal \ALU.mult_492_c_RNIGN2JECZ0\ : std_logic;
signal \ALU.dZ0Z_7\ : std_logic;
signal \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\ : std_logic;
signal \ALU.a_15_m3_sZ0Z_13\ : std_logic;
signal \ALU.mult_495_c_RNIKOB51JZ0\ : std_logic;
signal \ALU.dZ0Z_8\ : std_logic;
signal \ALU.mult_15\ : std_logic;
signal \ALU.a_15_1_15\ : std_logic;
signal \ALU.a_15_m1_9\ : std_logic;
signal \ALU.mult_546_c_RNIJOT4JZ0Z8\ : std_logic;
signal \ALU.dZ0Z_9\ : std_logic;
signal \ALU.N_835\ : std_logic;
signal \ALU.d_RNIPFFDD1_0Z0Z_6_cascade_\ : std_logic;
signal \ALU.N_863_cascade_\ : std_logic;
signal \ALU.d_RNIN3H0DZ0Z_3\ : std_logic;
signal \ALU.d_RNIGPBNB6Z0Z_2_cascade_\ : std_logic;
signal \ALU.a_15_m0_5\ : std_logic;
signal bus_5 : std_logic;
signal \ALU.c_RNINGV0T2Z0Z_15\ : std_logic;
signal \ALU.d_RNIPFFDD1Z0Z_6\ : std_logic;
signal \ALU.status_14_0_0_cascade_\ : std_logic;
signal \ALU.status_14_5_0\ : std_logic;
signal \ALU.status_14_7_0_cascade_\ : std_logic;
signal \ALU.status_14_13_0\ : std_logic;
signal \ALU.N_979\ : std_logic;
signal \ALU.N_979_cascade_\ : std_logic;
signal \ALU.combOperand2_a0_0Z0Z_6\ : std_logic;
signal \ALU.status_RNO_22Z0Z_0\ : std_logic;
signal \ALU.status_14_6_0\ : std_logic;
signal \ALU.status_17_I_21_c_RNOZ0\ : std_logic;
signal \ALU.status_e_0_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \ALU.N_570_cascade_\ : std_logic;
signal \ALU.status_e_0_RNO_1Z0Z_2\ : std_logic;
signal \aluStatus_2\ : std_logic;
signal \PROM_ROMDATA_dintern_9ro\ : std_logic;
signal \CONTROL.g3Z0Z_0\ : std_logic;
signal \ALU.bZ0Z_15\ : std_logic;
signal \aluOperand2_fast_2\ : std_logic;
signal f_15 : std_logic;
signal \aluOperand2_fast_1\ : std_logic;
signal \ALU.operand2_6_ns_1_15_cascade_\ : std_logic;
signal \aluOperand2_1_rep1\ : std_logic;
signal \ALU.dZ0Z_15\ : std_logic;
signal \ALU.dout_6_ns_1_15\ : std_logic;
signal \aluOperand1_1_rep2\ : std_logic;
signal h_15 : std_logic;
signal \ALU.N_1100\ : std_logic;
signal \ALU.N_1148_cascade_\ : std_logic;
signal \aluOperand1_0\ : std_logic;
signal \ALU.N_1260\ : std_logic;
signal \ALU.N_1212\ : std_logic;
signal \aluOperand2_0\ : std_logic;
signal \ALU.combOperand2_d_bmZ0Z_15\ : std_logic;
signal \ALU.c_RNI8VV95Z0Z_15_cascade_\ : std_logic;
signal \ALU.c_RNIJTKD7Z0Z_15\ : std_logic;
signal \PROM.ROMDATA.m320_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m410_am\ : std_logic;
signal \PROM.ROMDATA.m413_am_cascade_\ : std_logic;
signal \CONTROL.ctrlOut_2\ : std_logic;
signal \CONTROL.dout_reto_2\ : std_logic;
signal \CONTROL.N_136_0\ : std_logic;
signal \CONTROL.N_86_0\ : std_logic;
signal \CONTROL.N_98_0\ : std_logic;
signal \controlWord_4\ : std_logic;
signal \PROM.ROMDATA.m320_am\ : std_logic;
signal \PROM.ROMDATA.m150\ : std_logic;
signal \PROM.ROMDATA.N_558_mux\ : std_logic;
signal \PROM.ROMDATA.m49_cascade_\ : std_logic;
signal \PROM.ROMDATA.m229_1\ : std_logic;
signal \PROM.ROMDATA.m228_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m229\ : std_logic;
signal \PROM.ROMDATA.m437_ns\ : std_logic;
signal \PROM.ROMDATA.m312_bm\ : std_logic;
signal \PROM.ROMDATA.m312_am\ : std_logic;
signal \PROM.ROMDATA.m437_ns_1\ : std_logic;
signal \PROM.ROMDATA.m11_bm\ : std_logic;
signal \PROM.ROMDATA.m18_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m11_am\ : std_logic;
signal \PROM.ROMDATA.m19_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m18_am\ : std_logic;
signal \PROM.ROMDATA.m19_ns\ : std_logic;
signal \PROM.ROMDATA.m33\ : std_logic;
signal \CONTROL.dout_reto_1\ : std_logic;
signal \CONTROL.programCounter_1_reto_1\ : std_logic;
signal \CONTROL.programCounter_ret_1_RNIH68IZ0Z_1_cascade_\ : std_logic;
signal \CONTROL.programCounter_ret_19_RNIAK8JZ0Z_1\ : std_logic;
signal \progRomAddress_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m55\ : std_logic;
signal \CONTROL.programCounter_1_reto_4\ : std_logic;
signal \CONTROL_addrstack_reto_4\ : std_logic;
signal \CONTROL.programCounter11_reto_fast\ : std_logic;
signal \CONTROL.un1_programCounter9_reto_fast\ : std_logic;
signal \CONTROL.programCounter_ret_1_RNINC8IZ0Z_4_cascade_\ : std_logic;
signal \CONTROL.programCounter_ret_19_RNIGQ8JZ0Z_4\ : std_logic;
signal \PROM.ROMDATA.m143\ : std_logic;
signal \progRomAddress_4_cascade_\ : std_logic;
signal \PROM.ROMDATA.m145\ : std_logic;
signal \PROM.ROMDATA.m90\ : std_logic;
signal \PROM.ROMDATA.m92_bm\ : std_logic;
signal \PROM.ROMDATA.m183_cascade_\ : std_logic;
signal \PROM.ROMDATA.m185_bm\ : std_logic;
signal \PROM.ROMDATA.N_525_mux_cascade_\ : std_logic;
signal \PROM.ROMDATA.i4_mux\ : std_logic;
signal \PROM.ROMDATA.m103\ : std_logic;
signal \PROM.ROMDATA.m226\ : std_logic;
signal \PROM.ROMDATA.m92_am_1\ : std_logic;
signal \PROM.ROMDATA.m158\ : std_logic;
signal \PROM.ROMDATA.m158_cascade_\ : std_logic;
signal \PROM.ROMDATA.m196_ns\ : std_logic;
signal \PROM_ROMDATA_dintern_6ro\ : std_logic;
signal \CONTROL.ctrlOut_4\ : std_logic;
signal \CONTROL.dout_reto_4\ : std_logic;
signal \ALU.aluOut_i_0\ : std_logic;
signal \bfn_23_7_0_\ : std_logic;
signal \ALU.aluOut_i_1\ : std_logic;
signal \ALU.status_19_cry_0\ : std_logic;
signal \ALU.aluOut_i_2\ : std_logic;
signal \ALU.status_19_cry_1\ : std_logic;
signal \ALU.aluOut_i_3\ : std_logic;
signal \ALU.status_19_cry_2\ : std_logic;
signal \ALU.status_19_3\ : std_logic;
signal \ALU.aluOut_i_4\ : std_logic;
signal \ALU.status_19_cry_3\ : std_logic;
signal \ALU.status_19_4\ : std_logic;
signal \ALU.aluOut_i_5\ : std_logic;
signal \ALU.status_19_cry_4\ : std_logic;
signal \ALU.status_19_5\ : std_logic;
signal \ALU.aluOut_i_6\ : std_logic;
signal \ALU.status_19_cry_5\ : std_logic;
signal \ALU.status_19_6\ : std_logic;
signal \ALU.aluOut_i_7\ : std_logic;
signal \ALU.status_19_cry_6\ : std_logic;
signal \ALU.status_19_cry_7\ : std_logic;
signal \ALU.status_19_7\ : std_logic;
signal \ALU.aluOut_i_8\ : std_logic;
signal \bfn_23_8_0_\ : std_logic;
signal \ALU.status_19_8\ : std_logic;
signal \ALU.aluOut_i_9\ : std_logic;
signal \ALU.status_19_cry_8\ : std_logic;
signal \ALU.status_19_9\ : std_logic;
signal \ALU.aluOut_i_10\ : std_logic;
signal \ALU.status_19_cry_9\ : std_logic;
signal \ALU.status_19_10\ : std_logic;
signal \ALU.aluOut_i_11\ : std_logic;
signal \ALU.status_19_cry_10\ : std_logic;
signal \ALU.N_126\ : std_logic;
signal \ALU.aluOut_i_12\ : std_logic;
signal \ALU.status_19_cry_11\ : std_logic;
signal \ALU.N_125\ : std_logic;
signal \ALU.aluOut_i_13\ : std_logic;
signal \ALU.status_19_cry_12\ : std_logic;
signal \ALU.status_19_13\ : std_logic;
signal \ALU.aluOut_i_14\ : std_logic;
signal \ALU.status_19_cry_13\ : std_logic;
signal \ALU.aluOut_i_15\ : std_logic;
signal \ALU.status_19_cry_14\ : std_logic;
signal \ALU.status_19Z0Z_5\ : std_logic;
signal \bfn_23_9_0_\ : std_logic;
signal \aluStatus_5\ : std_logic;
signal \ALU.un1_a41_0\ : std_logic;
signal \ALU.aZ0Z32\ : std_logic;
signal \ALU.N_866\ : std_logic;
signal \ALU.N_967\ : std_logic;
signal \ALU.log_1_3\ : std_logic;
signal \ALU.lshift62_2\ : std_logic;
signal \ALU.mult_558_c_RNIB3E8DCZ0\ : std_logic;
signal \ALU.a_15_d_ns_1_13_cascade_\ : std_logic;
signal \ALU.mult_558_c_RNIB75F9GZ0_cascade_\ : std_logic;
signal \ALU.aZ0Z_13\ : std_logic;
signal \ALU.d_RNIJ7J1M5_0Z0Z_2\ : std_logic;
signal \ALU.a_15_m3_d_sZ0Z_8\ : std_logic;
signal bus_0_8 : std_logic;
signal \ALU.a_15_m3_d_sZ0Z_8_cascade_\ : std_logic;
signal \ALU.d_RNI12L8C5Z0Z_2\ : std_logic;
signal \ALU.d_RNIJ7J1M5Z0Z_2\ : std_logic;
signal f_12 : std_logic;
signal f_13 : std_logic;
signal f_14 : std_logic;
signal \ALU.log_1_14\ : std_logic;
signal \ALU.a_15_m0_14\ : std_logic;
signal \ALU.addsub_cry_13_c_RNIBVHEA1Z0Z_0_cascade_\ : std_logic;
signal \ALU.addsub_cry_13_c_RNIBVHEAZ0Z1\ : std_logic;
signal \ALU.addsub_cry_13_c_RNIJMTGAZ0Z5_cascade_\ : std_logic;
signal \ALU.mult_14\ : std_logic;
signal \ALU.a_15_ns_rn_0_14_cascade_\ : std_logic;
signal \ALU.aZ0Z_14\ : std_logic;
signal \ALU.a_15_sZ0Z_3\ : std_logic;
signal \ALU.a_15_m2_sZ0Z_15\ : std_logic;
signal \ALU.a_15_sm0\ : std_logic;
signal \aluOperation_1\ : std_logic;
signal \ALU.a_15_ns_1_7\ : std_logic;
signal \ALU.mult_388_c_RNIPGN6QZ0Z7\ : std_logic;
signal \ALU.rshift_3\ : std_logic;
signal \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\ : std_logic;
signal h_3 : std_logic;
signal \ALU.a_15_sZ0Z_13\ : std_logic;
signal \ALU.c_RNIO0KOKEZ0Z_10\ : std_logic;
signal \ALU.mult_549_c_RNIE7260OZ0\ : std_logic;
signal h_10 : std_logic;
signal \ALU.c_RNIBN2FN8Z0Z_11\ : std_logic;
signal \ALU.mult_552_c_RNIOT7VLFZ0Z_0\ : std_logic;
signal \ALU.mult_552_c_RNIOT7VLFZ0\ : std_logic;
signal h_11 : std_logic;
signal h_12 : std_logic;
signal h_13 : std_logic;
signal h_14 : std_logic;
signal \CONTROL.addrstack_1\ : std_logic;
signal \CONTROL.addrstackptrZ0Z_4\ : std_logic;
signal \CONTROL.addrstackptrZ0Z_2\ : std_logic;
signal \CONTROL.g1_1_3\ : std_logic;
signal \bfn_23_14_0_\ : std_logic;
signal \aluOut_0\ : std_logic;
signal \ALU.d_RNI27KBDZ0Z_0\ : std_logic;
signal \ALU.addsub_0\ : std_logic;
signal \ALU.addsub_cry_0_c_THRU_CO\ : std_logic;
signal \ALU.d_RNIIEOKOZ0Z_1\ : std_logic;
signal \ALU.addsub_1\ : std_logic;
signal \ALU.addsub_cry_0\ : std_logic;
signal \ALU.d_RNIN178LZ0Z_2\ : std_logic;
signal \ALU.addsub_2\ : std_logic;
signal \ALU.addsub_cry_1\ : std_logic;
signal \aluOut_3\ : std_logic;
signal \ALU.d_RNI04H8GZ0Z_3\ : std_logic;
signal \ALU.addsub_3\ : std_logic;
signal \ALU.addsub_cry_2\ : std_logic;
signal \aluOut_4\ : std_logic;
signal \ALU.d_RNI7BF7IZ0Z_4\ : std_logic;
signal \ALU.addsub_4\ : std_logic;
signal \ALU.addsub_cry_3\ : std_logic;
signal \aluOut_5\ : std_logic;
signal \ALU.d_RNI58QFIZ0Z_5\ : std_logic;
signal \ALU.addsub_5\ : std_logic;
signal \ALU.addsub_cry_4\ : std_logic;
signal \aluOut_6\ : std_logic;
signal \ALU.d_RNIALE3IZ0Z_6\ : std_logic;
signal \ALU.addsub_6\ : std_logic;
signal \ALU.addsub_cry_5\ : std_logic;
signal \ALU.addsub_cry_6\ : std_logic;
signal \aluOut_7\ : std_logic;
signal \ALU.d_RNI500DGZ0Z_7\ : std_logic;
signal \ALU.addsub_7\ : std_logic;
signal \bfn_23_15_0_\ : std_logic;
signal \aluOut_8\ : std_logic;
signal \ALU.d_RNIAJ1KHZ0Z_8\ : std_logic;
signal \ALU.addsub_8\ : std_logic;
signal \ALU.addsub_cry_7\ : std_logic;
signal \ALU.addsub_cry_8\ : std_logic;
signal \ALU.c_RNI1QK5KZ0Z_10\ : std_logic;
signal \aluOut_10\ : std_logic;
signal \ALU.addsub_10\ : std_logic;
signal \ALU.addsub_cry_9\ : std_logic;
signal \aluOut_11\ : std_logic;
signal \ALU.c_RNIRRB4IZ0Z_11\ : std_logic;
signal \ALU.addsub_11\ : std_logic;
signal \ALU.addsub_cry_10\ : std_logic;
signal \ALU.c_RNITVOEKZ0Z_12\ : std_logic;
signal \aluOut_12\ : std_logic;
signal \ALU.addsub_12\ : std_logic;
signal \ALU.addsub_cry_11\ : std_logic;
signal \ALU.c_RNIVHVMKZ0Z_13\ : std_logic;
signal \aluOut_13\ : std_logic;
signal \ALU.addsub_13\ : std_logic;
signal \ALU.addsub_cry_12\ : std_logic;
signal \ALU.c_RNIDDGOIZ0Z_14\ : std_logic;
signal \aluOut_14\ : std_logic;
signal \ALU.addsub_14\ : std_logic;
signal \ALU.addsub_cry_13\ : std_logic;
signal \ALU.addsub_cry_14\ : std_logic;
signal \ALU.c_RNI0NMSHZ0Z_15\ : std_logic;
signal \aluOut_15\ : std_logic;
signal \ALU.addsub_15\ : std_logic;
signal \bfn_23_16_0_\ : std_logic;
signal \aluStatus_1\ : std_logic;
signal \ALU.addsub_cry_15\ : std_logic;
signal \ALU.N_545\ : std_logic;
signal bus_6 : std_logic;
signal \ALU.c_RNIPBAG72Z0Z_14\ : std_logic;
signal \aluParams_0\ : std_logic;
signal \ALU.combOperand2_0_9\ : std_logic;
signal \aluOut_9\ : std_logic;
signal \ALU.d_RNI70I1IZ0Z_9\ : std_logic;
signal \ALU.N_980\ : std_logic;
signal \ALU.N_1029\ : std_logic;
signal \PROM.ROMDATA.m500_ns_1\ : std_logic;
signal \PROM.ROMDATA.m500_ns\ : std_logic;
signal \PROM.ROMDATA.m498_bm\ : std_logic;
signal \PROM.ROMDATA.m498_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m498_ns\ : std_logic;
signal \PROM.ROMDATA.m317_am\ : std_logic;
signal \PROM.ROMDATA.m317_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m312_ns\ : std_logic;
signal \PROM.ROMDATA.m317_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m325_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m320_ns\ : std_logic;
signal \PROM.ROMDATA.m325_ns\ : std_logic;
signal \PROM_ROMDATA_dintern_14ro_cascade_\ : std_logic;
signal \PROM.ROMDATA.m494_ns\ : std_logic;
signal \PROM.ROMDATA.m414_ns_1\ : std_logic;
signal \PROM.ROMDATA.m413_bm\ : std_logic;
signal \PROM.ROMDATA.m414_ns\ : std_logic;
signal \PROM.ROMDATA.m304\ : std_logic;
signal \PROM_ROMDATA_dintern_13ro_cascade_\ : std_logic;
signal \INVCONTROL.results_1C_net\ : std_logic;
signal \PROM.ROMDATA.m198\ : std_logic;
signal \PROM.ROMDATA.m16\ : std_logic;
signal \CONTROL.N_45_0\ : std_logic;
signal \PROM_ROMDATA_dintern_15ro_cascade_\ : std_logic;
signal \INVCONTROL.results_2C_net\ : std_logic;
signal \PROM.ROMDATA.m139\ : std_logic;
signal \PROM.ROMDATA.N_564_mux\ : std_logic;
signal \PROM.ROMDATA.m298_bm\ : std_logic;
signal \PROM.ROMDATA.N_72_i\ : std_logic;
signal \PROM.ROMDATA.N_565_mux\ : std_logic;
signal \PROM.ROMDATA.m287_cascade_\ : std_logic;
signal \PROM.ROMDATA.m410_bm\ : std_logic;
signal \PROM.ROMDATA.m66\ : std_logic;
signal \PROM.ROMDATA.m163\ : std_logic;
signal \PROM.ROMDATA.m490\ : std_logic;
signal \PROM.ROMDATA.m149\ : std_logic;
signal \PROM.ROMDATA.m118\ : std_logic;
signal \PROM.ROMDATA.m117\ : std_logic;
signal \PROM.ROMDATA.m157\ : std_logic;
signal \PROM.ROMDATA.m456_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m456_ns\ : std_logic;
signal \N_418\ : std_logic;
signal \CONTROL_addrstack_reto_3\ : std_logic;
signal \PROM.ROMDATA.m166_e\ : std_logic;
signal \PROM.ROMDATA.m104_ns_1\ : std_logic;
signal \PROM.ROMDATA.m107\ : std_logic;
signal \PROM.ROMDATA.m104_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m109_am\ : std_logic;
signal \PROM.ROMDATA.m109_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m121_ns\ : std_logic;
signal \PROM.ROMDATA.m114\ : std_logic;
signal \PROM.ROMDATA.m111\ : std_logic;
signal \PROM.ROMDATA.m120_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m120_bm\ : std_logic;
signal \PROM.ROMDATA.m121_ns_1\ : std_logic;
signal \PROM.ROMDATA.m140\ : std_logic;
signal \PROM.ROMDATA.m138_cascade_\ : std_logic;
signal \PROM.ROMDATA.m80_bm_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m80_bm\ : std_logic;
signal \N_417\ : std_logic;
signal \CONTROL_addrstack_reto_2\ : std_logic;
signal \CONTROL_programCounter11_reto_rep2\ : std_logic;
signal \PROM.ROMDATA.m135\ : std_logic;
signal \PROM.ROMDATA.m132\ : std_logic;
signal \PROM.ROMDATA.m83\ : std_logic;
signal \PROM.ROMDATA.m83_cascade_\ : std_logic;
signal \PROM.ROMDATA.m133\ : std_logic;
signal \PROM.ROMDATA.m161\ : std_logic;
signal \PROM.ROMDATA.m15\ : std_logic;
signal \PROM.ROMDATA.m171_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m162\ : std_logic;
signal \PROM.ROMDATA.m172\ : std_logic;
signal \PROM.ROMDATA.m20\ : std_logic;
signal \PROM.ROMDATA.m156\ : std_logic;
signal \PROM.ROMDATA.m171_bm\ : std_logic;
signal \PROM.ROMDATA.m383_cascade_\ : std_logic;
signal \PROM.ROMDATA.m427_bm\ : std_logic;
signal \PROM.ROMDATA.m427_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m427_ns\ : std_logic;
signal \PROM.ROMDATA.m492_am\ : std_logic;
signal \PROM.ROMDATA.m492_bm\ : std_logic;
signal \PROM.ROMDATA.m494_ns_1\ : std_logic;
signal \PROM.ROMDATA.m88\ : std_logic;
signal \PROM.ROMDATA.m514_ns_1\ : std_logic;
signal \PROM.ROMDATA.m181_cascade_\ : std_logic;
signal \PROM.ROMDATA.m514_ns\ : std_logic;
signal \PROM.ROMDATA.N_525_mux\ : std_logic;
signal \PROM.ROMDATA.m164\ : std_logic;
signal \PROM.ROMDATA.m171_am\ : std_logic;
signal \ALU.dZ0Z_12\ : std_logic;
signal \ALU.dZ0Z_13\ : std_logic;
signal \ALU.dZ0Z_14\ : std_logic;
signal \ALU.c_RNIBRG4Q9Z0Z_12\ : std_logic;
signal \ALU.c_RNIBRG4Q9_0Z0Z_12\ : std_logic;
signal \ALU.mult_555_c_RNIJF56AMZ0\ : std_logic;
signal \ALU.cZ0Z_12\ : std_logic;
signal \ALU.c_RNIO5N04A_0Z0Z_13\ : std_logic;
signal \ALU.c_RNIO5N04AZ0Z_13\ : std_logic;
signal \ALU.mult_558_c_RNIB75F9GZ0\ : std_logic;
signal \ALU.cZ0Z_13\ : std_logic;
signal \ALU.cZ0Z_14\ : std_logic;
signal \aluOperation_0\ : std_logic;
signal \ALU.a_15_d_sZ0Z_10\ : std_logic;
signal \ALU.addsub_9\ : std_logic;
signal \ALU.a_15_d_ns_sx_9\ : std_logic;
signal \ALU.status_19\ : std_logic;
signal \aluOut_2\ : std_logic;
signal \ALU.status_19_0\ : std_logic;
signal \aluOut_1\ : std_logic;
signal \ALU.d_RNIMGKJC1_0Z0Z_2\ : std_logic;
signal \ALU.d_RNIMGKJC1Z0Z_2_cascade_\ : std_logic;
signal \ALU.N_831\ : std_logic;
signal \ALU.N_863\ : std_logic;
signal \ALU.N_859_cascade_\ : std_logic;
signal \ALU.rshift_15_ns_1_1_cascade_\ : std_logic;
signal \ALU.a_15_m2_sZ0Z_1\ : std_logic;
signal \ALU.rshift_1_cascade_\ : std_logic;
signal bus_1 : std_logic;
signal \ALU.c_RNI98D92DZ0Z_15\ : std_logic;
signal \ALU.status_19_1\ : std_logic;
signal \ALU.N_968\ : std_logic;
signal \ALU.status_19_2\ : std_logic;
signal \ALU.N_867\ : std_logic;
signal \ALU.c_RNICBIG85Z0Z_15\ : std_logic;
signal \ALU.a_15_ns_snZ0Z_14\ : std_logic;
signal \ALU.lshift_14\ : std_logic;
signal \ALU.a_15_ns_rn_0_14\ : std_logic;
signal \ALU.bZ0Z_14\ : std_logic;
signal \ALU.un1_a41_8_0\ : std_logic;
signal \ALU.un1_a41_4_0\ : std_logic;
signal \ALU.un1_operation_5_0\ : std_logic;
signal \aluOperation_5\ : std_logic;
signal \ALU.un1_operation_10_0_cascade_\ : std_logic;
signal \ALU.un1_a41_7_0_2\ : std_logic;
signal \ALU.un1_operation_13Z0Z_2_cascade_\ : std_logic;
signal \ALU.un1_a41_4_0_2\ : std_logic;
signal \ALU.un1_a41_4_0_2_cascade_\ : std_logic;
signal \ALU.un1_a41_6_0\ : std_logic;
signal \aluOperation_2\ : std_logic;
signal \aluOperation_4\ : std_logic;
signal \aluOperation_3\ : std_logic;
signal \ALU.a32Z0Z_0\ : std_logic;
signal \ALU.un1_operationZ0Z_7\ : std_logic;
signal \ALU.un1_a41_2_0\ : std_logic;
signal \PROM.ROMDATA.m160\ : std_logic;
signal \aluOperation_6\ : std_logic;
signal \aluResults_0\ : std_logic;
signal \ALU.un1_a41_3_0_1_cascade_\ : std_logic;
signal \ALU.un1_a41_5_0\ : std_logic;
signal \ALU.un1_a41_7_0\ : std_logic;
signal \ALU.un1_operation_13Z0Z_2\ : std_logic;
signal \ALU.un1_operation_10_0\ : std_logic;
signal \aluReadBus\ : std_logic;
signal \ALU.un1_operation_13_0_cascade_\ : std_logic;
signal \ALU.un1_a41_9_0\ : std_logic;
signal \ALU.un1_a41_3_0_1\ : std_logic;
signal \ALU.un1_operation_13_0\ : std_logic;
signal \ALU.un1_a41_3_0\ : std_logic;
signal \aluResults_2\ : std_logic;
signal \aluResults_1\ : std_logic;
signal \ALU.un1_a41_2Z0Z_1\ : std_logic;
signal \controlWord_22\ : std_logic;
signal \CONTROL.un1_busState101_3_0_0_0\ : std_logic;
signal f_6 : std_logic;
signal \CONTROL.un1_busState101_3_0Z0Z_1\ : std_logic;
signal \A6_c\ : std_logic;
signal \INVCONTROL.ramAddReg_6C_net\ : std_logic;
signal \CONTROL.N_60\ : std_logic;
signal \PROM.ROMDATA.m281_cascade_\ : std_logic;
signal \PROM.ROMDATA.m60\ : std_logic;
signal \CONTROL.programCounter_1_7\ : std_logic;
signal \CONTROL.programCounter_1_reto_7\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \PROM.ROMDATA.m181\ : std_logic;
signal \PROM.ROMDATA.m480_bm\ : std_logic;
signal \PROM.ROMDATA.m480_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.N_551_mux\ : std_logic;
signal \progRomAddress_7\ : std_logic;
signal \PROM.ROMDATA.m480_ns_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_25ro\ : std_logic;
signal g_9 : std_logic;
signal \PROM_ROMDATA_dintern_adflt\ : std_logic;
signal \PROM_ROMDATA_dintern_25ro_cascade_\ : std_logic;
signal \PROM_ROMDATA_dintern_3ro\ : std_logic;
signal \CONTROL_romAddReg_7_9\ : std_logic;
signal \PROM.ROMDATA.m446_bm\ : std_logic;
signal \PROM.ROMDATA.m447_ns_1\ : std_logic;
signal \PROM.ROMDATA.m446_am\ : std_logic;
signal \PROM.ROMDATA.m447_ns\ : std_logic;
signal \PROM.ROMDATA.m488_ns_1\ : std_logic;
signal m125_e : std_logic;
signal \PROM.ROMDATA.N_570_mux\ : std_logic;
signal \PROM.ROMDATA.m2\ : std_logic;
signal \PROM.ROMDATA.m493_am\ : std_logic;
signal \CONTROL_addrstack_reto_1\ : std_logic;
signal \CONTROL_programCounter11_reto\ : std_logic;
signal \N_416\ : std_logic;
signal \PROM.ROMDATA.m1\ : std_logic;
signal \PROM.ROMDATA.m493_bm\ : std_logic;
signal \PROM.ROMDATA.m361_am\ : std_logic;
signal \PROM.ROMDATA.m211_ns_N_2L1\ : std_logic;
signal \PROM.ROMDATA.m211_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m221cf0_1\ : std_logic;
signal \PROM.ROMDATA.m211_ns\ : std_logic;
signal \PROM.ROMDATA.m221cf1_1\ : std_logic;
signal \PROM.ROMDATA.m369\ : std_logic;
signal \PROM.ROMDATA.m373\ : std_logic;
signal \PROM.ROMDATA.m298_ns\ : std_logic;
signal \PROM.ROMDATA.m303_ns\ : std_logic;
signal \PROM.ROMDATA.m262\ : std_logic;
signal \PROM.ROMDATA.m422_ns\ : std_logic;
signal \PROM.ROMDATA.m424\ : std_logic;
signal \PROM.ROMDATA.m361_bm\ : std_logic;
signal \PROM.ROMDATA.m127\ : std_logic;
signal \PROM.ROMDATA.m128\ : std_logic;
signal \PROM.ROMDATA.m137_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m137_bm\ : std_logic;
signal \PROM.ROMDATA.m147_am\ : std_logic;
signal \PROM.ROMDATA.m147_bm\ : std_logic;
signal \PROM.ROMDATA.m148_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m148_ns\ : std_logic;
signal \PROM.ROMDATA.m292\ : std_logic;
signal \PROM.ROMDATA.m299\ : std_logic;
signal \PROM.ROMDATA.m301\ : std_logic;
signal \PROM.ROMDATA.m357_bm\ : std_logic;
signal \PROM.ROMDATA.m357_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m178\ : std_logic;
signal \PROM.ROMDATA.m287\ : std_logic;
signal \PROM.ROMDATA.m294_ns\ : std_logic;
signal \PROM.ROMDATA.m290_cascade_\ : std_logic;
signal \PROM.ROMDATA.m303_ns_1\ : std_logic;
signal \PROM.ROMDATA.m361_ns\ : std_logic;
signal \PROM.ROMDATA.m357_ns\ : std_logic;
signal \PROM.ROMDATA.m363_ns\ : std_logic;
signal \PROM.ROMDATA.m353_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m353_bm\ : std_logic;
signal \PROM.ROMDATA.m353_ns_cascade_\ : std_logic;
signal \PROM.ROMDATA.m363_ns_1\ : std_logic;
signal \PROM.ROMDATA.m347\ : std_logic;
signal \PROM.ROMDATA.m112\ : std_logic;
signal \PROM.ROMDATA.m349_am\ : std_logic;
signal \PROM.ROMDATA.m349_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m349_ns\ : std_logic;
signal \PROM.ROMDATA.m331_bm_cascade_\ : std_logic;
signal \PROM.ROMDATA.m323_bm\ : std_logic;
signal \PROM.ROMDATA.m323_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m323_ns\ : std_logic;
signal \aluParams_1\ : std_logic;
signal \ALU.un14_log_0_0_15\ : std_logic;
signal \ALU.status_19_14\ : std_logic;
signal \ALU.N_586\ : std_logic;
signal \PROM.ROMDATA.m331_am\ : std_logic;
signal \PROM.ROMDATA.m331_ns\ : std_logic;
signal \progRomAddress_5\ : std_logic;
signal \progRomAddress_6\ : std_logic;
signal \PROM.ROMDATA.m343_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.m343_ns\ : std_logic;
signal \PROM.ROMDATA.m4\ : std_logic;
signal \PROM.ROMDATA.N_28_i\ : std_logic;
signal \PROM.ROMDATA.m183\ : std_logic;
signal \PROM.ROMDATA.m334_ns_1_cascade_\ : std_logic;
signal \PROM.ROMDATA.i3_mux_0\ : std_logic;
signal \progRomAddress_1\ : std_logic;
signal \progRomAddress_2\ : std_logic;
signal \progRomAddress_0\ : std_logic;
signal \PROM.ROMDATA.m338_bm\ : std_logic;
signal \PROM.ROMDATA.m338_am_cascade_\ : std_logic;
signal \PROM.ROMDATA.m338_ns\ : std_logic;
signal \PROM.ROMDATA.m246\ : std_logic;
signal \progRomAddress_4\ : std_logic;
signal \PROM.ROMDATA.m341_ns_1\ : std_logic;
signal \progRomAddress_3\ : std_logic;
signal \PROM.ROMDATA.m341_ns\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \BUFFER_ADDRESS_wire\ : std_logic_vector(15 downto 0);
signal \D3_wire\ : std_logic;
signal \BUFFER_DATA_IN_wire\ : std_logic_vector(15 downto 0);
signal \D10_wire\ : std_logic;
signal \D7_wire\ : std_logic;
signal \B_CE_wire\ : std_logic;
signal \D0_wire\ : std_logic;
signal \BUFFER_DATA_OUT_wire\ : std_logic_vector(15 downto 0);
signal \D9_in_wire\ : std_logic;
signal \D6_wire\ : std_logic;
signal \D10_in_wire\ : std_logic;
signal \D2_wire\ : std_logic;
signal \D4_in_wire\ : std_logic;
signal \A4_wire\ : std_logic;
signal \D0_in_wire\ : std_logic;
signal \A10_wire\ : std_logic;
signal \D3_in_wire\ : std_logic;
signal \UB_wire\ : std_logic;
signal \B_LB_wire\ : std_logic;
signal \D15_wire\ : std_logic;
signal \D14_in_wire\ : std_logic;
signal \A6_wire\ : std_logic;
signal \WR_wire\ : std_logic;
signal \D13_wire\ : std_logic;
signal \D11_in_wire\ : std_logic;
signal \A8_wire\ : std_logic;
signal \A9_wire\ : std_logic;
signal \LB_wire\ : std_logic;
signal \D8_wire\ : std_logic;
signal \A7_wire\ : std_logic;
signal \OE_wire\ : std_logic;
signal \GPIO3_wire\ : std_logic;
signal \D2_in_wire\ : std_logic;
signal \A14_wire\ : std_logic;
signal \A5_wire\ : std_logic;
signal \D9_wire\ : std_logic;
signal \D11_wire\ : std_logic;
signal \D12_in_wire\ : std_logic;
signal \A15_wire\ : std_logic;
signal \A13_wire\ : std_logic;
signal \A1_wire\ : std_logic;
signal \B_UB_wire\ : std_logic;
signal \D7_in_wire\ : std_logic;
signal \B_WR_wire\ : std_logic;
signal \GPIO11_wire\ : std_logic;
signal \A2_wire\ : std_logic;
signal \D5_wire\ : std_logic;
signal \D4_wire\ : std_logic;
signal \A3_wire\ : std_logic;
signal \A11_wire\ : std_logic;
signal \GPIO9_wire\ : std_logic;
signal \D5_in_wire\ : std_logic;
signal \D15_in_wire\ : std_logic;
signal \D1_in_wire\ : std_logic;
signal \B_OE_wire\ : std_logic;
signal \D12_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \D8_in_wire\ : std_logic;
signal \D6_in_wire\ : std_logic;
signal \D13_in_wire\ : std_logic;
signal \D1_wire\ : std_logic;
signal \A12_wire\ : std_logic;
signal \A0_wire\ : std_logic;
signal \CE_wire\ : std_logic;
signal \D14_wire\ : std_logic;
signal \DROM.ROMDATA.dintern_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \DROM.ROMDATA.dintern_0_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \DROM.ROMDATA.dintern_0_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \CONTROL.addrstack_addrstack_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \CONTROL.addrstack_addrstack_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \CONTROL.addrstack_addrstack_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \CONTROL.addrstack_addrstack_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \CLK_wire\ <= CLK;
    BUFFER_ADDRESS <= \BUFFER_ADDRESS_wire\;
    D3 <= \D3_wire\;
    \BUFFER_DATA_IN_wire\ <= BUFFER_DATA_IN;
    D10 <= \D10_wire\;
    D7 <= \D7_wire\;
    B_CE <= \B_CE_wire\;
    D0 <= \D0_wire\;
    BUFFER_DATA_OUT <= \BUFFER_DATA_OUT_wire\;
    \D9_in_wire\ <= D9_in;
    D6 <= \D6_wire\;
    \D10_in_wire\ <= D10_in;
    D2 <= \D2_wire\;
    \D4_in_wire\ <= D4_in;
    A4 <= \A4_wire\;
    \D0_in_wire\ <= D0_in;
    A10 <= \A10_wire\;
    \D3_in_wire\ <= D3_in;
    UB <= \UB_wire\;
    B_LB <= \B_LB_wire\;
    D15 <= \D15_wire\;
    \D14_in_wire\ <= D14_in;
    A6 <= \A6_wire\;
    WR <= \WR_wire\;
    D13 <= \D13_wire\;
    \D11_in_wire\ <= D11_in;
    A8 <= \A8_wire\;
    A9 <= \A9_wire\;
    LB <= \LB_wire\;
    D8 <= \D8_wire\;
    A7 <= \A7_wire\;
    OE <= \OE_wire\;
    GPIO3 <= \GPIO3_wire\;
    \D2_in_wire\ <= D2_in;
    A14 <= \A14_wire\;
    A5 <= \A5_wire\;
    D9 <= \D9_wire\;
    D11 <= \D11_wire\;
    \D12_in_wire\ <= D12_in;
    A15 <= \A15_wire\;
    A13 <= \A13_wire\;
    A1 <= \A1_wire\;
    B_UB <= \B_UB_wire\;
    \D7_in_wire\ <= D7_in;
    B_WR <= \B_WR_wire\;
    GPIO11 <= \GPIO11_wire\;
    A2 <= \A2_wire\;
    D5 <= \D5_wire\;
    D4 <= \D4_wire\;
    A3 <= \A3_wire\;
    A11 <= \A11_wire\;
    GPIO9 <= \GPIO9_wire\;
    \D5_in_wire\ <= D5_in;
    \D15_in_wire\ <= D15_in;
    \D1_in_wire\ <= D1_in;
    B_OE <= \B_OE_wire\;
    D12 <= \D12_wire\;
    TX <= \TX_wire\;
    \D8_in_wire\ <= D8_in;
    \D6_in_wire\ <= D6_in;
    \D13_in_wire\ <= D13_in;
    D1 <= \D1_wire\;
    A12 <= \A12_wire\;
    A0 <= \A0_wire\;
    CE <= \CE_wire\;
    D14 <= \D14_wire\;
    \DROM.ROMDATA.dintern_0_0_NEW_3\ <= \DROM.ROMDATA.dintern_0_0_physical_RDATA_wire\(13);
    \DROM.ROMDATA.dintern_0_0_NEW_2\ <= \DROM.ROMDATA.dintern_0_0_physical_RDATA_wire\(9);
    \DROM.ROMDATA.dintern_0_0_NEW_1\ <= \DROM.ROMDATA.dintern_0_0_physical_RDATA_wire\(5);
    \DROM.ROMDATA.dintern_0_0_NEW_0\ <= \DROM.ROMDATA.dintern_0_0_physical_RDATA_wire\(1);
    \DROM.ROMDATA.dintern_0_0_physical_RADDR_wire\ <= '0'&\N__71657\&\N__26564\&\N__26639\&\N__26606\&\N__26369\&\N__26537\&\N__26399\&\N__26432\&\N__33233\&\N__33293\;
    \DROM.ROMDATA.dintern_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_1_NEW_3\ <= \DROM.ROMDATA.dintern_0_1_physical_RDATA_wire\(13);
    \DROM.ROMDATA.dintern_0_1_NEW_2\ <= \DROM.ROMDATA.dintern_0_1_physical_RDATA_wire\(9);
    \DROM.ROMDATA.dintern_0_1_NEW_1\ <= \DROM.ROMDATA.dintern_0_1_physical_RDATA_wire\(5);
    \DROM.ROMDATA.dintern_0_1_NEW_0\ <= \DROM.ROMDATA.dintern_0_1_physical_RDATA_wire\(1);
    \DROM.ROMDATA.dintern_0_1_physical_RADDR_wire\ <= '0'&\N__71651\&\N__26558\&\N__26633\&\N__26600\&\N__26363\&\N__26531\&\N__26393\&\N__26426\&\N__33227\&\N__33287\;
    \DROM.ROMDATA.dintern_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_2_NEW_3\ <= \DROM.ROMDATA.dintern_0_2_physical_RDATA_wire\(13);
    \DROM.ROMDATA.dintern_0_2_NEW_2\ <= \DROM.ROMDATA.dintern_0_2_physical_RDATA_wire\(9);
    \DROM.ROMDATA.dintern_0_2_NEW_1\ <= \DROM.ROMDATA.dintern_0_2_physical_RDATA_wire\(5);
    \DROM.ROMDATA.dintern_0_2_NEW_0\ <= \DROM.ROMDATA.dintern_0_2_physical_RDATA_wire\(1);
    \DROM.ROMDATA.dintern_0_2_physical_RADDR_wire\ <= '0'&\N__71645\&\N__26552\&\N__26627\&\N__26594\&\N__26357\&\N__26525\&\N__26387\&\N__26420\&\N__33221\&\N__33281\;
    \DROM.ROMDATA.dintern_0_2_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_3_NEW_3\ <= \DROM.ROMDATA.dintern_0_3_physical_RDATA_wire\(13);
    \DROM.ROMDATA.dintern_0_3_NEW_2\ <= \DROM.ROMDATA.dintern_0_3_physical_RDATA_wire\(9);
    \DROM.ROMDATA.dintern_0_3_NEW_1\ <= \DROM.ROMDATA.dintern_0_3_physical_RDATA_wire\(5);
    \DROM.ROMDATA.dintern_0_3_NEW_0\ <= \DROM.ROMDATA.dintern_0_3_physical_RDATA_wire\(1);
    \DROM.ROMDATA.dintern_0_3_physical_RADDR_wire\ <= '0'&\N__71639\&\N__26546\&\N__26621\&\N__26588\&\N__26351\&\N__26519\&\N__26381\&\N__26414\&\N__33215\&\N__33275\;
    \DROM.ROMDATA.dintern_0_3_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \DROM.ROMDATA.dintern_0_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \CONTROL.addrstack_15\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(15);
    \CONTROL.addrstack_14\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(14);
    \CONTROL.addrstack_13\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(13);
    \CONTROL.addrstack_12\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(12);
    \CONTROL.addrstack_11\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(11);
    \CONTROL.addrstack_10\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(10);
    \CONTROL.addrstack_9\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(9);
    \CONTROL.addrstack_8\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(8);
    \CONTROL.addrstack_7\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(7);
    \CONTROL.addrstack_6\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(6);
    \CONTROL.addrstack_5\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(5);
    \CONTROL.addrstack_4\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(4);
    \CONTROL.addrstack_3\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(3);
    \CONTROL.addrstack_2\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(2);
    \CONTROL.addrstackZ0Z_1\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(1);
    \CONTROL.addrstack_0\ <= \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\(0);
    \CONTROL.addrstack_addrstack_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__41885\&\N__26690\&\N__27554\&\N__29663\&\N__34619\&\N__38369\&\N__29777\&\N__29765\;
    \CONTROL.addrstack_addrstack_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__42322\&\N__26724\&\N__27528\&\N__29700\&\N__34795\&\N__38461\&\N__31524\&\N__33797\;
    \CONTROL.addrstack_addrstack_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \CONTROL.addrstack_addrstack_0_0_physical_WDATA_wire\ <= \N__27725\&\N__27713\&\N__26657\&\N__33509\&\N__27737\&\N__28505\&\N__28481\&\N__33569\&\N__33524\&\N__26651\&\N__33620\&\N__33554\&\N__33605\&\N__33497\&\N__33539\&\N__33635\;

    \DROM.ROMDATA.dintern_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0001000100010001000000000000000100010001000100010000000000000001000100000000000100000001000000010000000000010000000000010001000000010001000000010001000100010001000100010001000000010000000000010001000100010000000000000001000000000001000000010001000100010001",
            INIT_E => "0001000100010000000000000000000100010001000100000001000100010001000100010001000000010001000100010001000100010001000000010001000000010001000100010000000000000000000000000000000000010001000100010001000000010001000000010000000000010001000100010001000100010001",
            INIT_D => "0000000000000000000100000000000000000000000000010001000100010001000000000000000100010001000100010000000100000000000100010001000100010001000000010000000100000001000100010001000000000001000000010000000100000001000100010001000100000001000000010000000100000001",
            INIT_C => "0001000100010001000100010001000000000000000000010001000100010001000000000000000100000000000000010001000100010000000100000001000000000001000000010001000100010001000100010001000000000001000000010001000100010000000000010001000000000001000000010001000100010000",
            INIT_B => "0000000000010001000000010000000100000000010001010000000101000100010100000001010001100000000000010011000000010000001100000001010000110000010100000000010001000101000100000001000000000101000000000100000000000000000101000001010000000100000000000000000000000000",
            INIT_A => "0001010000010000010001000100000000010001000101010000000100000001000001010001010100010101000100010100000100000101000100010101000100000000000100010000000101000101000100000000000100010101010001010100010101000001010100010001010001010000010001010000000101000001",
            INIT_9 => "0100010101010101000101010101010100000001000000000100000101010001000101000001010001000101000000010000000000000001010001000001010001000001000001010001000001000101010000000100000000010001000100010000010000010100000101010101000100000000000001010101000100010000",
            INIT_8 => "0000000000010001000001010100010001010100010001000100010001000000000000000000000001000000000001000000000101000100000001010000010001000001010001000100010001000000000100000000000000000000000000000100010101000100010101010101010000000001000000000000000100000001",
            INIT_7 => "0010001000110010001000110010001100100010001000100001000100010010000000000010001100000000001000010001001100010000001000000010001000000000000000100000000000010001001000000010001000010001000000000000000100010011001100010011001100000010000100000000001100100000",
            INIT_6 => "0011001000100001001000010010000100110011001100010011000000010000000100110011000100010000001100000011001100010001000000000011000100100010001000000010001000010001001000100010000000100011001100010010000000000000001000100010000000100010001000000000000000000000",
            INIT_5 => "0011001100110001000100010011000100110011001100110001000100110001001000000010000100110011001100010001001100010001000000000010000100010001001100010011001100010001001000100010000100010001001100010011001100010001001000100000000100010001001100010011001100110001",
            INIT_4 => "0010001000000001000100010011000100110011000100010010001000000001000100010011000100110011001100010010001000100001001100110011000100110011001100010000000000000001001100110011001100010001000100110000000000100001001100110001000100110011001100110010001000000011",
            INIT_3 => "0001000100010001000100010001000100000000000000010011001100010011000100010001000101100010000000010101000100110001011100110011001101100010001000010011000100110001001100110001000100000010000000110011001100110001000100110001000100000010001000010011000100110001",
            INIT_2 => "0011001100010001001000100010001100010001001100010011001100010001000000000010000100010001001100010011001100010001001000100000000100010001001100010011001100110011001000100000000100010011001100010011000100110001000000000000000100010001001100010001000100010011",
            INIT_1 => "0000000000000001000100010001000100010001000100010000000000100001000100010001001100010001001100010010001000100011000100010001001100010001000100110010000000000001000100110001000100010001001100010000000000000011000100010001001100110011001100110000000000100011",
            INIT_0 => "0001001100010011001100010001001100000000001000110011001100010001000100010011001100100000001000110001001100010001001100010011001100100010001000110011001100010001001100110011001100000010001000110011000100010001000100110011001100100010001000110001000100010001"
        )
    port map (
            RDATA => \DROM.ROMDATA.dintern_0_0_physical_RDATA_wire\,
            RADDR => \DROM.ROMDATA.dintern_0_0_physical_RADDR_wire\,
            WADDR => \DROM.ROMDATA.dintern_0_0_physical_WADDR_wire\,
            MASK => \DROM.ROMDATA.dintern_0_0_physical_MASK_wire\,
            WDATA => \DROM.ROMDATA.dintern_0_0_physical_WDATA_wire\,
            RCLKE => \N__28122\,
            RCLK => \INVDROM.ROMDATA.dintern_0_0RCLKN_net\,
            RE => \N__32495\,
            WCLKE => \N__35927\,
            WCLK => \GNDG0\,
            WE => 'L'
        );

    \DROM.ROMDATA.dintern_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000010010001000000001000000100000000100100010000000000010000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000001",
            INIT_E => "0000000000000000000000000000000100000000000000000000000000000001000000000000000000100010001000010000000000100001001000100010000000100010001000010010001000000001001000000000000100000000000000010000000000000001000000000000000000000000000000010000000000000000",
            INIT_D => "0000000000000001000000000000000000000000000000010000000000000001000000000000000100100010001000110010000000000010001000100010001100100010001000110010001000100001001000100000000000000000000000000000000000000000000000000000000100000000000000010000000000000001",
            INIT_C => "0000000000000001000000000000000000000000000000010000000000000001000000000000000100100010001000110010000000000010001000100010001000000010001000110010001000100001001000100000000100000000000000000000000000000001000000000000000100000000000000010000000000000000",
            INIT_B => "0000000000000000000000000000000100000100010001000000010001000000000001000100000000000110011000110010011001000100000001100110001000100100011001100010011001100011001000100110000000000100010001000000010001000100000001000100000000000100010001010000000001000000",
            INIT_A => "0000010001000000000001000100000000000100010000000000000001000001000001000100000100100110011001110010010001000011001001100110011100000110011001100010011001100100001000100100000100000100010000010000010001000001000001000100000100000100010000000000010001000101",
            INIT_9 => "0000010001000001000001000100010100000000010000000000000001000000000001000100000000100110011000010000010001100101001001100110000100100110011000010010011001000101000000000100000000000000010000010000010001000000000001000100010000000100010000010000010001000001",
            INIT_8 => "0000000001000000000001000100010000000100010000010000010001000000000000000100000100100110001000000000000001100100011001100010000001100010011000000010011001000000000000000100000000000000010000010100010001000100010001000100010000000000000000000000000000000000",
            INIT_7 => "0000000000000010000000000000001000000000000000100000000000000000000000000000000100000000000000010000000000000000000000000000001000000000000000100000000000000000000000000000001000000000000000010000000000000011000000000000001000000000000000010000000000000010",
            INIT_6 => "0000000000000010000000000000001000000000000000110000000000100000000000000000000100000000000000100000000000000001000000000000001000000000000000100000000000000010000000000000001000000000000000010000000000000010000000000000000000000000000000100000000000000010",
            INIT_5 => "0000000000000001000000000000001100000000000000110000000000000001000000000000000100000000010000110100010001000011000000000100000101000100010000010100010000000011010001000010001101000000000000110100000000000001010000000000000100000000000000110000000000100011",
            INIT_4 => "0000000000000001000000000000001101000100000000010100010000000011010001000000000101000000000001110100010001000111010000000000010101000100010001110100010001000011010001000100001101000100010000110100010000000011010001000000000101000100000000110000000000000011",
            INIT_3 => "0000000000100001000000000000001101000100000000010100010000000011010001000000000101000100000000110100010001000101010001000000001101000100010001110100010001100101010001000100010100000100010000010000010001000011010001000000000101000100000000110000000000000011",
            INIT_2 => "0000000000000001000000000000001100000000000000110100000000000001010000000000001101000000000001110100010001000101010000000000010101000100010001110100010001000011010001000100001101000100000000110100010000000011010000000000000100000000000000010000000000000001",
            INIT_1 => "0000000000000011000000000000001100000000000000110000000000000001000000000000000100000000010000010100010001000011000000000100001101000100010000110100010000000001010000000000000100000000000000010000000000000011000000000000001100000000000000110000000000000011",
            INIT_0 => "0000000000000011000000000000001100000000000000010000000000000011000000000000000100000100010000110100010001000001000001000100001101000100010000110100010000000001010000000000001100000000000000010000000000000011000000000000000100000000000000110000000000000011"
        )
    port map (
            RDATA => \DROM.ROMDATA.dintern_0_1_physical_RDATA_wire\,
            RADDR => \DROM.ROMDATA.dintern_0_1_physical_RADDR_wire\,
            WADDR => \DROM.ROMDATA.dintern_0_1_physical_WADDR_wire\,
            MASK => \DROM.ROMDATA.dintern_0_1_physical_MASK_wire\,
            WDATA => \DROM.ROMDATA.dintern_0_1_physical_WDATA_wire\,
            RCLKE => \N__28112\,
            RCLK => \INVDROM.ROMDATA.dintern_0_1RCLKN_net\,
            RE => \N__32513\,
            WCLKE => \N__35928\,
            WCLK => \GNDG0\,
            WE => 'L'
        );

    \DROM.ROMDATA.dintern_0_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000010001000100010001000100010000000100010001000100010001000100010000000100010001000100010001000000010001000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000001000100010001000100010001000100010001000100000000000100010000000100010001000000010001000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000010001000100010000000100010001000100010000000000010001000100010001000000010001000000000001000100000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000010000000000000001000100000000000100010001000000010001000100010001000100000000000100010001000100010000000100010001000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000010001000000000001000100010000000100010001000100000001000100010000000100010000000000010001000100010001000000010001000100000001000100000000000000010000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000010000000000000001000100000000000100010001000100000001000100010000000100000001000100000001000000010000000100010001000000010001000100000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000001000000000000000100010001000100010001000100010001000100010001000100000000000100000001000100010000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001000100010001000100010000000100110001000100010001000100110010000100110000000100010001000000010001000100000001000100000010001000100010000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000010000000000000001000100000001000100010001000100010001000100010001000100010001000100010001000100010001000100000001000100010000000000010001000000000000000100000000000000010000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000100000001000100010001000100010001000100010001000000010001000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000010000000000000001000100000000000100010000000100010001000100010001000100010001000100010001000100000001000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000100000000000000010001000000010001000100000001000100010001000100010001000100010001000100010001000100010000000000000000000000000001000000000000000100000000000000010000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000100010000000100010001000000010001000100010001000100010001000100010001000100010001000100000000000100010000000000010001000000010001000000000001000100000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000000000010001000100010001000100000001000100010001000100010001000100000000000100010000000100010001000100010001000000010001000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \DROM.ROMDATA.dintern_0_2_physical_RDATA_wire\,
            RADDR => \DROM.ROMDATA.dintern_0_2_physical_RADDR_wire\,
            WADDR => \DROM.ROMDATA.dintern_0_2_physical_WADDR_wire\,
            MASK => \DROM.ROMDATA.dintern_0_2_physical_MASK_wire\,
            WDATA => \DROM.ROMDATA.dintern_0_2_physical_WDATA_wire\,
            RCLKE => \N__28123\,
            RCLK => \INVDROM.ROMDATA.dintern_0_2RCLKN_net\,
            RE => \N__32514\,
            WCLKE => \N__35929\,
            WCLK => \GNDG0\,
            WE => 'L'
        );

    \DROM.ROMDATA.dintern_0_3_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001000100010001000000010001000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000001000100000001000100000000000100010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100010001000100000001000100000001000000000000000100000000000100010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000001000100000000000100010001000100010001000100010000000000010001000000000000000000000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000001000100010000000100010001000000000001000100000000000000010000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000001000100000000000100010000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000010000000000010001000000000001000100000001000100000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000100001000000000000000000000010001100110000000100010001000100010011000000000001000000000010001000100010000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000001000100000000000100010001000000000000000100000000000000010000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000001000100000000000100010000000000010001000000000000000100000000000000010000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000100010000000000010001000000000001000100000000000000010000000000000001000000000000000000000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000100000000000100010000000000000001000000000001000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \DROM.ROMDATA.dintern_0_3_physical_RDATA_wire\,
            RADDR => \DROM.ROMDATA.dintern_0_3_physical_RADDR_wire\,
            WADDR => \DROM.ROMDATA.dintern_0_3_physical_WADDR_wire\,
            MASK => \DROM.ROMDATA.dintern_0_3_physical_MASK_wire\,
            WDATA => \DROM.ROMDATA.dintern_0_3_physical_WDATA_wire\,
            RCLKE => \N__28124\,
            RCLK => \INVDROM.ROMDATA.dintern_0_3RCLKN_net\,
            RE => \N__32530\,
            WCLKE => \N__35930\,
            WCLK => \GNDG0\,
            WE => 'L'
        );

    \CONTROL.addrstack_addrstack_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \CONTROL.addrstack_addrstack_0_0_physical_RDATA_wire\,
            RADDR => \CONTROL.addrstack_addrstack_0_0_physical_RADDR_wire\,
            WADDR => \CONTROL.addrstack_addrstack_0_0_physical_WADDR_wire\,
            MASK => \CONTROL.addrstack_addrstack_0_0_physical_MASK_wire\,
            WDATA => \CONTROL.addrstack_addrstack_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \INVCONTROL.addrstack_addrstack_0_0RCLKN_net\,
            RE => \N__32544\,
            WCLKE => \N__28367\,
            WCLK => \N__73292\,
            WE => \N__32563\
        );

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__80916\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80918\,
            DIN => \N__80917\,
            DOUT => \N__80916\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80918\,
            PADOUT => \N__80917\,
            PADIN => \N__80916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80907\,
            DIN => \N__80906\,
            DOUT => \N__80905\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(15)
        );

    \BUFFER_ADDRESS_obuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80907\,
            PADOUT => \N__80906\,
            PADIN => \N__80905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26453\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D3_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80898\,
            DIN => \N__80897\,
            DOUT => \N__80896\,
            PACKAGEPIN => \D3_wire\
        );

    \D3_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80898\,
            PADOUT => \N__80897\,
            PADIN => \N__80896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35113\,
            DIN0 => OPEN,
            DOUT0 => \N__34244\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80889\,
            DIN => \N__80888\,
            DOUT => \N__80887\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(12)
        );

    \BUFFER_DATA_IN_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80889\,
            PADOUT => \N__80888\,
            PADIN => \N__80887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80880\,
            DIN => \N__80879\,
            DOUT => \N__80878\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(4)
        );

    \BUFFER_ADDRESS_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80880\,
            PADOUT => \N__80879\,
            PADIN => \N__80878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29312\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D10_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80871\,
            DIN => \N__80870\,
            DOUT => \N__80869\,
            PACKAGEPIN => \D10_wire\
        );

    \D10_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80871\,
            PADOUT => \N__80870\,
            PADIN => \N__80869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35050\,
            DIN0 => OPEN,
            DOUT0 => \N__26228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D7_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80862\,
            DIN => \N__80861\,
            DOUT => \N__80860\,
            PACKAGEPIN => \D7_wire\
        );

    \D7_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80862\,
            PADOUT => \N__80861\,
            PADIN => \N__80860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35102\,
            DIN0 => OPEN,
            DOUT0 => \N__46043\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80853\,
            DIN => \N__80852\,
            DOUT => \N__80851\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(2)
        );

    \BUFFER_DATA_IN_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80853\,
            PADOUT => \N__80852\,
            PADIN => \N__80851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_CE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80844\,
            DIN => \N__80843\,
            DOUT => \N__80842\,
            PACKAGEPIN => \B_CE_wire\
        );

    \B_CE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80844\,
            PADOUT => \N__80843\,
            PADIN => \N__80842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32493\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D0_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80835\,
            DIN => \N__80834\,
            DOUT => \N__80833\,
            PACKAGEPIN => \D0_wire\
        );

    \D0_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80835\,
            PADOUT => \N__80834\,
            PADIN => \N__80833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35117\,
            DIN0 => OPEN,
            DOUT0 => \N__37688\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80826\,
            DIN => \N__80825\,
            DOUT => \N__80824\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(8)
        );

    \BUFFER_DATA_OUT_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80826\,
            PADOUT => \N__80825\,
            PADIN => \N__80824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26131\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D9_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80817\,
            DIN => \N__80816\,
            DOUT => \N__80815\,
            PACKAGEPIN => \D9_in_wire\
        );

    \D9_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80817\,
            PADOUT => \N__80816\,
            PADIN => \N__80815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D9_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80808\,
            DIN => \N__80807\,
            DOUT => \N__80806\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(13)
        );

    \BUFFER_DATA_OUT_obuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80808\,
            PADOUT => \N__80807\,
            PADIN => \N__80806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80799\,
            DIN => \N__80798\,
            DOUT => \N__80797\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(8)
        );

    \BUFFER_DATA_IN_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80799\,
            PADOUT => \N__80798\,
            PADIN => \N__80797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80790\,
            DIN => \N__80789\,
            DOUT => \N__80788\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(8)
        );

    \BUFFER_ADDRESS_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80790\,
            PADOUT => \N__80789\,
            PADIN => \N__80788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29234\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80781\,
            DIN => \N__80780\,
            DOUT => \N__80779\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(12)
        );

    \BUFFER_ADDRESS_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80781\,
            PADOUT => \N__80780\,
            PADIN => \N__80779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26492\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D6_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80772\,
            DIN => \N__80771\,
            DOUT => \N__80770\,
            PACKAGEPIN => \D6_wire\
        );

    \D6_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80772\,
            PADOUT => \N__80771\,
            PADIN => \N__80770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35071\,
            DIN0 => OPEN,
            DOUT0 => \N__63380\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D10_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80763\,
            DIN => \N__80762\,
            DOUT => \N__80761\,
            PACKAGEPIN => \D10_in_wire\
        );

    \D10_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80763\,
            PADOUT => \N__80762\,
            PADIN => \N__80761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D10_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D2_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80754\,
            DIN => \N__80753\,
            DOUT => \N__80752\,
            PACKAGEPIN => \D2_wire\
        );

    \D2_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80754\,
            PADOUT => \N__80753\,
            PADIN => \N__80752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35099\,
            DIN0 => OPEN,
            DOUT0 => \N__43481\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D4_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80745\,
            DIN => \N__80744\,
            DOUT => \N__80743\,
            PACKAGEPIN => \D4_in_wire\
        );

    \D4_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80745\,
            PADOUT => \N__80744\,
            PADIN => \N__80743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D4_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80736\,
            DIN => \N__80735\,
            DOUT => \N__80734\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(13)
        );

    \BUFFER_DATA_IN_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80736\,
            PADOUT => \N__80735\,
            PADIN => \N__80734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80727\,
            DIN => \N__80726\,
            DOUT => \N__80725\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(5)
        );

    \BUFFER_DATA_OUT_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80727\,
            PADOUT => \N__80726\,
            PADIN => \N__80725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__52531\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80718\,
            DIN => \N__80717\,
            DOUT => \N__80716\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(7)
        );

    \BUFFER_DATA_IN_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80718\,
            PADOUT => \N__80717\,
            PADIN => \N__80716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80709\,
            DIN => \N__80708\,
            DOUT => \N__80707\,
            PACKAGEPIN => \A4_wire\
        );

    \A4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80709\,
            PADOUT => \N__80708\,
            PADIN => \N__80707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__44072\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80700\,
            DIN => \N__80699\,
            DOUT => \N__80698\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(7)
        );

    \BUFFER_ADDRESS_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80700\,
            PADOUT => \N__80699\,
            PADIN => \N__80698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29252\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D0_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80691\,
            DIN => \N__80690\,
            DOUT => \N__80689\,
            PACKAGEPIN => \D0_in_wire\
        );

    \D0_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80691\,
            PADOUT => \N__80690\,
            PADIN => \N__80689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D0_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A10_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80682\,
            DIN => \N__80681\,
            DOUT => \N__80680\,
            PACKAGEPIN => \A10_wire\
        );

    \A10_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80682\,
            PADOUT => \N__80681\,
            PADIN => \N__80680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31202\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80673\,
            DIN => \N__80672\,
            DOUT => \N__80671\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(9)
        );

    \BUFFER_DATA_OUT_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80673\,
            PADOUT => \N__80672\,
            PADIN => \N__80671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__40385\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80664\,
            DIN => \N__80663\,
            DOUT => \N__80662\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(12)
        );

    \BUFFER_DATA_OUT_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80664\,
            PADOUT => \N__80663\,
            PADIN => \N__80662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26320\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D3_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80655\,
            DIN => \N__80654\,
            DOUT => \N__80653\,
            PACKAGEPIN => \D3_in_wire\
        );

    \D3_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80655\,
            PADOUT => \N__80654\,
            PADIN => \N__80653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D3_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80646\,
            DIN => \N__80645\,
            DOUT => \N__80644\,
            PACKAGEPIN => \UB_wire\
        );

    \UB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80646\,
            PADOUT => \N__80645\,
            PADIN => \N__80644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25684\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_LB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80637\,
            DIN => \N__80636\,
            DOUT => \N__80635\,
            PACKAGEPIN => \B_LB_wire\
        );

    \B_LB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80637\,
            PADOUT => \N__80636\,
            PADIN => \N__80635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25791\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D15_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80628\,
            DIN => \N__80627\,
            DOUT => \N__80626\,
            PACKAGEPIN => \D15_wire\
        );

    \D15_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80628\,
            PADOUT => \N__80627\,
            PADIN => \N__80626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35025\,
            DIN0 => OPEN,
            DOUT0 => \N__49219\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80619\,
            DIN => \N__80618\,
            DOUT => \N__80617\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(13)
        );

    \BUFFER_ADDRESS_obuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80619\,
            PADOUT => \N__80618\,
            PADIN => \N__80617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26474\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D14_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80610\,
            DIN => \N__80609\,
            DOUT => \N__80608\,
            PACKAGEPIN => \D14_in_wire\
        );

    \D14_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80610\,
            PADOUT => \N__80609\,
            PADIN => \N__80608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D14_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A6_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80601\,
            DIN => \N__80600\,
            DOUT => \N__80599\,
            PACKAGEPIN => \A6_wire\
        );

    \A6_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80601\,
            PADOUT => \N__80600\,
            PADIN => \N__80599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__70373\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80592\,
            DIN => \N__80591\,
            DOUT => \N__80590\,
            PACKAGEPIN => \WR_wire\
        );

    \WR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80592\,
            PADOUT => \N__80591\,
            PADIN => \N__80590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25672\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D13_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80583\,
            DIN => \N__80582\,
            DOUT => \N__80581\,
            PACKAGEPIN => \D13_wire\
        );

    \D13_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80583\,
            PADOUT => \N__80582\,
            PADIN => \N__80581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35007\,
            DIN0 => OPEN,
            DOUT0 => \N__27242\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80574\,
            DIN => \N__80573\,
            DOUT => \N__80572\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(10)
        );

    \BUFFER_DATA_IN_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80574\,
            PADOUT => \N__80573\,
            PADIN => \N__80572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D11_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80565\,
            DIN => \N__80564\,
            DOUT => \N__80563\,
            PACKAGEPIN => \D11_in_wire\
        );

    \D11_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80565\,
            PADOUT => \N__80564\,
            PADIN => \N__80563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D11_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A8_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80556\,
            DIN => \N__80555\,
            DOUT => \N__80554\,
            PACKAGEPIN => \A8_wire\
        );

    \A8_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80556\,
            PADOUT => \N__80555\,
            PADIN => \N__80554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31058\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80547\,
            DIN => \N__80546\,
            DOUT => \N__80545\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(2)
        );

    \BUFFER_DATA_OUT_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80547\,
            PADOUT => \N__80546\,
            PADIN => \N__80545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__43474\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80538\,
            DIN => \N__80537\,
            DOUT => \N__80536\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(6)
        );

    \BUFFER_DATA_IN_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80538\,
            PADOUT => \N__80537\,
            PADIN => \N__80536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80529\,
            DIN => \N__80528\,
            DOUT => \N__80527\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(6)
        );

    \BUFFER_ADDRESS_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80529\,
            PADOUT => \N__80528\,
            PADIN => \N__80527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29267\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A9_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80520\,
            DIN => \N__80519\,
            DOUT => \N__80518\,
            PACKAGEPIN => \A9_wire\
        );

    \A9_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80520\,
            PADOUT => \N__80519\,
            PADIN => \N__80518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31112\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80511\,
            DIN => \N__80510\,
            DOUT => \N__80509\,
            PACKAGEPIN => \LB_wire\
        );

    \LB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80511\,
            PADOUT => \N__80510\,
            PADIN => \N__80509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25688\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80502\,
            DIN => \N__80501\,
            DOUT => \N__80500\,
            PACKAGEPIN => \D8_wire\
        );

    \D8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80502\,
            PADOUT => \N__80501\,
            PADIN => \N__80500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35100\,
            DIN0 => OPEN,
            DOUT0 => \N__26138\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80493\,
            DIN => \N__80492\,
            DOUT => \N__80491\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(11)
        );

    \BUFFER_DATA_OUT_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80493\,
            PADOUT => \N__80492\,
            PADIN => \N__80491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37354\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80484\,
            DIN => \N__80483\,
            DOUT => \N__80482\,
            PACKAGEPIN => \A7_wire\
        );

    \A7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80484\,
            PADOUT => \N__80483\,
            PADIN => \N__80482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29354\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80475\,
            DIN => \N__80474\,
            DOUT => \N__80473\,
            PACKAGEPIN => \OE_wire\
        );

    \OE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80475\,
            PADOUT => \N__80474\,
            PADIN => \N__80473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25703\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80466\,
            DIN => \N__80465\,
            DOUT => \N__80464\,
            PACKAGEPIN => \GPIO3_wire\
        );

    \GPIO3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80466\,
            PADOUT => \N__80465\,
            PADIN => \N__80464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25811\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80457\,
            DIN => \N__80456\,
            DOUT => \N__80455\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(10)
        );

    \BUFFER_ADDRESS_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80457\,
            PADOUT => \N__80456\,
            PADIN => \N__80455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26510\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D2_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80448\,
            DIN => \N__80447\,
            DOUT => \N__80446\,
            PACKAGEPIN => \D2_in_wire\
        );

    \D2_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80448\,
            PADOUT => \N__80447\,
            PADIN => \N__80446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D2_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80439\,
            DIN => \N__80438\,
            DOUT => \N__80437\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(11)
        );

    \BUFFER_DATA_IN_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80439\,
            PADOUT => \N__80438\,
            PADIN => \N__80437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A14_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80430\,
            DIN => \N__80429\,
            DOUT => \N__80428\,
            PACKAGEPIN => \A14_wire\
        );

    \A14_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80430\,
            PADOUT => \N__80429\,
            PADIN => \N__80428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__44111\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A5_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80421\,
            DIN => \N__80420\,
            DOUT => \N__80419\,
            PACKAGEPIN => \A5_wire\
        );

    \A5_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80421\,
            PADOUT => \N__80420\,
            PADIN => \N__80419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80412\,
            DIN => \N__80411\,
            DOUT => \N__80410\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(3)
        );

    \BUFFER_DATA_OUT_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80412\,
            PADOUT => \N__80411\,
            PADIN => \N__80410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80403\,
            DIN => \N__80402\,
            DOUT => \N__80401\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(1)
        );

    \BUFFER_DATA_IN_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80403\,
            PADOUT => \N__80402\,
            PADIN => \N__80401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D9_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80394\,
            DIN => \N__80393\,
            DOUT => \N__80392\,
            PACKAGEPIN => \D9_wire\
        );

    \D9_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80394\,
            PADOUT => \N__80393\,
            PADIN => \N__80392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35097\,
            DIN0 => OPEN,
            DOUT0 => \N__40384\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80385\,
            DIN => \N__80384\,
            DOUT => \N__80383\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(1)
        );

    \BUFFER_ADDRESS_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80385\,
            PADOUT => \N__80384\,
            PADIN => \N__80383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26159\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D11_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80376\,
            DIN => \N__80375\,
            DOUT => \N__80374\,
            PACKAGEPIN => \D11_wire\
        );

    \D11_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80376\,
            PADOUT => \N__80375\,
            PADIN => \N__80374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35098\,
            DIN0 => OPEN,
            DOUT0 => \N__37358\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D12_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80367\,
            DIN => \N__80366\,
            DOUT => \N__80365\,
            PACKAGEPIN => \D12_in_wire\
        );

    \D12_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80367\,
            PADOUT => \N__80366\,
            PADIN => \N__80365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D12_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A15_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80358\,
            DIN => \N__80357\,
            DOUT => \N__80356\,
            PACKAGEPIN => \A15_wire\
        );

    \A15_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80358\,
            PADOUT => \N__80357\,
            PADIN => \N__80356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__44978\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A13_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80349\,
            DIN => \N__80348\,
            DOUT => \N__80347\,
            PACKAGEPIN => \A13_wire\
        );

    \A13_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80349\,
            PADOUT => \N__80348\,
            PADIN => \N__80347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28175\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80340\,
            DIN => \N__80339\,
            DOUT => \N__80338\,
            PACKAGEPIN => \A1_wire\
        );

    \A1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80340\,
            PADOUT => \N__80339\,
            PADIN => \N__80338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31310\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80331\,
            DIN => \N__80330\,
            DOUT => \N__80329\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(10)
        );

    \BUFFER_DATA_OUT_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80331\,
            PADOUT => \N__80330\,
            PADIN => \N__80329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26224\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_UB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80322\,
            DIN => \N__80321\,
            DOUT => \N__80320\,
            PACKAGEPIN => \B_UB_wire\
        );

    \B_UB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80322\,
            PADOUT => \N__80321\,
            PADIN => \N__80320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25792\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D7_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80313\,
            DIN => \N__80312\,
            DOUT => \N__80311\,
            PACKAGEPIN => \D7_in_wire\
        );

    \D7_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80313\,
            PADOUT => \N__80312\,
            PADIN => \N__80311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D7_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_WR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80304\,
            DIN => \N__80303\,
            DOUT => \N__80302\,
            PACKAGEPIN => \B_WR_wire\
        );

    \B_WR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80304\,
            PADOUT => \N__80303\,
            PADIN => \N__80302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25793\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80295\,
            DIN => \N__80294\,
            DOUT => \N__80293\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(14)
        );

    \BUFFER_DATA_IN_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80295\,
            PADOUT => \N__80294\,
            PADIN => \N__80293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80286\,
            DIN => \N__80285\,
            DOUT => \N__80284\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(11)
        );

    \BUFFER_ADDRESS_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80286\,
            PADOUT => \N__80285\,
            PADIN => \N__80284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25748\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO11_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80277\,
            DIN => \N__80276\,
            DOUT => \N__80275\,
            PACKAGEPIN => \GPIO11_wire\
        );

    \GPIO11_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80277\,
            PADOUT => \N__80276\,
            PADIN => \N__80275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80268\,
            DIN => \N__80267\,
            DOUT => \N__80266\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(6)
        );

    \BUFFER_DATA_OUT_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80268\,
            PADOUT => \N__80267\,
            PADIN => \N__80266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__63370\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80259\,
            DIN => \N__80258\,
            DOUT => \N__80257\,
            PACKAGEPIN => \A2_wire\
        );

    \A2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80259\,
            PADOUT => \N__80258\,
            PADIN => \N__80257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29576\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D5_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80250\,
            DIN => \N__80249\,
            DOUT => \N__80248\,
            PACKAGEPIN => \D5_wire\
        );

    \D5_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80250\,
            PADOUT => \N__80249\,
            PADIN => \N__80248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35052\,
            DIN0 => OPEN,
            DOUT0 => \N__52541\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D4_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80241\,
            DIN => \N__80240\,
            DOUT => \N__80239\,
            PACKAGEPIN => \D4_wire\
        );

    \D4_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80241\,
            PADOUT => \N__80240\,
            PADIN => \N__80239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35101\,
            DIN0 => OPEN,
            DOUT0 => \N__33764\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80232\,
            DIN => \N__80231\,
            DOUT => \N__80230\,
            PACKAGEPIN => \A3_wire\
        );

    \A3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80232\,
            PADOUT => \N__80231\,
            PADIN => \N__80230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__44048\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80223\,
            DIN => \N__80222\,
            DOUT => \N__80221\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(0)
        );

    \BUFFER_DATA_OUT_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80223\,
            PADOUT => \N__80222\,
            PADIN => \N__80221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37684\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80214\,
            DIN => \N__80213\,
            DOUT => \N__80212\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(0)
        );

    \BUFFER_DATA_IN_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80214\,
            PADOUT => \N__80213\,
            PADIN => \N__80212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80205\,
            DIN => \N__80204\,
            DOUT => \N__80203\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(0)
        );

    \BUFFER_ADDRESS_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80205\,
            PADOUT => \N__80204\,
            PADIN => \N__80203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26177\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80196\,
            DIN => \N__80195\,
            DOUT => \N__80194\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(15)
        );

    \BUFFER_DATA_OUT_obuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80196\,
            PADOUT => \N__80195\,
            PADIN => \N__80194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__49232\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A11_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80187\,
            DIN => \N__80186\,
            DOUT => \N__80185\,
            PACKAGEPIN => \A11_wire\
        );

    \A11_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80187\,
            PADOUT => \N__80186\,
            PADIN => \N__80185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31181\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO9_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80178\,
            DIN => \N__80177\,
            DOUT => \N__80176\,
            PACKAGEPIN => \GPIO9_wire\
        );

    \GPIO9_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80178\,
            PADOUT => \N__80177\,
            PADIN => \N__80176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32573\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D5_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80169\,
            DIN => \N__80168\,
            DOUT => \N__80167\,
            PACKAGEPIN => \D5_in_wire\
        );

    \D5_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80169\,
            PADOUT => \N__80168\,
            PADIN => \N__80167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D5_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80160\,
            DIN => \N__80159\,
            DOUT => \N__80158\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(14)
        );

    \BUFFER_ADDRESS_obuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80160\,
            PADOUT => \N__80159\,
            PADIN => \N__80158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25733\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D15_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80151\,
            DIN => \N__80150\,
            DOUT => \N__80149\,
            PACKAGEPIN => \D15_in_wire\
        );

    \D15_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80151\,
            PADOUT => \N__80150\,
            PADIN => \N__80149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D15_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D1_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80142\,
            DIN => \N__80141\,
            DOUT => \N__80140\,
            PACKAGEPIN => \D1_in_wire\
        );

    \D1_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80142\,
            PADOUT => \N__80141\,
            PADIN => \N__80140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D1_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \B_OE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80133\,
            DIN => \N__80132\,
            DOUT => \N__80131\,
            PACKAGEPIN => \B_OE_wire\
        );

    \B_OE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80133\,
            PADOUT => \N__80132\,
            PADIN => \N__80131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25775\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80124\,
            DIN => \N__80123\,
            DOUT => \N__80122\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(15)
        );

    \BUFFER_DATA_IN_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80124\,
            PADOUT => \N__80123\,
            PADIN => \N__80122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80115\,
            DIN => \N__80114\,
            DOUT => \N__80113\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(7)
        );

    \BUFFER_DATA_OUT_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80115\,
            PADOUT => \N__80114\,
            PADIN => \N__80113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__46039\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80106\,
            DIN => \N__80105\,
            DOUT => \N__80104\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(5)
        );

    \BUFFER_DATA_IN_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80106\,
            PADOUT => \N__80105\,
            PADIN => \N__80104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D12_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80097\,
            DIN => \N__80096\,
            DOUT => \N__80095\,
            PACKAGEPIN => \D12_wire\
        );

    \D12_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80097\,
            PADOUT => \N__80096\,
            PADIN => \N__80095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35051\,
            DIN0 => OPEN,
            DOUT0 => \N__26327\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80088\,
            DIN => \N__80087\,
            DOUT => \N__80086\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(5)
        );

    \BUFFER_ADDRESS_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80088\,
            PADOUT => \N__80087\,
            PADIN => \N__80086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29288\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TX_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80079\,
            DIN => \N__80078\,
            DOUT => \N__80077\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__80079\,
            PADOUT => \N__80078\,
            PADIN => \N__80077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D8_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80070\,
            DIN => \N__80069\,
            DOUT => \N__80068\,
            PACKAGEPIN => \D8_in_wire\
        );

    \D8_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80070\,
            PADOUT => \N__80069\,
            PADIN => \N__80068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D8_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80061\,
            DIN => \N__80060\,
            DOUT => \N__80059\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(1)
        );

    \BUFFER_DATA_OUT_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80061\,
            PADOUT => \N__80060\,
            PADIN => \N__80059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__69070\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D6_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80052\,
            DIN => \N__80051\,
            DOUT => \N__80050\,
            PACKAGEPIN => \D6_in_wire\
        );

    \D6_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80052\,
            PADOUT => \N__80051\,
            PADIN => \N__80050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D6_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80043\,
            DIN => \N__80042\,
            DOUT => \N__80041\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(3)
        );

    \BUFFER_DATA_IN_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80043\,
            PADOUT => \N__80042\,
            PADIN => \N__80041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D13_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80034\,
            DIN => \N__80033\,
            DOUT => \N__80032\,
            PACKAGEPIN => \D13_in_wire\
        );

    \D13_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80034\,
            PADOUT => \N__80033\,
            PADIN => \N__80032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \D13_in_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80025\,
            DIN => \N__80024\,
            DOUT => \N__80023\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(3)
        );

    \BUFFER_ADDRESS_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80025\,
            PADOUT => \N__80024\,
            PADIN => \N__80023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29333\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80016\,
            DIN => \N__80015\,
            DOUT => \N__80014\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(14)
        );

    \BUFFER_DATA_OUT_obuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__80016\,
            PADOUT => \N__80015\,
            PADIN => \N__80014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__39752\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__80007\,
            DIN => \N__80006\,
            DOUT => \N__80005\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(9)
        );

    \BUFFER_DATA_IN_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__80007\,
            PADOUT => \N__80006\,
            PADIN => \N__80005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79998\,
            DIN => \N__79997\,
            DOUT => \N__79996\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(9)
        );

    \BUFFER_ADDRESS_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__79998\,
            PADOUT => \N__79997\,
            PADIN => \N__79996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25715\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D1_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79989\,
            DIN => \N__79988\,
            DOUT => \N__79987\,
            PACKAGEPIN => \D1_wire\
        );

    \D1_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__79989\,
            PADOUT => \N__79988\,
            PADIN => \N__79987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35112\,
            DIN0 => OPEN,
            DOUT0 => \N__69074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79980\,
            DIN => \N__79979\,
            DOUT => \N__79978\,
            PACKAGEPIN => \A12_wire\
        );

    \A12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__79980\,
            PADOUT => \N__79979\,
            PADIN => \N__79978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_OUT_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79971\,
            DIN => \N__79970\,
            DOUT => \N__79969\,
            PACKAGEPIN => \BUFFER_DATA_OUT_wire\(4)
        );

    \BUFFER_DATA_OUT_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__79971\,
            PADOUT => \N__79970\,
            PADIN => \N__79969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33763\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_DATA_IN_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79962\,
            DIN => \N__79961\,
            DOUT => \N__79960\,
            PACKAGEPIN => \BUFFER_DATA_IN_wire\(4)
        );

    \BUFFER_DATA_IN_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__79962\,
            PADOUT => \N__79961\,
            PADIN => \N__79960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \gpuOut_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79953\,
            DIN => \N__79952\,
            DOUT => \N__79951\,
            PACKAGEPIN => \A0_wire\
        );

    \A0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__79953\,
            PADOUT => \N__79952\,
            PADIN => \N__79951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31334\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79944\,
            DIN => \N__79943\,
            DOUT => \N__79942\,
            PACKAGEPIN => \CE_wire\
        );

    \CE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__79944\,
            PADOUT => \N__79943\,
            PADIN => \N__79942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32494\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D14_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79935\,
            DIN => \N__79934\,
            DOUT => \N__79933\,
            PACKAGEPIN => \D14_wire\
        );

    \D14_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__79935\,
            PADOUT => \N__79934\,
            PADIN => \N__79933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__35026\,
            DIN0 => OPEN,
            DOUT0 => \N__39751\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFFER_ADDRESS_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__79926\,
            DIN => \N__79925\,
            DOUT => \N__79924\,
            PACKAGEPIN => \BUFFER_ADDRESS_wire\(2)
        );

    \BUFFER_ADDRESS_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__79926\,
            PADOUT => \N__79925\,
            PADIN => \N__79924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29108\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__20304\ : InMux
    port map (
            O => \N__79907\,
            I => \N__79904\
        );

    \I__20303\ : LocalMux
    port map (
            O => \N__79904\,
            I => \N__79901\
        );

    \I__20302\ : Odrv4
    port map (
            O => \N__79901\,
            I => \PROM.ROMDATA.m331_ns\
        );

    \I__20301\ : InMux
    port map (
            O => \N__79898\,
            I => \N__79892\
        );

    \I__20300\ : InMux
    port map (
            O => \N__79897\,
            I => \N__79887\
        );

    \I__20299\ : InMux
    port map (
            O => \N__79896\,
            I => \N__79884\
        );

    \I__20298\ : InMux
    port map (
            O => \N__79895\,
            I => \N__79875\
        );

    \I__20297\ : LocalMux
    port map (
            O => \N__79892\,
            I => \N__79867\
        );

    \I__20296\ : CascadeMux
    port map (
            O => \N__79891\,
            I => \N__79863\
        );

    \I__20295\ : CascadeMux
    port map (
            O => \N__79890\,
            I => \N__79854\
        );

    \I__20294\ : LocalMux
    port map (
            O => \N__79887\,
            I => \N__79851\
        );

    \I__20293\ : LocalMux
    port map (
            O => \N__79884\,
            I => \N__79847\
        );

    \I__20292\ : InMux
    port map (
            O => \N__79883\,
            I => \N__79835\
        );

    \I__20291\ : InMux
    port map (
            O => \N__79882\,
            I => \N__79819\
        );

    \I__20290\ : InMux
    port map (
            O => \N__79881\,
            I => \N__79819\
        );

    \I__20289\ : InMux
    port map (
            O => \N__79880\,
            I => \N__79819\
        );

    \I__20288\ : InMux
    port map (
            O => \N__79879\,
            I => \N__79819\
        );

    \I__20287\ : InMux
    port map (
            O => \N__79878\,
            I => \N__79819\
        );

    \I__20286\ : LocalMux
    port map (
            O => \N__79875\,
            I => \N__79815\
        );

    \I__20285\ : InMux
    port map (
            O => \N__79874\,
            I => \N__79812\
        );

    \I__20284\ : InMux
    port map (
            O => \N__79873\,
            I => \N__79809\
        );

    \I__20283\ : InMux
    port map (
            O => \N__79872\,
            I => \N__79801\
        );

    \I__20282\ : InMux
    port map (
            O => \N__79871\,
            I => \N__79801\
        );

    \I__20281\ : InMux
    port map (
            O => \N__79870\,
            I => \N__79801\
        );

    \I__20280\ : Span4Mux_v
    port map (
            O => \N__79867\,
            I => \N__79798\
        );

    \I__20279\ : InMux
    port map (
            O => \N__79866\,
            I => \N__79795\
        );

    \I__20278\ : InMux
    port map (
            O => \N__79863\,
            I => \N__79792\
        );

    \I__20277\ : InMux
    port map (
            O => \N__79862\,
            I => \N__79789\
        );

    \I__20276\ : CascadeMux
    port map (
            O => \N__79861\,
            I => \N__79784\
        );

    \I__20275\ : InMux
    port map (
            O => \N__79860\,
            I => \N__79778\
        );

    \I__20274\ : InMux
    port map (
            O => \N__79859\,
            I => \N__79778\
        );

    \I__20273\ : InMux
    port map (
            O => \N__79858\,
            I => \N__79775\
        );

    \I__20272\ : InMux
    port map (
            O => \N__79857\,
            I => \N__79772\
        );

    \I__20271\ : InMux
    port map (
            O => \N__79854\,
            I => \N__79769\
        );

    \I__20270\ : Span4Mux_v
    port map (
            O => \N__79851\,
            I => \N__79766\
        );

    \I__20269\ : InMux
    port map (
            O => \N__79850\,
            I => \N__79763\
        );

    \I__20268\ : Span4Mux_v
    port map (
            O => \N__79847\,
            I => \N__79758\
        );

    \I__20267\ : InMux
    port map (
            O => \N__79846\,
            I => \N__79755\
        );

    \I__20266\ : InMux
    port map (
            O => \N__79845\,
            I => \N__79752\
        );

    \I__20265\ : InMux
    port map (
            O => \N__79844\,
            I => \N__79748\
        );

    \I__20264\ : InMux
    port map (
            O => \N__79843\,
            I => \N__79744\
        );

    \I__20263\ : InMux
    port map (
            O => \N__79842\,
            I => \N__79741\
        );

    \I__20262\ : InMux
    port map (
            O => \N__79841\,
            I => \N__79738\
        );

    \I__20261\ : InMux
    port map (
            O => \N__79840\,
            I => \N__79735\
        );

    \I__20260\ : InMux
    port map (
            O => \N__79839\,
            I => \N__79732\
        );

    \I__20259\ : InMux
    port map (
            O => \N__79838\,
            I => \N__79729\
        );

    \I__20258\ : LocalMux
    port map (
            O => \N__79835\,
            I => \N__79726\
        );

    \I__20257\ : InMux
    port map (
            O => \N__79834\,
            I => \N__79723\
        );

    \I__20256\ : InMux
    port map (
            O => \N__79833\,
            I => \N__79716\
        );

    \I__20255\ : InMux
    port map (
            O => \N__79832\,
            I => \N__79716\
        );

    \I__20254\ : InMux
    port map (
            O => \N__79831\,
            I => \N__79716\
        );

    \I__20253\ : CascadeMux
    port map (
            O => \N__79830\,
            I => \N__79711\
        );

    \I__20252\ : LocalMux
    port map (
            O => \N__79819\,
            I => \N__79708\
        );

    \I__20251\ : InMux
    port map (
            O => \N__79818\,
            I => \N__79705\
        );

    \I__20250\ : Span4Mux_v
    port map (
            O => \N__79815\,
            I => \N__79698\
        );

    \I__20249\ : LocalMux
    port map (
            O => \N__79812\,
            I => \N__79698\
        );

    \I__20248\ : LocalMux
    port map (
            O => \N__79809\,
            I => \N__79698\
        );

    \I__20247\ : InMux
    port map (
            O => \N__79808\,
            I => \N__79695\
        );

    \I__20246\ : LocalMux
    port map (
            O => \N__79801\,
            I => \N__79692\
        );

    \I__20245\ : Sp12to4
    port map (
            O => \N__79798\,
            I => \N__79683\
        );

    \I__20244\ : LocalMux
    port map (
            O => \N__79795\,
            I => \N__79683\
        );

    \I__20243\ : LocalMux
    port map (
            O => \N__79792\,
            I => \N__79683\
        );

    \I__20242\ : LocalMux
    port map (
            O => \N__79789\,
            I => \N__79683\
        );

    \I__20241\ : InMux
    port map (
            O => \N__79788\,
            I => \N__79678\
        );

    \I__20240\ : InMux
    port map (
            O => \N__79787\,
            I => \N__79678\
        );

    \I__20239\ : InMux
    port map (
            O => \N__79784\,
            I => \N__79675\
        );

    \I__20238\ : InMux
    port map (
            O => \N__79783\,
            I => \N__79672\
        );

    \I__20237\ : LocalMux
    port map (
            O => \N__79778\,
            I => \N__79667\
        );

    \I__20236\ : LocalMux
    port map (
            O => \N__79775\,
            I => \N__79667\
        );

    \I__20235\ : LocalMux
    port map (
            O => \N__79772\,
            I => \N__79662\
        );

    \I__20234\ : LocalMux
    port map (
            O => \N__79769\,
            I => \N__79662\
        );

    \I__20233\ : Span4Mux_h
    port map (
            O => \N__79766\,
            I => \N__79657\
        );

    \I__20232\ : LocalMux
    port map (
            O => \N__79763\,
            I => \N__79657\
        );

    \I__20231\ : InMux
    port map (
            O => \N__79762\,
            I => \N__79652\
        );

    \I__20230\ : InMux
    port map (
            O => \N__79761\,
            I => \N__79652\
        );

    \I__20229\ : Span4Mux_h
    port map (
            O => \N__79758\,
            I => \N__79649\
        );

    \I__20228\ : LocalMux
    port map (
            O => \N__79755\,
            I => \N__79644\
        );

    \I__20227\ : LocalMux
    port map (
            O => \N__79752\,
            I => \N__79644\
        );

    \I__20226\ : InMux
    port map (
            O => \N__79751\,
            I => \N__79641\
        );

    \I__20225\ : LocalMux
    port map (
            O => \N__79748\,
            I => \N__79638\
        );

    \I__20224\ : InMux
    port map (
            O => \N__79747\,
            I => \N__79635\
        );

    \I__20223\ : LocalMux
    port map (
            O => \N__79744\,
            I => \N__79628\
        );

    \I__20222\ : LocalMux
    port map (
            O => \N__79741\,
            I => \N__79628\
        );

    \I__20221\ : LocalMux
    port map (
            O => \N__79738\,
            I => \N__79628\
        );

    \I__20220\ : LocalMux
    port map (
            O => \N__79735\,
            I => \N__79621\
        );

    \I__20219\ : LocalMux
    port map (
            O => \N__79732\,
            I => \N__79621\
        );

    \I__20218\ : LocalMux
    port map (
            O => \N__79729\,
            I => \N__79621\
        );

    \I__20217\ : Span4Mux_v
    port map (
            O => \N__79726\,
            I => \N__79614\
        );

    \I__20216\ : LocalMux
    port map (
            O => \N__79723\,
            I => \N__79614\
        );

    \I__20215\ : LocalMux
    port map (
            O => \N__79716\,
            I => \N__79614\
        );

    \I__20214\ : InMux
    port map (
            O => \N__79715\,
            I => \N__79610\
        );

    \I__20213\ : InMux
    port map (
            O => \N__79714\,
            I => \N__79605\
        );

    \I__20212\ : InMux
    port map (
            O => \N__79711\,
            I => \N__79605\
        );

    \I__20211\ : Span4Mux_v
    port map (
            O => \N__79708\,
            I => \N__79598\
        );

    \I__20210\ : LocalMux
    port map (
            O => \N__79705\,
            I => \N__79598\
        );

    \I__20209\ : Span4Mux_h
    port map (
            O => \N__79698\,
            I => \N__79598\
        );

    \I__20208\ : LocalMux
    port map (
            O => \N__79695\,
            I => \N__79591\
        );

    \I__20207\ : Span12Mux_h
    port map (
            O => \N__79692\,
            I => \N__79591\
        );

    \I__20206\ : Span12Mux_h
    port map (
            O => \N__79683\,
            I => \N__79591\
        );

    \I__20205\ : LocalMux
    port map (
            O => \N__79678\,
            I => \N__79584\
        );

    \I__20204\ : LocalMux
    port map (
            O => \N__79675\,
            I => \N__79584\
        );

    \I__20203\ : LocalMux
    port map (
            O => \N__79672\,
            I => \N__79584\
        );

    \I__20202\ : Span12Mux_s11_v
    port map (
            O => \N__79667\,
            I => \N__79581\
        );

    \I__20201\ : Span4Mux_v
    port map (
            O => \N__79662\,
            I => \N__79578\
        );

    \I__20200\ : Span4Mux_v
    port map (
            O => \N__79657\,
            I => \N__79573\
        );

    \I__20199\ : LocalMux
    port map (
            O => \N__79652\,
            I => \N__79573\
        );

    \I__20198\ : Span4Mux_h
    port map (
            O => \N__79649\,
            I => \N__79556\
        );

    \I__20197\ : Span4Mux_v
    port map (
            O => \N__79644\,
            I => \N__79556\
        );

    \I__20196\ : LocalMux
    port map (
            O => \N__79641\,
            I => \N__79556\
        );

    \I__20195\ : Span4Mux_v
    port map (
            O => \N__79638\,
            I => \N__79556\
        );

    \I__20194\ : LocalMux
    port map (
            O => \N__79635\,
            I => \N__79556\
        );

    \I__20193\ : Span4Mux_v
    port map (
            O => \N__79628\,
            I => \N__79556\
        );

    \I__20192\ : Span4Mux_v
    port map (
            O => \N__79621\,
            I => \N__79556\
        );

    \I__20191\ : Span4Mux_h
    port map (
            O => \N__79614\,
            I => \N__79556\
        );

    \I__20190\ : InMux
    port map (
            O => \N__79613\,
            I => \N__79553\
        );

    \I__20189\ : LocalMux
    port map (
            O => \N__79610\,
            I => \progRomAddress_5\
        );

    \I__20188\ : LocalMux
    port map (
            O => \N__79605\,
            I => \progRomAddress_5\
        );

    \I__20187\ : Odrv4
    port map (
            O => \N__79598\,
            I => \progRomAddress_5\
        );

    \I__20186\ : Odrv12
    port map (
            O => \N__79591\,
            I => \progRomAddress_5\
        );

    \I__20185\ : Odrv4
    port map (
            O => \N__79584\,
            I => \progRomAddress_5\
        );

    \I__20184\ : Odrv12
    port map (
            O => \N__79581\,
            I => \progRomAddress_5\
        );

    \I__20183\ : Odrv4
    port map (
            O => \N__79578\,
            I => \progRomAddress_5\
        );

    \I__20182\ : Odrv4
    port map (
            O => \N__79573\,
            I => \progRomAddress_5\
        );

    \I__20181\ : Odrv4
    port map (
            O => \N__79556\,
            I => \progRomAddress_5\
        );

    \I__20180\ : LocalMux
    port map (
            O => \N__79553\,
            I => \progRomAddress_5\
        );

    \I__20179\ : CascadeMux
    port map (
            O => \N__79532\,
            I => \N__79524\
        );

    \I__20178\ : CascadeMux
    port map (
            O => \N__79531\,
            I => \N__79519\
        );

    \I__20177\ : CascadeMux
    port map (
            O => \N__79530\,
            I => \N__79516\
        );

    \I__20176\ : CascadeMux
    port map (
            O => \N__79529\,
            I => \N__79511\
        );

    \I__20175\ : CascadeMux
    port map (
            O => \N__79528\,
            I => \N__79508\
        );

    \I__20174\ : CascadeMux
    port map (
            O => \N__79527\,
            I => \N__79504\
        );

    \I__20173\ : InMux
    port map (
            O => \N__79524\,
            I => \N__79490\
        );

    \I__20172\ : InMux
    port map (
            O => \N__79523\,
            I => \N__79490\
        );

    \I__20171\ : InMux
    port map (
            O => \N__79522\,
            I => \N__79483\
        );

    \I__20170\ : InMux
    port map (
            O => \N__79519\,
            I => \N__79474\
        );

    \I__20169\ : InMux
    port map (
            O => \N__79516\,
            I => \N__79474\
        );

    \I__20168\ : InMux
    port map (
            O => \N__79515\,
            I => \N__79474\
        );

    \I__20167\ : InMux
    port map (
            O => \N__79514\,
            I => \N__79474\
        );

    \I__20166\ : InMux
    port map (
            O => \N__79511\,
            I => \N__79469\
        );

    \I__20165\ : InMux
    port map (
            O => \N__79508\,
            I => \N__79469\
        );

    \I__20164\ : InMux
    port map (
            O => \N__79507\,
            I => \N__79464\
        );

    \I__20163\ : InMux
    port map (
            O => \N__79504\,
            I => \N__79464\
        );

    \I__20162\ : InMux
    port map (
            O => \N__79503\,
            I => \N__79461\
        );

    \I__20161\ : InMux
    port map (
            O => \N__79502\,
            I => \N__79458\
        );

    \I__20160\ : InMux
    port map (
            O => \N__79501\,
            I => \N__79447\
        );

    \I__20159\ : InMux
    port map (
            O => \N__79500\,
            I => \N__79447\
        );

    \I__20158\ : InMux
    port map (
            O => \N__79499\,
            I => \N__79440\
        );

    \I__20157\ : InMux
    port map (
            O => \N__79498\,
            I => \N__79440\
        );

    \I__20156\ : InMux
    port map (
            O => \N__79497\,
            I => \N__79440\
        );

    \I__20155\ : CascadeMux
    port map (
            O => \N__79496\,
            I => \N__79437\
        );

    \I__20154\ : CascadeMux
    port map (
            O => \N__79495\,
            I => \N__79434\
        );

    \I__20153\ : LocalMux
    port map (
            O => \N__79490\,
            I => \N__79428\
        );

    \I__20152\ : CascadeMux
    port map (
            O => \N__79489\,
            I => \N__79425\
        );

    \I__20151\ : CascadeMux
    port map (
            O => \N__79488\,
            I => \N__79422\
        );

    \I__20150\ : InMux
    port map (
            O => \N__79487\,
            I => \N__79408\
        );

    \I__20149\ : InMux
    port map (
            O => \N__79486\,
            I => \N__79405\
        );

    \I__20148\ : LocalMux
    port map (
            O => \N__79483\,
            I => \N__79398\
        );

    \I__20147\ : LocalMux
    port map (
            O => \N__79474\,
            I => \N__79398\
        );

    \I__20146\ : LocalMux
    port map (
            O => \N__79469\,
            I => \N__79398\
        );

    \I__20145\ : LocalMux
    port map (
            O => \N__79464\,
            I => \N__79395\
        );

    \I__20144\ : LocalMux
    port map (
            O => \N__79461\,
            I => \N__79392\
        );

    \I__20143\ : LocalMux
    port map (
            O => \N__79458\,
            I => \N__79388\
        );

    \I__20142\ : InMux
    port map (
            O => \N__79457\,
            I => \N__79381\
        );

    \I__20141\ : InMux
    port map (
            O => \N__79456\,
            I => \N__79381\
        );

    \I__20140\ : InMux
    port map (
            O => \N__79455\,
            I => \N__79381\
        );

    \I__20139\ : InMux
    port map (
            O => \N__79454\,
            I => \N__79378\
        );

    \I__20138\ : InMux
    port map (
            O => \N__79453\,
            I => \N__79373\
        );

    \I__20137\ : InMux
    port map (
            O => \N__79452\,
            I => \N__79373\
        );

    \I__20136\ : LocalMux
    port map (
            O => \N__79447\,
            I => \N__79370\
        );

    \I__20135\ : LocalMux
    port map (
            O => \N__79440\,
            I => \N__79367\
        );

    \I__20134\ : InMux
    port map (
            O => \N__79437\,
            I => \N__79358\
        );

    \I__20133\ : InMux
    port map (
            O => \N__79434\,
            I => \N__79358\
        );

    \I__20132\ : InMux
    port map (
            O => \N__79433\,
            I => \N__79358\
        );

    \I__20131\ : InMux
    port map (
            O => \N__79432\,
            I => \N__79358\
        );

    \I__20130\ : InMux
    port map (
            O => \N__79431\,
            I => \N__79355\
        );

    \I__20129\ : Span4Mux_v
    port map (
            O => \N__79428\,
            I => \N__79352\
        );

    \I__20128\ : InMux
    port map (
            O => \N__79425\,
            I => \N__79343\
        );

    \I__20127\ : InMux
    port map (
            O => \N__79422\,
            I => \N__79343\
        );

    \I__20126\ : InMux
    port map (
            O => \N__79421\,
            I => \N__79343\
        );

    \I__20125\ : InMux
    port map (
            O => \N__79420\,
            I => \N__79343\
        );

    \I__20124\ : InMux
    port map (
            O => \N__79419\,
            I => \N__79336\
        );

    \I__20123\ : InMux
    port map (
            O => \N__79418\,
            I => \N__79336\
        );

    \I__20122\ : CascadeMux
    port map (
            O => \N__79417\,
            I => \N__79333\
        );

    \I__20121\ : InMux
    port map (
            O => \N__79416\,
            I => \N__79328\
        );

    \I__20120\ : InMux
    port map (
            O => \N__79415\,
            I => \N__79328\
        );

    \I__20119\ : CascadeMux
    port map (
            O => \N__79414\,
            I => \N__79324\
        );

    \I__20118\ : CascadeMux
    port map (
            O => \N__79413\,
            I => \N__79315\
        );

    \I__20117\ : InMux
    port map (
            O => \N__79412\,
            I => \N__79309\
        );

    \I__20116\ : InMux
    port map (
            O => \N__79411\,
            I => \N__79309\
        );

    \I__20115\ : LocalMux
    port map (
            O => \N__79408\,
            I => \N__79306\
        );

    \I__20114\ : LocalMux
    port map (
            O => \N__79405\,
            I => \N__79301\
        );

    \I__20113\ : Span4Mux_v
    port map (
            O => \N__79398\,
            I => \N__79301\
        );

    \I__20112\ : Span4Mux_v
    port map (
            O => \N__79395\,
            I => \N__79294\
        );

    \I__20111\ : Span4Mux_v
    port map (
            O => \N__79392\,
            I => \N__79290\
        );

    \I__20110\ : InMux
    port map (
            O => \N__79391\,
            I => \N__79287\
        );

    \I__20109\ : Span4Mux_h
    port map (
            O => \N__79388\,
            I => \N__79277\
        );

    \I__20108\ : LocalMux
    port map (
            O => \N__79381\,
            I => \N__79277\
        );

    \I__20107\ : LocalMux
    port map (
            O => \N__79378\,
            I => \N__79277\
        );

    \I__20106\ : LocalMux
    port map (
            O => \N__79373\,
            I => \N__79277\
        );

    \I__20105\ : Span4Mux_v
    port map (
            O => \N__79370\,
            I => \N__79274\
        );

    \I__20104\ : Span4Mux_h
    port map (
            O => \N__79367\,
            I => \N__79269\
        );

    \I__20103\ : LocalMux
    port map (
            O => \N__79358\,
            I => \N__79269\
        );

    \I__20102\ : LocalMux
    port map (
            O => \N__79355\,
            I => \N__79262\
        );

    \I__20101\ : Span4Mux_h
    port map (
            O => \N__79352\,
            I => \N__79262\
        );

    \I__20100\ : LocalMux
    port map (
            O => \N__79343\,
            I => \N__79262\
        );

    \I__20099\ : InMux
    port map (
            O => \N__79342\,
            I => \N__79259\
        );

    \I__20098\ : InMux
    port map (
            O => \N__79341\,
            I => \N__79256\
        );

    \I__20097\ : LocalMux
    port map (
            O => \N__79336\,
            I => \N__79253\
        );

    \I__20096\ : InMux
    port map (
            O => \N__79333\,
            I => \N__79250\
        );

    \I__20095\ : LocalMux
    port map (
            O => \N__79328\,
            I => \N__79245\
        );

    \I__20094\ : InMux
    port map (
            O => \N__79327\,
            I => \N__79238\
        );

    \I__20093\ : InMux
    port map (
            O => \N__79324\,
            I => \N__79238\
        );

    \I__20092\ : InMux
    port map (
            O => \N__79323\,
            I => \N__79238\
        );

    \I__20091\ : InMux
    port map (
            O => \N__79322\,
            I => \N__79233\
        );

    \I__20090\ : InMux
    port map (
            O => \N__79321\,
            I => \N__79233\
        );

    \I__20089\ : InMux
    port map (
            O => \N__79320\,
            I => \N__79228\
        );

    \I__20088\ : InMux
    port map (
            O => \N__79319\,
            I => \N__79228\
        );

    \I__20087\ : InMux
    port map (
            O => \N__79318\,
            I => \N__79223\
        );

    \I__20086\ : InMux
    port map (
            O => \N__79315\,
            I => \N__79223\
        );

    \I__20085\ : InMux
    port map (
            O => \N__79314\,
            I => \N__79220\
        );

    \I__20084\ : LocalMux
    port map (
            O => \N__79309\,
            I => \N__79217\
        );

    \I__20083\ : Span4Mux_v
    port map (
            O => \N__79306\,
            I => \N__79214\
        );

    \I__20082\ : Span4Mux_h
    port map (
            O => \N__79301\,
            I => \N__79211\
        );

    \I__20081\ : InMux
    port map (
            O => \N__79300\,
            I => \N__79204\
        );

    \I__20080\ : InMux
    port map (
            O => \N__79299\,
            I => \N__79201\
        );

    \I__20079\ : InMux
    port map (
            O => \N__79298\,
            I => \N__79196\
        );

    \I__20078\ : InMux
    port map (
            O => \N__79297\,
            I => \N__79196\
        );

    \I__20077\ : Span4Mux_h
    port map (
            O => \N__79294\,
            I => \N__79193\
        );

    \I__20076\ : InMux
    port map (
            O => \N__79293\,
            I => \N__79190\
        );

    \I__20075\ : Span4Mux_h
    port map (
            O => \N__79290\,
            I => \N__79185\
        );

    \I__20074\ : LocalMux
    port map (
            O => \N__79287\,
            I => \N__79185\
        );

    \I__20073\ : InMux
    port map (
            O => \N__79286\,
            I => \N__79182\
        );

    \I__20072\ : Span4Mux_v
    port map (
            O => \N__79277\,
            I => \N__79179\
        );

    \I__20071\ : Span4Mux_h
    port map (
            O => \N__79274\,
            I => \N__79176\
        );

    \I__20070\ : Span4Mux_h
    port map (
            O => \N__79269\,
            I => \N__79171\
        );

    \I__20069\ : Span4Mux_h
    port map (
            O => \N__79262\,
            I => \N__79171\
        );

    \I__20068\ : LocalMux
    port map (
            O => \N__79259\,
            I => \N__79162\
        );

    \I__20067\ : LocalMux
    port map (
            O => \N__79256\,
            I => \N__79162\
        );

    \I__20066\ : Span4Mux_h
    port map (
            O => \N__79253\,
            I => \N__79162\
        );

    \I__20065\ : LocalMux
    port map (
            O => \N__79250\,
            I => \N__79162\
        );

    \I__20064\ : InMux
    port map (
            O => \N__79249\,
            I => \N__79157\
        );

    \I__20063\ : InMux
    port map (
            O => \N__79248\,
            I => \N__79157\
        );

    \I__20062\ : Span4Mux_v
    port map (
            O => \N__79245\,
            I => \N__79150\
        );

    \I__20061\ : LocalMux
    port map (
            O => \N__79238\,
            I => \N__79150\
        );

    \I__20060\ : LocalMux
    port map (
            O => \N__79233\,
            I => \N__79150\
        );

    \I__20059\ : LocalMux
    port map (
            O => \N__79228\,
            I => \N__79143\
        );

    \I__20058\ : LocalMux
    port map (
            O => \N__79223\,
            I => \N__79143\
        );

    \I__20057\ : LocalMux
    port map (
            O => \N__79220\,
            I => \N__79143\
        );

    \I__20056\ : Span4Mux_v
    port map (
            O => \N__79217\,
            I => \N__79139\
        );

    \I__20055\ : Span4Mux_h
    port map (
            O => \N__79214\,
            I => \N__79134\
        );

    \I__20054\ : Span4Mux_h
    port map (
            O => \N__79211\,
            I => \N__79134\
        );

    \I__20053\ : InMux
    port map (
            O => \N__79210\,
            I => \N__79131\
        );

    \I__20052\ : InMux
    port map (
            O => \N__79209\,
            I => \N__79126\
        );

    \I__20051\ : InMux
    port map (
            O => \N__79208\,
            I => \N__79126\
        );

    \I__20050\ : InMux
    port map (
            O => \N__79207\,
            I => \N__79123\
        );

    \I__20049\ : LocalMux
    port map (
            O => \N__79204\,
            I => \N__79116\
        );

    \I__20048\ : LocalMux
    port map (
            O => \N__79201\,
            I => \N__79116\
        );

    \I__20047\ : LocalMux
    port map (
            O => \N__79196\,
            I => \N__79116\
        );

    \I__20046\ : Span4Mux_h
    port map (
            O => \N__79193\,
            I => \N__79111\
        );

    \I__20045\ : LocalMux
    port map (
            O => \N__79190\,
            I => \N__79111\
        );

    \I__20044\ : Span4Mux_v
    port map (
            O => \N__79185\,
            I => \N__79104\
        );

    \I__20043\ : LocalMux
    port map (
            O => \N__79182\,
            I => \N__79104\
        );

    \I__20042\ : Span4Mux_h
    port map (
            O => \N__79179\,
            I => \N__79104\
        );

    \I__20041\ : Span4Mux_h
    port map (
            O => \N__79176\,
            I => \N__79091\
        );

    \I__20040\ : Span4Mux_v
    port map (
            O => \N__79171\,
            I => \N__79091\
        );

    \I__20039\ : Span4Mux_v
    port map (
            O => \N__79162\,
            I => \N__79091\
        );

    \I__20038\ : LocalMux
    port map (
            O => \N__79157\,
            I => \N__79091\
        );

    \I__20037\ : Span4Mux_h
    port map (
            O => \N__79150\,
            I => \N__79091\
        );

    \I__20036\ : Span4Mux_v
    port map (
            O => \N__79143\,
            I => \N__79091\
        );

    \I__20035\ : InMux
    port map (
            O => \N__79142\,
            I => \N__79088\
        );

    \I__20034\ : Odrv4
    port map (
            O => \N__79139\,
            I => \progRomAddress_6\
        );

    \I__20033\ : Odrv4
    port map (
            O => \N__79134\,
            I => \progRomAddress_6\
        );

    \I__20032\ : LocalMux
    port map (
            O => \N__79131\,
            I => \progRomAddress_6\
        );

    \I__20031\ : LocalMux
    port map (
            O => \N__79126\,
            I => \progRomAddress_6\
        );

    \I__20030\ : LocalMux
    port map (
            O => \N__79123\,
            I => \progRomAddress_6\
        );

    \I__20029\ : Odrv4
    port map (
            O => \N__79116\,
            I => \progRomAddress_6\
        );

    \I__20028\ : Odrv4
    port map (
            O => \N__79111\,
            I => \progRomAddress_6\
        );

    \I__20027\ : Odrv4
    port map (
            O => \N__79104\,
            I => \progRomAddress_6\
        );

    \I__20026\ : Odrv4
    port map (
            O => \N__79091\,
            I => \progRomAddress_6\
        );

    \I__20025\ : LocalMux
    port map (
            O => \N__79088\,
            I => \progRomAddress_6\
        );

    \I__20024\ : CascadeMux
    port map (
            O => \N__79067\,
            I => \PROM.ROMDATA.m343_ns_1_cascade_\
        );

    \I__20023\ : CascadeMux
    port map (
            O => \N__79064\,
            I => \N__79061\
        );

    \I__20022\ : InMux
    port map (
            O => \N__79061\,
            I => \N__79058\
        );

    \I__20021\ : LocalMux
    port map (
            O => \N__79058\,
            I => \N__79055\
        );

    \I__20020\ : Span4Mux_h
    port map (
            O => \N__79055\,
            I => \N__79052\
        );

    \I__20019\ : Odrv4
    port map (
            O => \N__79052\,
            I => \PROM.ROMDATA.m343_ns\
        );

    \I__20018\ : CascadeMux
    port map (
            O => \N__79049\,
            I => \N__79045\
        );

    \I__20017\ : CascadeMux
    port map (
            O => \N__79048\,
            I => \N__79040\
        );

    \I__20016\ : InMux
    port map (
            O => \N__79045\,
            I => \N__79037\
        );

    \I__20015\ : InMux
    port map (
            O => \N__79044\,
            I => \N__79034\
        );

    \I__20014\ : CascadeMux
    port map (
            O => \N__79043\,
            I => \N__79030\
        );

    \I__20013\ : InMux
    port map (
            O => \N__79040\,
            I => \N__79027\
        );

    \I__20012\ : LocalMux
    port map (
            O => \N__79037\,
            I => \N__79024\
        );

    \I__20011\ : LocalMux
    port map (
            O => \N__79034\,
            I => \N__79021\
        );

    \I__20010\ : InMux
    port map (
            O => \N__79033\,
            I => \N__79016\
        );

    \I__20009\ : InMux
    port map (
            O => \N__79030\,
            I => \N__79016\
        );

    \I__20008\ : LocalMux
    port map (
            O => \N__79027\,
            I => \N__79011\
        );

    \I__20007\ : Span4Mux_h
    port map (
            O => \N__79024\,
            I => \N__79011\
        );

    \I__20006\ : Span4Mux_v
    port map (
            O => \N__79021\,
            I => \N__79006\
        );

    \I__20005\ : LocalMux
    port map (
            O => \N__79016\,
            I => \N__79006\
        );

    \I__20004\ : Span4Mux_v
    port map (
            O => \N__79011\,
            I => \N__79001\
        );

    \I__20003\ : Span4Mux_h
    port map (
            O => \N__79006\,
            I => \N__79001\
        );

    \I__20002\ : Odrv4
    port map (
            O => \N__79001\,
            I => \PROM.ROMDATA.m4\
        );

    \I__20001\ : InMux
    port map (
            O => \N__78998\,
            I => \N__78990\
        );

    \I__20000\ : InMux
    port map (
            O => \N__78997\,
            I => \N__78985\
        );

    \I__19999\ : InMux
    port map (
            O => \N__78996\,
            I => \N__78981\
        );

    \I__19998\ : InMux
    port map (
            O => \N__78995\,
            I => \N__78977\
        );

    \I__19997\ : InMux
    port map (
            O => \N__78994\,
            I => \N__78972\
        );

    \I__19996\ : InMux
    port map (
            O => \N__78993\,
            I => \N__78972\
        );

    \I__19995\ : LocalMux
    port map (
            O => \N__78990\,
            I => \N__78969\
        );

    \I__19994\ : InMux
    port map (
            O => \N__78989\,
            I => \N__78966\
        );

    \I__19993\ : InMux
    port map (
            O => \N__78988\,
            I => \N__78963\
        );

    \I__19992\ : LocalMux
    port map (
            O => \N__78985\,
            I => \N__78960\
        );

    \I__19991\ : InMux
    port map (
            O => \N__78984\,
            I => \N__78957\
        );

    \I__19990\ : LocalMux
    port map (
            O => \N__78981\,
            I => \N__78952\
        );

    \I__19989\ : InMux
    port map (
            O => \N__78980\,
            I => \N__78949\
        );

    \I__19988\ : LocalMux
    port map (
            O => \N__78977\,
            I => \N__78944\
        );

    \I__19987\ : LocalMux
    port map (
            O => \N__78972\,
            I => \N__78944\
        );

    \I__19986\ : Span4Mux_v
    port map (
            O => \N__78969\,
            I => \N__78940\
        );

    \I__19985\ : LocalMux
    port map (
            O => \N__78966\,
            I => \N__78937\
        );

    \I__19984\ : LocalMux
    port map (
            O => \N__78963\,
            I => \N__78934\
        );

    \I__19983\ : Span4Mux_v
    port map (
            O => \N__78960\,
            I => \N__78929\
        );

    \I__19982\ : LocalMux
    port map (
            O => \N__78957\,
            I => \N__78929\
        );

    \I__19981\ : InMux
    port map (
            O => \N__78956\,
            I => \N__78924\
        );

    \I__19980\ : InMux
    port map (
            O => \N__78955\,
            I => \N__78924\
        );

    \I__19979\ : Span4Mux_h
    port map (
            O => \N__78952\,
            I => \N__78921\
        );

    \I__19978\ : LocalMux
    port map (
            O => \N__78949\,
            I => \N__78918\
        );

    \I__19977\ : Span4Mux_v
    port map (
            O => \N__78944\,
            I => \N__78915\
        );

    \I__19976\ : InMux
    port map (
            O => \N__78943\,
            I => \N__78912\
        );

    \I__19975\ : Span4Mux_h
    port map (
            O => \N__78940\,
            I => \N__78905\
        );

    \I__19974\ : Span4Mux_v
    port map (
            O => \N__78937\,
            I => \N__78905\
        );

    \I__19973\ : Span4Mux_v
    port map (
            O => \N__78934\,
            I => \N__78905\
        );

    \I__19972\ : Span4Mux_h
    port map (
            O => \N__78929\,
            I => \N__78900\
        );

    \I__19971\ : LocalMux
    port map (
            O => \N__78924\,
            I => \N__78900\
        );

    \I__19970\ : Odrv4
    port map (
            O => \N__78921\,
            I => \PROM.ROMDATA.N_28_i\
        );

    \I__19969\ : Odrv4
    port map (
            O => \N__78918\,
            I => \PROM.ROMDATA.N_28_i\
        );

    \I__19968\ : Odrv4
    port map (
            O => \N__78915\,
            I => \PROM.ROMDATA.N_28_i\
        );

    \I__19967\ : LocalMux
    port map (
            O => \N__78912\,
            I => \PROM.ROMDATA.N_28_i\
        );

    \I__19966\ : Odrv4
    port map (
            O => \N__78905\,
            I => \PROM.ROMDATA.N_28_i\
        );

    \I__19965\ : Odrv4
    port map (
            O => \N__78900\,
            I => \PROM.ROMDATA.N_28_i\
        );

    \I__19964\ : InMux
    port map (
            O => \N__78887\,
            I => \N__78884\
        );

    \I__19963\ : LocalMux
    port map (
            O => \N__78884\,
            I => \N__78881\
        );

    \I__19962\ : Span12Mux_s10_h
    port map (
            O => \N__78881\,
            I => \N__78878\
        );

    \I__19961\ : Odrv12
    port map (
            O => \N__78878\,
            I => \PROM.ROMDATA.m183\
        );

    \I__19960\ : CascadeMux
    port map (
            O => \N__78875\,
            I => \PROM.ROMDATA.m334_ns_1_cascade_\
        );

    \I__19959\ : CascadeMux
    port map (
            O => \N__78872\,
            I => \N__78869\
        );

    \I__19958\ : InMux
    port map (
            O => \N__78869\,
            I => \N__78866\
        );

    \I__19957\ : LocalMux
    port map (
            O => \N__78866\,
            I => \PROM.ROMDATA.i3_mux_0\
        );

    \I__19956\ : CascadeMux
    port map (
            O => \N__78863\,
            I => \N__78846\
        );

    \I__19955\ : CascadeMux
    port map (
            O => \N__78862\,
            I => \N__78824\
        );

    \I__19954\ : CascadeMux
    port map (
            O => \N__78861\,
            I => \N__78820\
        );

    \I__19953\ : CascadeMux
    port map (
            O => \N__78860\,
            I => \N__78815\
        );

    \I__19952\ : InMux
    port map (
            O => \N__78859\,
            I => \N__78799\
        );

    \I__19951\ : InMux
    port map (
            O => \N__78858\,
            I => \N__78799\
        );

    \I__19950\ : InMux
    port map (
            O => \N__78857\,
            I => \N__78799\
        );

    \I__19949\ : InMux
    port map (
            O => \N__78856\,
            I => \N__78780\
        );

    \I__19948\ : InMux
    port map (
            O => \N__78855\,
            I => \N__78780\
        );

    \I__19947\ : InMux
    port map (
            O => \N__78854\,
            I => \N__78780\
        );

    \I__19946\ : InMux
    port map (
            O => \N__78853\,
            I => \N__78770\
        );

    \I__19945\ : InMux
    port map (
            O => \N__78852\,
            I => \N__78761\
        );

    \I__19944\ : InMux
    port map (
            O => \N__78851\,
            I => \N__78761\
        );

    \I__19943\ : InMux
    port map (
            O => \N__78850\,
            I => \N__78754\
        );

    \I__19942\ : InMux
    port map (
            O => \N__78849\,
            I => \N__78754\
        );

    \I__19941\ : InMux
    port map (
            O => \N__78846\,
            I => \N__78754\
        );

    \I__19940\ : CascadeMux
    port map (
            O => \N__78845\,
            I => \N__78750\
        );

    \I__19939\ : CascadeMux
    port map (
            O => \N__78844\,
            I => \N__78747\
        );

    \I__19938\ : InMux
    port map (
            O => \N__78843\,
            I => \N__78741\
        );

    \I__19937\ : InMux
    port map (
            O => \N__78842\,
            I => \N__78738\
        );

    \I__19936\ : InMux
    port map (
            O => \N__78841\,
            I => \N__78724\
        );

    \I__19935\ : InMux
    port map (
            O => \N__78840\,
            I => \N__78721\
        );

    \I__19934\ : CascadeMux
    port map (
            O => \N__78839\,
            I => \N__78715\
        );

    \I__19933\ : InMux
    port map (
            O => \N__78838\,
            I => \N__78705\
        );

    \I__19932\ : InMux
    port map (
            O => \N__78837\,
            I => \N__78705\
        );

    \I__19931\ : InMux
    port map (
            O => \N__78836\,
            I => \N__78705\
        );

    \I__19930\ : CascadeMux
    port map (
            O => \N__78835\,
            I => \N__78701\
        );

    \I__19929\ : CascadeMux
    port map (
            O => \N__78834\,
            I => \N__78697\
        );

    \I__19928\ : CascadeMux
    port map (
            O => \N__78833\,
            I => \N__78689\
        );

    \I__19927\ : InMux
    port map (
            O => \N__78832\,
            I => \N__78680\
        );

    \I__19926\ : InMux
    port map (
            O => \N__78831\,
            I => \N__78680\
        );

    \I__19925\ : InMux
    port map (
            O => \N__78830\,
            I => \N__78672\
        );

    \I__19924\ : InMux
    port map (
            O => \N__78829\,
            I => \N__78672\
        );

    \I__19923\ : InMux
    port map (
            O => \N__78828\,
            I => \N__78663\
        );

    \I__19922\ : InMux
    port map (
            O => \N__78827\,
            I => \N__78663\
        );

    \I__19921\ : InMux
    port map (
            O => \N__78824\,
            I => \N__78663\
        );

    \I__19920\ : InMux
    port map (
            O => \N__78823\,
            I => \N__78663\
        );

    \I__19919\ : InMux
    port map (
            O => \N__78820\,
            I => \N__78652\
        );

    \I__19918\ : InMux
    port map (
            O => \N__78819\,
            I => \N__78652\
        );

    \I__19917\ : InMux
    port map (
            O => \N__78818\,
            I => \N__78652\
        );

    \I__19916\ : InMux
    port map (
            O => \N__78815\,
            I => \N__78652\
        );

    \I__19915\ : InMux
    port map (
            O => \N__78814\,
            I => \N__78652\
        );

    \I__19914\ : InMux
    port map (
            O => \N__78813\,
            I => \N__78641\
        );

    \I__19913\ : InMux
    port map (
            O => \N__78812\,
            I => \N__78641\
        );

    \I__19912\ : InMux
    port map (
            O => \N__78811\,
            I => \N__78641\
        );

    \I__19911\ : InMux
    port map (
            O => \N__78810\,
            I => \N__78641\
        );

    \I__19910\ : InMux
    port map (
            O => \N__78809\,
            I => \N__78641\
        );

    \I__19909\ : InMux
    port map (
            O => \N__78808\,
            I => \N__78631\
        );

    \I__19908\ : InMux
    port map (
            O => \N__78807\,
            I => \N__78626\
        );

    \I__19907\ : InMux
    port map (
            O => \N__78806\,
            I => \N__78626\
        );

    \I__19906\ : LocalMux
    port map (
            O => \N__78799\,
            I => \N__78622\
        );

    \I__19905\ : InMux
    port map (
            O => \N__78798\,
            I => \N__78613\
        );

    \I__19904\ : InMux
    port map (
            O => \N__78797\,
            I => \N__78613\
        );

    \I__19903\ : InMux
    port map (
            O => \N__78796\,
            I => \N__78613\
        );

    \I__19902\ : InMux
    port map (
            O => \N__78795\,
            I => \N__78613\
        );

    \I__19901\ : InMux
    port map (
            O => \N__78794\,
            I => \N__78606\
        );

    \I__19900\ : InMux
    port map (
            O => \N__78793\,
            I => \N__78606\
        );

    \I__19899\ : InMux
    port map (
            O => \N__78792\,
            I => \N__78606\
        );

    \I__19898\ : InMux
    port map (
            O => \N__78791\,
            I => \N__78597\
        );

    \I__19897\ : InMux
    port map (
            O => \N__78790\,
            I => \N__78597\
        );

    \I__19896\ : InMux
    port map (
            O => \N__78789\,
            I => \N__78597\
        );

    \I__19895\ : InMux
    port map (
            O => \N__78788\,
            I => \N__78597\
        );

    \I__19894\ : InMux
    port map (
            O => \N__78787\,
            I => \N__78594\
        );

    \I__19893\ : LocalMux
    port map (
            O => \N__78780\,
            I => \N__78591\
        );

    \I__19892\ : InMux
    port map (
            O => \N__78779\,
            I => \N__78588\
        );

    \I__19891\ : InMux
    port map (
            O => \N__78778\,
            I => \N__78583\
        );

    \I__19890\ : InMux
    port map (
            O => \N__78777\,
            I => \N__78583\
        );

    \I__19889\ : InMux
    port map (
            O => \N__78776\,
            I => \N__78574\
        );

    \I__19888\ : InMux
    port map (
            O => \N__78775\,
            I => \N__78574\
        );

    \I__19887\ : InMux
    port map (
            O => \N__78774\,
            I => \N__78574\
        );

    \I__19886\ : InMux
    port map (
            O => \N__78773\,
            I => \N__78574\
        );

    \I__19885\ : LocalMux
    port map (
            O => \N__78770\,
            I => \N__78570\
        );

    \I__19884\ : InMux
    port map (
            O => \N__78769\,
            I => \N__78560\
        );

    \I__19883\ : InMux
    port map (
            O => \N__78768\,
            I => \N__78560\
        );

    \I__19882\ : InMux
    port map (
            O => \N__78767\,
            I => \N__78560\
        );

    \I__19881\ : InMux
    port map (
            O => \N__78766\,
            I => \N__78560\
        );

    \I__19880\ : LocalMux
    port map (
            O => \N__78761\,
            I => \N__78555\
        );

    \I__19879\ : LocalMux
    port map (
            O => \N__78754\,
            I => \N__78555\
        );

    \I__19878\ : InMux
    port map (
            O => \N__78753\,
            I => \N__78552\
        );

    \I__19877\ : InMux
    port map (
            O => \N__78750\,
            I => \N__78547\
        );

    \I__19876\ : InMux
    port map (
            O => \N__78747\,
            I => \N__78547\
        );

    \I__19875\ : InMux
    port map (
            O => \N__78746\,
            I => \N__78544\
        );

    \I__19874\ : InMux
    port map (
            O => \N__78745\,
            I => \N__78537\
        );

    \I__19873\ : InMux
    port map (
            O => \N__78744\,
            I => \N__78537\
        );

    \I__19872\ : LocalMux
    port map (
            O => \N__78741\,
            I => \N__78532\
        );

    \I__19871\ : LocalMux
    port map (
            O => \N__78738\,
            I => \N__78532\
        );

    \I__19870\ : InMux
    port map (
            O => \N__78737\,
            I => \N__78523\
        );

    \I__19869\ : InMux
    port map (
            O => \N__78736\,
            I => \N__78523\
        );

    \I__19868\ : InMux
    port map (
            O => \N__78735\,
            I => \N__78523\
        );

    \I__19867\ : InMux
    port map (
            O => \N__78734\,
            I => \N__78523\
        );

    \I__19866\ : InMux
    port map (
            O => \N__78733\,
            I => \N__78516\
        );

    \I__19865\ : InMux
    port map (
            O => \N__78732\,
            I => \N__78516\
        );

    \I__19864\ : InMux
    port map (
            O => \N__78731\,
            I => \N__78516\
        );

    \I__19863\ : InMux
    port map (
            O => \N__78730\,
            I => \N__78507\
        );

    \I__19862\ : InMux
    port map (
            O => \N__78729\,
            I => \N__78507\
        );

    \I__19861\ : InMux
    port map (
            O => \N__78728\,
            I => \N__78507\
        );

    \I__19860\ : InMux
    port map (
            O => \N__78727\,
            I => \N__78507\
        );

    \I__19859\ : LocalMux
    port map (
            O => \N__78724\,
            I => \N__78502\
        );

    \I__19858\ : LocalMux
    port map (
            O => \N__78721\,
            I => \N__78499\
        );

    \I__19857\ : InMux
    port map (
            O => \N__78720\,
            I => \N__78496\
        );

    \I__19856\ : InMux
    port map (
            O => \N__78719\,
            I => \N__78489\
        );

    \I__19855\ : InMux
    port map (
            O => \N__78718\,
            I => \N__78489\
        );

    \I__19854\ : InMux
    port map (
            O => \N__78715\,
            I => \N__78489\
        );

    \I__19853\ : InMux
    port map (
            O => \N__78714\,
            I => \N__78484\
        );

    \I__19852\ : InMux
    port map (
            O => \N__78713\,
            I => \N__78484\
        );

    \I__19851\ : InMux
    port map (
            O => \N__78712\,
            I => \N__78479\
        );

    \I__19850\ : LocalMux
    port map (
            O => \N__78705\,
            I => \N__78476\
        );

    \I__19849\ : CascadeMux
    port map (
            O => \N__78704\,
            I => \N__78469\
        );

    \I__19848\ : InMux
    port map (
            O => \N__78701\,
            I => \N__78457\
        );

    \I__19847\ : InMux
    port map (
            O => \N__78700\,
            I => \N__78457\
        );

    \I__19846\ : InMux
    port map (
            O => \N__78697\,
            I => \N__78457\
        );

    \I__19845\ : InMux
    port map (
            O => \N__78696\,
            I => \N__78457\
        );

    \I__19844\ : InMux
    port map (
            O => \N__78695\,
            I => \N__78457\
        );

    \I__19843\ : InMux
    port map (
            O => \N__78694\,
            I => \N__78454\
        );

    \I__19842\ : InMux
    port map (
            O => \N__78693\,
            I => \N__78447\
        );

    \I__19841\ : InMux
    port map (
            O => \N__78692\,
            I => \N__78447\
        );

    \I__19840\ : InMux
    port map (
            O => \N__78689\,
            I => \N__78447\
        );

    \I__19839\ : InMux
    port map (
            O => \N__78688\,
            I => \N__78442\
        );

    \I__19838\ : InMux
    port map (
            O => \N__78687\,
            I => \N__78442\
        );

    \I__19837\ : InMux
    port map (
            O => \N__78686\,
            I => \N__78437\
        );

    \I__19836\ : InMux
    port map (
            O => \N__78685\,
            I => \N__78437\
        );

    \I__19835\ : LocalMux
    port map (
            O => \N__78680\,
            I => \N__78434\
        );

    \I__19834\ : InMux
    port map (
            O => \N__78679\,
            I => \N__78431\
        );

    \I__19833\ : InMux
    port map (
            O => \N__78678\,
            I => \N__78426\
        );

    \I__19832\ : InMux
    port map (
            O => \N__78677\,
            I => \N__78426\
        );

    \I__19831\ : LocalMux
    port map (
            O => \N__78672\,
            I => \N__78417\
        );

    \I__19830\ : LocalMux
    port map (
            O => \N__78663\,
            I => \N__78417\
        );

    \I__19829\ : LocalMux
    port map (
            O => \N__78652\,
            I => \N__78417\
        );

    \I__19828\ : LocalMux
    port map (
            O => \N__78641\,
            I => \N__78417\
        );

    \I__19827\ : InMux
    port map (
            O => \N__78640\,
            I => \N__78410\
        );

    \I__19826\ : InMux
    port map (
            O => \N__78639\,
            I => \N__78410\
        );

    \I__19825\ : InMux
    port map (
            O => \N__78638\,
            I => \N__78410\
        );

    \I__19824\ : InMux
    port map (
            O => \N__78637\,
            I => \N__78407\
        );

    \I__19823\ : InMux
    port map (
            O => \N__78636\,
            I => \N__78399\
        );

    \I__19822\ : InMux
    port map (
            O => \N__78635\,
            I => \N__78399\
        );

    \I__19821\ : InMux
    port map (
            O => \N__78634\,
            I => \N__78396\
        );

    \I__19820\ : LocalMux
    port map (
            O => \N__78631\,
            I => \N__78391\
        );

    \I__19819\ : LocalMux
    port map (
            O => \N__78626\,
            I => \N__78391\
        );

    \I__19818\ : InMux
    port map (
            O => \N__78625\,
            I => \N__78388\
        );

    \I__19817\ : Span4Mux_h
    port map (
            O => \N__78622\,
            I => \N__78379\
        );

    \I__19816\ : LocalMux
    port map (
            O => \N__78613\,
            I => \N__78379\
        );

    \I__19815\ : LocalMux
    port map (
            O => \N__78606\,
            I => \N__78379\
        );

    \I__19814\ : LocalMux
    port map (
            O => \N__78597\,
            I => \N__78379\
        );

    \I__19813\ : LocalMux
    port map (
            O => \N__78594\,
            I => \N__78372\
        );

    \I__19812\ : Span4Mux_v
    port map (
            O => \N__78591\,
            I => \N__78372\
        );

    \I__19811\ : LocalMux
    port map (
            O => \N__78588\,
            I => \N__78372\
        );

    \I__19810\ : LocalMux
    port map (
            O => \N__78583\,
            I => \N__78369\
        );

    \I__19809\ : LocalMux
    port map (
            O => \N__78574\,
            I => \N__78366\
        );

    \I__19808\ : CascadeMux
    port map (
            O => \N__78573\,
            I => \N__78363\
        );

    \I__19807\ : Span4Mux_v
    port map (
            O => \N__78570\,
            I => \N__78355\
        );

    \I__19806\ : InMux
    port map (
            O => \N__78569\,
            I => \N__78352\
        );

    \I__19805\ : LocalMux
    port map (
            O => \N__78560\,
            I => \N__78345\
        );

    \I__19804\ : Span4Mux_h
    port map (
            O => \N__78555\,
            I => \N__78345\
        );

    \I__19803\ : LocalMux
    port map (
            O => \N__78552\,
            I => \N__78345\
        );

    \I__19802\ : LocalMux
    port map (
            O => \N__78547\,
            I => \N__78340\
        );

    \I__19801\ : LocalMux
    port map (
            O => \N__78544\,
            I => \N__78340\
        );

    \I__19800\ : CascadeMux
    port map (
            O => \N__78543\,
            I => \N__78316\
        );

    \I__19799\ : InMux
    port map (
            O => \N__78542\,
            I => \N__78312\
        );

    \I__19798\ : LocalMux
    port map (
            O => \N__78537\,
            I => \N__78305\
        );

    \I__19797\ : Span4Mux_h
    port map (
            O => \N__78532\,
            I => \N__78305\
        );

    \I__19796\ : LocalMux
    port map (
            O => \N__78523\,
            I => \N__78305\
        );

    \I__19795\ : LocalMux
    port map (
            O => \N__78516\,
            I => \N__78300\
        );

    \I__19794\ : LocalMux
    port map (
            O => \N__78507\,
            I => \N__78300\
        );

    \I__19793\ : InMux
    port map (
            O => \N__78506\,
            I => \N__78295\
        );

    \I__19792\ : InMux
    port map (
            O => \N__78505\,
            I => \N__78295\
        );

    \I__19791\ : Span4Mux_h
    port map (
            O => \N__78502\,
            I => \N__78290\
        );

    \I__19790\ : Span4Mux_h
    port map (
            O => \N__78499\,
            I => \N__78290\
        );

    \I__19789\ : LocalMux
    port map (
            O => \N__78496\,
            I => \N__78287\
        );

    \I__19788\ : LocalMux
    port map (
            O => \N__78489\,
            I => \N__78282\
        );

    \I__19787\ : LocalMux
    port map (
            O => \N__78484\,
            I => \N__78282\
        );

    \I__19786\ : InMux
    port map (
            O => \N__78483\,
            I => \N__78277\
        );

    \I__19785\ : InMux
    port map (
            O => \N__78482\,
            I => \N__78277\
        );

    \I__19784\ : LocalMux
    port map (
            O => \N__78479\,
            I => \N__78272\
        );

    \I__19783\ : Span4Mux_v
    port map (
            O => \N__78476\,
            I => \N__78272\
        );

    \I__19782\ : InMux
    port map (
            O => \N__78475\,
            I => \N__78265\
        );

    \I__19781\ : InMux
    port map (
            O => \N__78474\,
            I => \N__78265\
        );

    \I__19780\ : InMux
    port map (
            O => \N__78473\,
            I => \N__78265\
        );

    \I__19779\ : InMux
    port map (
            O => \N__78472\,
            I => \N__78258\
        );

    \I__19778\ : InMux
    port map (
            O => \N__78469\,
            I => \N__78258\
        );

    \I__19777\ : InMux
    port map (
            O => \N__78468\,
            I => \N__78258\
        );

    \I__19776\ : LocalMux
    port map (
            O => \N__78457\,
            I => \N__78237\
        );

    \I__19775\ : LocalMux
    port map (
            O => \N__78454\,
            I => \N__78237\
        );

    \I__19774\ : LocalMux
    port map (
            O => \N__78447\,
            I => \N__78237\
        );

    \I__19773\ : LocalMux
    port map (
            O => \N__78442\,
            I => \N__78237\
        );

    \I__19772\ : LocalMux
    port map (
            O => \N__78437\,
            I => \N__78237\
        );

    \I__19771\ : Span4Mux_h
    port map (
            O => \N__78434\,
            I => \N__78237\
        );

    \I__19770\ : LocalMux
    port map (
            O => \N__78431\,
            I => \N__78237\
        );

    \I__19769\ : LocalMux
    port map (
            O => \N__78426\,
            I => \N__78237\
        );

    \I__19768\ : Span4Mux_v
    port map (
            O => \N__78417\,
            I => \N__78237\
        );

    \I__19767\ : LocalMux
    port map (
            O => \N__78410\,
            I => \N__78237\
        );

    \I__19766\ : LocalMux
    port map (
            O => \N__78407\,
            I => \N__78234\
        );

    \I__19765\ : InMux
    port map (
            O => \N__78406\,
            I => \N__78227\
        );

    \I__19764\ : InMux
    port map (
            O => \N__78405\,
            I => \N__78227\
        );

    \I__19763\ : InMux
    port map (
            O => \N__78404\,
            I => \N__78227\
        );

    \I__19762\ : LocalMux
    port map (
            O => \N__78399\,
            I => \N__78214\
        );

    \I__19761\ : LocalMux
    port map (
            O => \N__78396\,
            I => \N__78214\
        );

    \I__19760\ : Span4Mux_v
    port map (
            O => \N__78391\,
            I => \N__78214\
        );

    \I__19759\ : LocalMux
    port map (
            O => \N__78388\,
            I => \N__78214\
        );

    \I__19758\ : Span4Mux_v
    port map (
            O => \N__78379\,
            I => \N__78214\
        );

    \I__19757\ : Span4Mux_h
    port map (
            O => \N__78372\,
            I => \N__78214\
        );

    \I__19756\ : Span4Mux_h
    port map (
            O => \N__78369\,
            I => \N__78209\
        );

    \I__19755\ : Span4Mux_v
    port map (
            O => \N__78366\,
            I => \N__78209\
        );

    \I__19754\ : InMux
    port map (
            O => \N__78363\,
            I => \N__78206\
        );

    \I__19753\ : InMux
    port map (
            O => \N__78362\,
            I => \N__78203\
        );

    \I__19752\ : InMux
    port map (
            O => \N__78361\,
            I => \N__78194\
        );

    \I__19751\ : InMux
    port map (
            O => \N__78360\,
            I => \N__78194\
        );

    \I__19750\ : InMux
    port map (
            O => \N__78359\,
            I => \N__78194\
        );

    \I__19749\ : InMux
    port map (
            O => \N__78358\,
            I => \N__78194\
        );

    \I__19748\ : Span4Mux_h
    port map (
            O => \N__78355\,
            I => \N__78185\
        );

    \I__19747\ : LocalMux
    port map (
            O => \N__78352\,
            I => \N__78185\
        );

    \I__19746\ : Span4Mux_v
    port map (
            O => \N__78345\,
            I => \N__78185\
        );

    \I__19745\ : Span4Mux_v
    port map (
            O => \N__78340\,
            I => \N__78185\
        );

    \I__19744\ : InMux
    port map (
            O => \N__78339\,
            I => \N__78178\
        );

    \I__19743\ : InMux
    port map (
            O => \N__78338\,
            I => \N__78178\
        );

    \I__19742\ : InMux
    port map (
            O => \N__78337\,
            I => \N__78178\
        );

    \I__19741\ : InMux
    port map (
            O => \N__78336\,
            I => \N__78169\
        );

    \I__19740\ : InMux
    port map (
            O => \N__78335\,
            I => \N__78169\
        );

    \I__19739\ : InMux
    port map (
            O => \N__78334\,
            I => \N__78169\
        );

    \I__19738\ : InMux
    port map (
            O => \N__78333\,
            I => \N__78169\
        );

    \I__19737\ : InMux
    port map (
            O => \N__78332\,
            I => \N__78160\
        );

    \I__19736\ : InMux
    port map (
            O => \N__78331\,
            I => \N__78160\
        );

    \I__19735\ : InMux
    port map (
            O => \N__78330\,
            I => \N__78160\
        );

    \I__19734\ : InMux
    port map (
            O => \N__78329\,
            I => \N__78160\
        );

    \I__19733\ : InMux
    port map (
            O => \N__78328\,
            I => \N__78151\
        );

    \I__19732\ : InMux
    port map (
            O => \N__78327\,
            I => \N__78151\
        );

    \I__19731\ : InMux
    port map (
            O => \N__78326\,
            I => \N__78151\
        );

    \I__19730\ : InMux
    port map (
            O => \N__78325\,
            I => \N__78151\
        );

    \I__19729\ : InMux
    port map (
            O => \N__78324\,
            I => \N__78142\
        );

    \I__19728\ : InMux
    port map (
            O => \N__78323\,
            I => \N__78142\
        );

    \I__19727\ : InMux
    port map (
            O => \N__78322\,
            I => \N__78142\
        );

    \I__19726\ : InMux
    port map (
            O => \N__78321\,
            I => \N__78142\
        );

    \I__19725\ : InMux
    port map (
            O => \N__78320\,
            I => \N__78133\
        );

    \I__19724\ : InMux
    port map (
            O => \N__78319\,
            I => \N__78133\
        );

    \I__19723\ : InMux
    port map (
            O => \N__78316\,
            I => \N__78133\
        );

    \I__19722\ : InMux
    port map (
            O => \N__78315\,
            I => \N__78133\
        );

    \I__19721\ : LocalMux
    port map (
            O => \N__78312\,
            I => \N__78124\
        );

    \I__19720\ : Span4Mux_v
    port map (
            O => \N__78305\,
            I => \N__78124\
        );

    \I__19719\ : Span4Mux_h
    port map (
            O => \N__78300\,
            I => \N__78124\
        );

    \I__19718\ : LocalMux
    port map (
            O => \N__78295\,
            I => \N__78124\
        );

    \I__19717\ : Span4Mux_v
    port map (
            O => \N__78290\,
            I => \N__78107\
        );

    \I__19716\ : Span4Mux_v
    port map (
            O => \N__78287\,
            I => \N__78107\
        );

    \I__19715\ : Span4Mux_v
    port map (
            O => \N__78282\,
            I => \N__78107\
        );

    \I__19714\ : LocalMux
    port map (
            O => \N__78277\,
            I => \N__78107\
        );

    \I__19713\ : Span4Mux_h
    port map (
            O => \N__78272\,
            I => \N__78107\
        );

    \I__19712\ : LocalMux
    port map (
            O => \N__78265\,
            I => \N__78107\
        );

    \I__19711\ : LocalMux
    port map (
            O => \N__78258\,
            I => \N__78107\
        );

    \I__19710\ : Span4Mux_v
    port map (
            O => \N__78237\,
            I => \N__78107\
        );

    \I__19709\ : Span4Mux_h
    port map (
            O => \N__78234\,
            I => \N__78100\
        );

    \I__19708\ : LocalMux
    port map (
            O => \N__78227\,
            I => \N__78100\
        );

    \I__19707\ : Span4Mux_h
    port map (
            O => \N__78214\,
            I => \N__78100\
        );

    \I__19706\ : Odrv4
    port map (
            O => \N__78209\,
            I => \progRomAddress_1\
        );

    \I__19705\ : LocalMux
    port map (
            O => \N__78206\,
            I => \progRomAddress_1\
        );

    \I__19704\ : LocalMux
    port map (
            O => \N__78203\,
            I => \progRomAddress_1\
        );

    \I__19703\ : LocalMux
    port map (
            O => \N__78194\,
            I => \progRomAddress_1\
        );

    \I__19702\ : Odrv4
    port map (
            O => \N__78185\,
            I => \progRomAddress_1\
        );

    \I__19701\ : LocalMux
    port map (
            O => \N__78178\,
            I => \progRomAddress_1\
        );

    \I__19700\ : LocalMux
    port map (
            O => \N__78169\,
            I => \progRomAddress_1\
        );

    \I__19699\ : LocalMux
    port map (
            O => \N__78160\,
            I => \progRomAddress_1\
        );

    \I__19698\ : LocalMux
    port map (
            O => \N__78151\,
            I => \progRomAddress_1\
        );

    \I__19697\ : LocalMux
    port map (
            O => \N__78142\,
            I => \progRomAddress_1\
        );

    \I__19696\ : LocalMux
    port map (
            O => \N__78133\,
            I => \progRomAddress_1\
        );

    \I__19695\ : Odrv4
    port map (
            O => \N__78124\,
            I => \progRomAddress_1\
        );

    \I__19694\ : Odrv4
    port map (
            O => \N__78107\,
            I => \progRomAddress_1\
        );

    \I__19693\ : Odrv4
    port map (
            O => \N__78100\,
            I => \progRomAddress_1\
        );

    \I__19692\ : CascadeMux
    port map (
            O => \N__78071\,
            I => \N__78056\
        );

    \I__19691\ : CascadeMux
    port map (
            O => \N__78070\,
            I => \N__78051\
        );

    \I__19690\ : InMux
    port map (
            O => \N__78069\,
            I => \N__78044\
        );

    \I__19689\ : InMux
    port map (
            O => \N__78068\,
            I => \N__78044\
        );

    \I__19688\ : InMux
    port map (
            O => \N__78067\,
            I => \N__78032\
        );

    \I__19687\ : InMux
    port map (
            O => \N__78066\,
            I => \N__78029\
        );

    \I__19686\ : InMux
    port map (
            O => \N__78065\,
            I => \N__78017\
        );

    \I__19685\ : InMux
    port map (
            O => \N__78064\,
            I => \N__78012\
        );

    \I__19684\ : InMux
    port map (
            O => \N__78063\,
            I => \N__78012\
        );

    \I__19683\ : InMux
    port map (
            O => \N__78062\,
            I => \N__78006\
        );

    \I__19682\ : InMux
    port map (
            O => \N__78061\,
            I => \N__78006\
        );

    \I__19681\ : InMux
    port map (
            O => \N__78060\,
            I => \N__78003\
        );

    \I__19680\ : InMux
    port map (
            O => \N__78059\,
            I => \N__77996\
        );

    \I__19679\ : InMux
    port map (
            O => \N__78056\,
            I => \N__77996\
        );

    \I__19678\ : InMux
    port map (
            O => \N__78055\,
            I => \N__77996\
        );

    \I__19677\ : CascadeMux
    port map (
            O => \N__78054\,
            I => \N__77990\
        );

    \I__19676\ : InMux
    port map (
            O => \N__78051\,
            I => \N__77983\
        );

    \I__19675\ : InMux
    port map (
            O => \N__78050\,
            I => \N__77983\
        );

    \I__19674\ : CascadeMux
    port map (
            O => \N__78049\,
            I => \N__77978\
        );

    \I__19673\ : LocalMux
    port map (
            O => \N__78044\,
            I => \N__77970\
        );

    \I__19672\ : CascadeMux
    port map (
            O => \N__78043\,
            I => \N__77967\
        );

    \I__19671\ : CascadeMux
    port map (
            O => \N__78042\,
            I => \N__77962\
        );

    \I__19670\ : InMux
    port map (
            O => \N__78041\,
            I => \N__77958\
        );

    \I__19669\ : CascadeMux
    port map (
            O => \N__78040\,
            I => \N__77950\
        );

    \I__19668\ : CascadeMux
    port map (
            O => \N__78039\,
            I => \N__77947\
        );

    \I__19667\ : CascadeMux
    port map (
            O => \N__78038\,
            I => \N__77944\
        );

    \I__19666\ : CascadeMux
    port map (
            O => \N__78037\,
            I => \N__77941\
        );

    \I__19665\ : CascadeMux
    port map (
            O => \N__78036\,
            I => \N__77937\
        );

    \I__19664\ : CascadeMux
    port map (
            O => \N__78035\,
            I => \N__77934\
        );

    \I__19663\ : LocalMux
    port map (
            O => \N__78032\,
            I => \N__77929\
        );

    \I__19662\ : LocalMux
    port map (
            O => \N__78029\,
            I => \N__77926\
        );

    \I__19661\ : InMux
    port map (
            O => \N__78028\,
            I => \N__77921\
        );

    \I__19660\ : InMux
    port map (
            O => \N__78027\,
            I => \N__77921\
        );

    \I__19659\ : InMux
    port map (
            O => \N__78026\,
            I => \N__77912\
        );

    \I__19658\ : InMux
    port map (
            O => \N__78025\,
            I => \N__77912\
        );

    \I__19657\ : InMux
    port map (
            O => \N__78024\,
            I => \N__77912\
        );

    \I__19656\ : InMux
    port map (
            O => \N__78023\,
            I => \N__77912\
        );

    \I__19655\ : CascadeMux
    port map (
            O => \N__78022\,
            I => \N__77903\
        );

    \I__19654\ : CascadeMux
    port map (
            O => \N__78021\,
            I => \N__77900\
        );

    \I__19653\ : CascadeMux
    port map (
            O => \N__78020\,
            I => \N__77889\
        );

    \I__19652\ : LocalMux
    port map (
            O => \N__78017\,
            I => \N__77870\
        );

    \I__19651\ : LocalMux
    port map (
            O => \N__78012\,
            I => \N__77867\
        );

    \I__19650\ : InMux
    port map (
            O => \N__78011\,
            I => \N__77859\
        );

    \I__19649\ : LocalMux
    port map (
            O => \N__78006\,
            I => \N__77856\
        );

    \I__19648\ : LocalMux
    port map (
            O => \N__78003\,
            I => \N__77853\
        );

    \I__19647\ : LocalMux
    port map (
            O => \N__77996\,
            I => \N__77850\
        );

    \I__19646\ : InMux
    port map (
            O => \N__77995\,
            I => \N__77847\
        );

    \I__19645\ : CascadeMux
    port map (
            O => \N__77994\,
            I => \N__77844\
        );

    \I__19644\ : InMux
    port map (
            O => \N__77993\,
            I => \N__77829\
        );

    \I__19643\ : InMux
    port map (
            O => \N__77990\,
            I => \N__77829\
        );

    \I__19642\ : InMux
    port map (
            O => \N__77989\,
            I => \N__77829\
        );

    \I__19641\ : InMux
    port map (
            O => \N__77988\,
            I => \N__77829\
        );

    \I__19640\ : LocalMux
    port map (
            O => \N__77983\,
            I => \N__77826\
        );

    \I__19639\ : InMux
    port map (
            O => \N__77982\,
            I => \N__77817\
        );

    \I__19638\ : InMux
    port map (
            O => \N__77981\,
            I => \N__77817\
        );

    \I__19637\ : InMux
    port map (
            O => \N__77978\,
            I => \N__77817\
        );

    \I__19636\ : InMux
    port map (
            O => \N__77977\,
            I => \N__77817\
        );

    \I__19635\ : CascadeMux
    port map (
            O => \N__77976\,
            I => \N__77813\
        );

    \I__19634\ : CascadeMux
    port map (
            O => \N__77975\,
            I => \N__77809\
        );

    \I__19633\ : CascadeMux
    port map (
            O => \N__77974\,
            I => \N__77800\
        );

    \I__19632\ : CascadeMux
    port map (
            O => \N__77973\,
            I => \N__77797\
        );

    \I__19631\ : Span4Mux_h
    port map (
            O => \N__77970\,
            I => \N__77790\
        );

    \I__19630\ : InMux
    port map (
            O => \N__77967\,
            I => \N__77785\
        );

    \I__19629\ : InMux
    port map (
            O => \N__77966\,
            I => \N__77785\
        );

    \I__19628\ : InMux
    port map (
            O => \N__77965\,
            I => \N__77778\
        );

    \I__19627\ : InMux
    port map (
            O => \N__77962\,
            I => \N__77778\
        );

    \I__19626\ : InMux
    port map (
            O => \N__77961\,
            I => \N__77778\
        );

    \I__19625\ : LocalMux
    port map (
            O => \N__77958\,
            I => \N__77775\
        );

    \I__19624\ : InMux
    port map (
            O => \N__77957\,
            I => \N__77766\
        );

    \I__19623\ : InMux
    port map (
            O => \N__77956\,
            I => \N__77766\
        );

    \I__19622\ : InMux
    port map (
            O => \N__77955\,
            I => \N__77766\
        );

    \I__19621\ : InMux
    port map (
            O => \N__77954\,
            I => \N__77766\
        );

    \I__19620\ : InMux
    port map (
            O => \N__77953\,
            I => \N__77755\
        );

    \I__19619\ : InMux
    port map (
            O => \N__77950\,
            I => \N__77755\
        );

    \I__19618\ : InMux
    port map (
            O => \N__77947\,
            I => \N__77755\
        );

    \I__19617\ : InMux
    port map (
            O => \N__77944\,
            I => \N__77755\
        );

    \I__19616\ : InMux
    port map (
            O => \N__77941\,
            I => \N__77755\
        );

    \I__19615\ : InMux
    port map (
            O => \N__77940\,
            I => \N__77752\
        );

    \I__19614\ : InMux
    port map (
            O => \N__77937\,
            I => \N__77745\
        );

    \I__19613\ : InMux
    port map (
            O => \N__77934\,
            I => \N__77745\
        );

    \I__19612\ : InMux
    port map (
            O => \N__77933\,
            I => \N__77745\
        );

    \I__19611\ : InMux
    port map (
            O => \N__77932\,
            I => \N__77740\
        );

    \I__19610\ : Span4Mux_h
    port map (
            O => \N__77929\,
            I => \N__77733\
        );

    \I__19609\ : Span4Mux_v
    port map (
            O => \N__77926\,
            I => \N__77733\
        );

    \I__19608\ : LocalMux
    port map (
            O => \N__77921\,
            I => \N__77733\
        );

    \I__19607\ : LocalMux
    port map (
            O => \N__77912\,
            I => \N__77730\
        );

    \I__19606\ : InMux
    port map (
            O => \N__77911\,
            I => \N__77723\
        );

    \I__19605\ : InMux
    port map (
            O => \N__77910\,
            I => \N__77723\
        );

    \I__19604\ : InMux
    port map (
            O => \N__77909\,
            I => \N__77723\
        );

    \I__19603\ : InMux
    port map (
            O => \N__77908\,
            I => \N__77720\
        );

    \I__19602\ : InMux
    port map (
            O => \N__77907\,
            I => \N__77715\
        );

    \I__19601\ : InMux
    port map (
            O => \N__77906\,
            I => \N__77715\
        );

    \I__19600\ : InMux
    port map (
            O => \N__77903\,
            I => \N__77708\
        );

    \I__19599\ : InMux
    port map (
            O => \N__77900\,
            I => \N__77708\
        );

    \I__19598\ : InMux
    port map (
            O => \N__77899\,
            I => \N__77708\
        );

    \I__19597\ : InMux
    port map (
            O => \N__77898\,
            I => \N__77701\
        );

    \I__19596\ : InMux
    port map (
            O => \N__77897\,
            I => \N__77701\
        );

    \I__19595\ : InMux
    port map (
            O => \N__77896\,
            I => \N__77701\
        );

    \I__19594\ : CascadeMux
    port map (
            O => \N__77895\,
            I => \N__77697\
        );

    \I__19593\ : CascadeMux
    port map (
            O => \N__77894\,
            I => \N__77694\
        );

    \I__19592\ : CascadeMux
    port map (
            O => \N__77893\,
            I => \N__77685\
        );

    \I__19591\ : InMux
    port map (
            O => \N__77892\,
            I => \N__77682\
        );

    \I__19590\ : InMux
    port map (
            O => \N__77889\,
            I => \N__77675\
        );

    \I__19589\ : InMux
    port map (
            O => \N__77888\,
            I => \N__77675\
        );

    \I__19588\ : InMux
    port map (
            O => \N__77887\,
            I => \N__77675\
        );

    \I__19587\ : InMux
    port map (
            O => \N__77886\,
            I => \N__77668\
        );

    \I__19586\ : InMux
    port map (
            O => \N__77885\,
            I => \N__77668\
        );

    \I__19585\ : InMux
    port map (
            O => \N__77884\,
            I => \N__77668\
        );

    \I__19584\ : InMux
    port map (
            O => \N__77883\,
            I => \N__77659\
        );

    \I__19583\ : InMux
    port map (
            O => \N__77882\,
            I => \N__77659\
        );

    \I__19582\ : InMux
    port map (
            O => \N__77881\,
            I => \N__77659\
        );

    \I__19581\ : InMux
    port map (
            O => \N__77880\,
            I => \N__77659\
        );

    \I__19580\ : InMux
    port map (
            O => \N__77879\,
            I => \N__77654\
        );

    \I__19579\ : InMux
    port map (
            O => \N__77878\,
            I => \N__77654\
        );

    \I__19578\ : InMux
    port map (
            O => \N__77877\,
            I => \N__77647\
        );

    \I__19577\ : InMux
    port map (
            O => \N__77876\,
            I => \N__77647\
        );

    \I__19576\ : InMux
    port map (
            O => \N__77875\,
            I => \N__77647\
        );

    \I__19575\ : InMux
    port map (
            O => \N__77874\,
            I => \N__77642\
        );

    \I__19574\ : InMux
    port map (
            O => \N__77873\,
            I => \N__77642\
        );

    \I__19573\ : Span4Mux_v
    port map (
            O => \N__77870\,
            I => \N__77639\
        );

    \I__19572\ : Span4Mux_v
    port map (
            O => \N__77867\,
            I => \N__77636\
        );

    \I__19571\ : InMux
    port map (
            O => \N__77866\,
            I => \N__77627\
        );

    \I__19570\ : InMux
    port map (
            O => \N__77865\,
            I => \N__77627\
        );

    \I__19569\ : InMux
    port map (
            O => \N__77864\,
            I => \N__77627\
        );

    \I__19568\ : InMux
    port map (
            O => \N__77863\,
            I => \N__77627\
        );

    \I__19567\ : InMux
    port map (
            O => \N__77862\,
            I => \N__77624\
        );

    \I__19566\ : LocalMux
    port map (
            O => \N__77859\,
            I => \N__77621\
        );

    \I__19565\ : Span4Mux_h
    port map (
            O => \N__77856\,
            I => \N__77605\
        );

    \I__19564\ : Span4Mux_h
    port map (
            O => \N__77853\,
            I => \N__77598\
        );

    \I__19563\ : Span4Mux_v
    port map (
            O => \N__77850\,
            I => \N__77598\
        );

    \I__19562\ : LocalMux
    port map (
            O => \N__77847\,
            I => \N__77598\
        );

    \I__19561\ : InMux
    port map (
            O => \N__77844\,
            I => \N__77591\
        );

    \I__19560\ : InMux
    port map (
            O => \N__77843\,
            I => \N__77591\
        );

    \I__19559\ : InMux
    port map (
            O => \N__77842\,
            I => \N__77591\
        );

    \I__19558\ : CascadeMux
    port map (
            O => \N__77841\,
            I => \N__77587\
        );

    \I__19557\ : CascadeMux
    port map (
            O => \N__77840\,
            I => \N__77584\
        );

    \I__19556\ : CascadeMux
    port map (
            O => \N__77839\,
            I => \N__77580\
        );

    \I__19555\ : CascadeMux
    port map (
            O => \N__77838\,
            I => \N__77577\
        );

    \I__19554\ : LocalMux
    port map (
            O => \N__77829\,
            I => \N__77568\
        );

    \I__19553\ : Span4Mux_h
    port map (
            O => \N__77826\,
            I => \N__77568\
        );

    \I__19552\ : LocalMux
    port map (
            O => \N__77817\,
            I => \N__77568\
        );

    \I__19551\ : InMux
    port map (
            O => \N__77816\,
            I => \N__77559\
        );

    \I__19550\ : InMux
    port map (
            O => \N__77813\,
            I => \N__77559\
        );

    \I__19549\ : InMux
    port map (
            O => \N__77812\,
            I => \N__77559\
        );

    \I__19548\ : InMux
    port map (
            O => \N__77809\,
            I => \N__77559\
        );

    \I__19547\ : InMux
    port map (
            O => \N__77808\,
            I => \N__77548\
        );

    \I__19546\ : InMux
    port map (
            O => \N__77807\,
            I => \N__77548\
        );

    \I__19545\ : InMux
    port map (
            O => \N__77806\,
            I => \N__77548\
        );

    \I__19544\ : InMux
    port map (
            O => \N__77805\,
            I => \N__77548\
        );

    \I__19543\ : InMux
    port map (
            O => \N__77804\,
            I => \N__77548\
        );

    \I__19542\ : InMux
    port map (
            O => \N__77803\,
            I => \N__77539\
        );

    \I__19541\ : InMux
    port map (
            O => \N__77800\,
            I => \N__77539\
        );

    \I__19540\ : InMux
    port map (
            O => \N__77797\,
            I => \N__77539\
        );

    \I__19539\ : InMux
    port map (
            O => \N__77796\,
            I => \N__77539\
        );

    \I__19538\ : InMux
    port map (
            O => \N__77795\,
            I => \N__77532\
        );

    \I__19537\ : InMux
    port map (
            O => \N__77794\,
            I => \N__77532\
        );

    \I__19536\ : InMux
    port map (
            O => \N__77793\,
            I => \N__77532\
        );

    \I__19535\ : Span4Mux_v
    port map (
            O => \N__77790\,
            I => \N__77525\
        );

    \I__19534\ : LocalMux
    port map (
            O => \N__77785\,
            I => \N__77525\
        );

    \I__19533\ : LocalMux
    port map (
            O => \N__77778\,
            I => \N__77525\
        );

    \I__19532\ : Span4Mux_h
    port map (
            O => \N__77775\,
            I => \N__77518\
        );

    \I__19531\ : LocalMux
    port map (
            O => \N__77766\,
            I => \N__77518\
        );

    \I__19530\ : LocalMux
    port map (
            O => \N__77755\,
            I => \N__77518\
        );

    \I__19529\ : LocalMux
    port map (
            O => \N__77752\,
            I => \N__77515\
        );

    \I__19528\ : LocalMux
    port map (
            O => \N__77745\,
            I => \N__77512\
        );

    \I__19527\ : InMux
    port map (
            O => \N__77744\,
            I => \N__77507\
        );

    \I__19526\ : InMux
    port map (
            O => \N__77743\,
            I => \N__77507\
        );

    \I__19525\ : LocalMux
    port map (
            O => \N__77740\,
            I => \N__77498\
        );

    \I__19524\ : Span4Mux_h
    port map (
            O => \N__77733\,
            I => \N__77498\
        );

    \I__19523\ : Span4Mux_h
    port map (
            O => \N__77730\,
            I => \N__77498\
        );

    \I__19522\ : LocalMux
    port map (
            O => \N__77723\,
            I => \N__77498\
        );

    \I__19521\ : LocalMux
    port map (
            O => \N__77720\,
            I => \N__77489\
        );

    \I__19520\ : LocalMux
    port map (
            O => \N__77715\,
            I => \N__77489\
        );

    \I__19519\ : LocalMux
    port map (
            O => \N__77708\,
            I => \N__77489\
        );

    \I__19518\ : LocalMux
    port map (
            O => \N__77701\,
            I => \N__77489\
        );

    \I__19517\ : InMux
    port map (
            O => \N__77700\,
            I => \N__77480\
        );

    \I__19516\ : InMux
    port map (
            O => \N__77697\,
            I => \N__77480\
        );

    \I__19515\ : InMux
    port map (
            O => \N__77694\,
            I => \N__77480\
        );

    \I__19514\ : InMux
    port map (
            O => \N__77693\,
            I => \N__77480\
        );

    \I__19513\ : InMux
    port map (
            O => \N__77692\,
            I => \N__77473\
        );

    \I__19512\ : InMux
    port map (
            O => \N__77691\,
            I => \N__77473\
        );

    \I__19511\ : InMux
    port map (
            O => \N__77690\,
            I => \N__77473\
        );

    \I__19510\ : InMux
    port map (
            O => \N__77689\,
            I => \N__77466\
        );

    \I__19509\ : InMux
    port map (
            O => \N__77688\,
            I => \N__77466\
        );

    \I__19508\ : InMux
    port map (
            O => \N__77685\,
            I => \N__77466\
        );

    \I__19507\ : LocalMux
    port map (
            O => \N__77682\,
            I => \N__77459\
        );

    \I__19506\ : LocalMux
    port map (
            O => \N__77675\,
            I => \N__77459\
        );

    \I__19505\ : LocalMux
    port map (
            O => \N__77668\,
            I => \N__77459\
        );

    \I__19504\ : LocalMux
    port map (
            O => \N__77659\,
            I => \N__77450\
        );

    \I__19503\ : LocalMux
    port map (
            O => \N__77654\,
            I => \N__77450\
        );

    \I__19502\ : LocalMux
    port map (
            O => \N__77647\,
            I => \N__77450\
        );

    \I__19501\ : LocalMux
    port map (
            O => \N__77642\,
            I => \N__77450\
        );

    \I__19500\ : Span4Mux_h
    port map (
            O => \N__77639\,
            I => \N__77441\
        );

    \I__19499\ : Span4Mux_v
    port map (
            O => \N__77636\,
            I => \N__77441\
        );

    \I__19498\ : LocalMux
    port map (
            O => \N__77627\,
            I => \N__77441\
        );

    \I__19497\ : LocalMux
    port map (
            O => \N__77624\,
            I => \N__77441\
        );

    \I__19496\ : Span12Mux_s11_h
    port map (
            O => \N__77621\,
            I => \N__77438\
        );

    \I__19495\ : InMux
    port map (
            O => \N__77620\,
            I => \N__77427\
        );

    \I__19494\ : InMux
    port map (
            O => \N__77619\,
            I => \N__77427\
        );

    \I__19493\ : InMux
    port map (
            O => \N__77618\,
            I => \N__77427\
        );

    \I__19492\ : InMux
    port map (
            O => \N__77617\,
            I => \N__77427\
        );

    \I__19491\ : InMux
    port map (
            O => \N__77616\,
            I => \N__77427\
        );

    \I__19490\ : InMux
    port map (
            O => \N__77615\,
            I => \N__77420\
        );

    \I__19489\ : InMux
    port map (
            O => \N__77614\,
            I => \N__77420\
        );

    \I__19488\ : InMux
    port map (
            O => \N__77613\,
            I => \N__77420\
        );

    \I__19487\ : InMux
    port map (
            O => \N__77612\,
            I => \N__77415\
        );

    \I__19486\ : InMux
    port map (
            O => \N__77611\,
            I => \N__77415\
        );

    \I__19485\ : InMux
    port map (
            O => \N__77610\,
            I => \N__77408\
        );

    \I__19484\ : InMux
    port map (
            O => \N__77609\,
            I => \N__77408\
        );

    \I__19483\ : InMux
    port map (
            O => \N__77608\,
            I => \N__77408\
        );

    \I__19482\ : Span4Mux_h
    port map (
            O => \N__77605\,
            I => \N__77401\
        );

    \I__19481\ : Span4Mux_h
    port map (
            O => \N__77598\,
            I => \N__77401\
        );

    \I__19480\ : LocalMux
    port map (
            O => \N__77591\,
            I => \N__77401\
        );

    \I__19479\ : InMux
    port map (
            O => \N__77590\,
            I => \N__77392\
        );

    \I__19478\ : InMux
    port map (
            O => \N__77587\,
            I => \N__77392\
        );

    \I__19477\ : InMux
    port map (
            O => \N__77584\,
            I => \N__77392\
        );

    \I__19476\ : InMux
    port map (
            O => \N__77583\,
            I => \N__77392\
        );

    \I__19475\ : InMux
    port map (
            O => \N__77580\,
            I => \N__77383\
        );

    \I__19474\ : InMux
    port map (
            O => \N__77577\,
            I => \N__77383\
        );

    \I__19473\ : InMux
    port map (
            O => \N__77576\,
            I => \N__77383\
        );

    \I__19472\ : InMux
    port map (
            O => \N__77575\,
            I => \N__77383\
        );

    \I__19471\ : Span4Mux_v
    port map (
            O => \N__77568\,
            I => \N__77378\
        );

    \I__19470\ : LocalMux
    port map (
            O => \N__77559\,
            I => \N__77378\
        );

    \I__19469\ : LocalMux
    port map (
            O => \N__77548\,
            I => \N__77373\
        );

    \I__19468\ : LocalMux
    port map (
            O => \N__77539\,
            I => \N__77373\
        );

    \I__19467\ : LocalMux
    port map (
            O => \N__77532\,
            I => \N__77366\
        );

    \I__19466\ : Span4Mux_h
    port map (
            O => \N__77525\,
            I => \N__77366\
        );

    \I__19465\ : Span4Mux_v
    port map (
            O => \N__77518\,
            I => \N__77366\
        );

    \I__19464\ : Span4Mux_v
    port map (
            O => \N__77515\,
            I => \N__77343\
        );

    \I__19463\ : Span4Mux_h
    port map (
            O => \N__77512\,
            I => \N__77343\
        );

    \I__19462\ : LocalMux
    port map (
            O => \N__77507\,
            I => \N__77343\
        );

    \I__19461\ : Span4Mux_v
    port map (
            O => \N__77498\,
            I => \N__77343\
        );

    \I__19460\ : Span4Mux_v
    port map (
            O => \N__77489\,
            I => \N__77343\
        );

    \I__19459\ : LocalMux
    port map (
            O => \N__77480\,
            I => \N__77343\
        );

    \I__19458\ : LocalMux
    port map (
            O => \N__77473\,
            I => \N__77343\
        );

    \I__19457\ : LocalMux
    port map (
            O => \N__77466\,
            I => \N__77343\
        );

    \I__19456\ : Span4Mux_v
    port map (
            O => \N__77459\,
            I => \N__77343\
        );

    \I__19455\ : Span4Mux_v
    port map (
            O => \N__77450\,
            I => \N__77343\
        );

    \I__19454\ : Span4Mux_h
    port map (
            O => \N__77441\,
            I => \N__77343\
        );

    \I__19453\ : Odrv12
    port map (
            O => \N__77438\,
            I => \progRomAddress_2\
        );

    \I__19452\ : LocalMux
    port map (
            O => \N__77427\,
            I => \progRomAddress_2\
        );

    \I__19451\ : LocalMux
    port map (
            O => \N__77420\,
            I => \progRomAddress_2\
        );

    \I__19450\ : LocalMux
    port map (
            O => \N__77415\,
            I => \progRomAddress_2\
        );

    \I__19449\ : LocalMux
    port map (
            O => \N__77408\,
            I => \progRomAddress_2\
        );

    \I__19448\ : Odrv4
    port map (
            O => \N__77401\,
            I => \progRomAddress_2\
        );

    \I__19447\ : LocalMux
    port map (
            O => \N__77392\,
            I => \progRomAddress_2\
        );

    \I__19446\ : LocalMux
    port map (
            O => \N__77383\,
            I => \progRomAddress_2\
        );

    \I__19445\ : Odrv4
    port map (
            O => \N__77378\,
            I => \progRomAddress_2\
        );

    \I__19444\ : Odrv4
    port map (
            O => \N__77373\,
            I => \progRomAddress_2\
        );

    \I__19443\ : Odrv4
    port map (
            O => \N__77366\,
            I => \progRomAddress_2\
        );

    \I__19442\ : Odrv4
    port map (
            O => \N__77343\,
            I => \progRomAddress_2\
        );

    \I__19441\ : InMux
    port map (
            O => \N__77318\,
            I => \N__77305\
        );

    \I__19440\ : InMux
    port map (
            O => \N__77317\,
            I => \N__77298\
        );

    \I__19439\ : InMux
    port map (
            O => \N__77316\,
            I => \N__77287\
        );

    \I__19438\ : InMux
    port map (
            O => \N__77315\,
            I => \N__77287\
        );

    \I__19437\ : CascadeMux
    port map (
            O => \N__77314\,
            I => \N__77284\
        );

    \I__19436\ : InMux
    port map (
            O => \N__77313\,
            I => \N__77275\
        );

    \I__19435\ : InMux
    port map (
            O => \N__77312\,
            I => \N__77275\
        );

    \I__19434\ : InMux
    port map (
            O => \N__77311\,
            I => \N__77268\
        );

    \I__19433\ : InMux
    port map (
            O => \N__77310\,
            I => \N__77265\
        );

    \I__19432\ : InMux
    port map (
            O => \N__77309\,
            I => \N__77262\
        );

    \I__19431\ : InMux
    port map (
            O => \N__77308\,
            I => \N__77259\
        );

    \I__19430\ : LocalMux
    port map (
            O => \N__77305\,
            I => \N__77231\
        );

    \I__19429\ : InMux
    port map (
            O => \N__77304\,
            I => \N__77222\
        );

    \I__19428\ : InMux
    port map (
            O => \N__77303\,
            I => \N__77222\
        );

    \I__19427\ : InMux
    port map (
            O => \N__77302\,
            I => \N__77222\
        );

    \I__19426\ : InMux
    port map (
            O => \N__77301\,
            I => \N__77222\
        );

    \I__19425\ : LocalMux
    port map (
            O => \N__77298\,
            I => \N__77219\
        );

    \I__19424\ : InMux
    port map (
            O => \N__77297\,
            I => \N__77214\
        );

    \I__19423\ : InMux
    port map (
            O => \N__77296\,
            I => \N__77214\
        );

    \I__19422\ : InMux
    port map (
            O => \N__77295\,
            I => \N__77205\
        );

    \I__19421\ : InMux
    port map (
            O => \N__77294\,
            I => \N__77205\
        );

    \I__19420\ : InMux
    port map (
            O => \N__77293\,
            I => \N__77205\
        );

    \I__19419\ : InMux
    port map (
            O => \N__77292\,
            I => \N__77205\
        );

    \I__19418\ : LocalMux
    port map (
            O => \N__77287\,
            I => \N__77202\
        );

    \I__19417\ : InMux
    port map (
            O => \N__77284\,
            I => \N__77193\
        );

    \I__19416\ : InMux
    port map (
            O => \N__77283\,
            I => \N__77176\
        );

    \I__19415\ : InMux
    port map (
            O => \N__77282\,
            I => \N__77176\
        );

    \I__19414\ : InMux
    port map (
            O => \N__77281\,
            I => \N__77166\
        );

    \I__19413\ : InMux
    port map (
            O => \N__77280\,
            I => \N__77166\
        );

    \I__19412\ : LocalMux
    port map (
            O => \N__77275\,
            I => \N__77161\
        );

    \I__19411\ : InMux
    port map (
            O => \N__77274\,
            I => \N__77152\
        );

    \I__19410\ : InMux
    port map (
            O => \N__77273\,
            I => \N__77152\
        );

    \I__19409\ : InMux
    port map (
            O => \N__77272\,
            I => \N__77152\
        );

    \I__19408\ : InMux
    port map (
            O => \N__77271\,
            I => \N__77152\
        );

    \I__19407\ : LocalMux
    port map (
            O => \N__77268\,
            I => \N__77137\
        );

    \I__19406\ : LocalMux
    port map (
            O => \N__77265\,
            I => \N__77132\
        );

    \I__19405\ : LocalMux
    port map (
            O => \N__77262\,
            I => \N__77132\
        );

    \I__19404\ : LocalMux
    port map (
            O => \N__77259\,
            I => \N__77129\
        );

    \I__19403\ : InMux
    port map (
            O => \N__77258\,
            I => \N__77126\
        );

    \I__19402\ : InMux
    port map (
            O => \N__77257\,
            I => \N__77109\
        );

    \I__19401\ : InMux
    port map (
            O => \N__77256\,
            I => \N__77109\
        );

    \I__19400\ : InMux
    port map (
            O => \N__77255\,
            I => \N__77100\
        );

    \I__19399\ : InMux
    port map (
            O => \N__77254\,
            I => \N__77100\
        );

    \I__19398\ : InMux
    port map (
            O => \N__77253\,
            I => \N__77100\
        );

    \I__19397\ : InMux
    port map (
            O => \N__77252\,
            I => \N__77100\
        );

    \I__19396\ : InMux
    port map (
            O => \N__77251\,
            I => \N__77093\
        );

    \I__19395\ : InMux
    port map (
            O => \N__77250\,
            I => \N__77093\
        );

    \I__19394\ : InMux
    port map (
            O => \N__77249\,
            I => \N__77093\
        );

    \I__19393\ : InMux
    port map (
            O => \N__77248\,
            I => \N__77088\
        );

    \I__19392\ : InMux
    port map (
            O => \N__77247\,
            I => \N__77088\
        );

    \I__19391\ : InMux
    port map (
            O => \N__77246\,
            I => \N__77081\
        );

    \I__19390\ : InMux
    port map (
            O => \N__77245\,
            I => \N__77081\
        );

    \I__19389\ : InMux
    port map (
            O => \N__77244\,
            I => \N__77081\
        );

    \I__19388\ : InMux
    port map (
            O => \N__77243\,
            I => \N__77074\
        );

    \I__19387\ : InMux
    port map (
            O => \N__77242\,
            I => \N__77074\
        );

    \I__19386\ : InMux
    port map (
            O => \N__77241\,
            I => \N__77074\
        );

    \I__19385\ : InMux
    port map (
            O => \N__77240\,
            I => \N__77062\
        );

    \I__19384\ : InMux
    port map (
            O => \N__77239\,
            I => \N__77055\
        );

    \I__19383\ : InMux
    port map (
            O => \N__77238\,
            I => \N__77055\
        );

    \I__19382\ : InMux
    port map (
            O => \N__77237\,
            I => \N__77055\
        );

    \I__19381\ : InMux
    port map (
            O => \N__77236\,
            I => \N__77048\
        );

    \I__19380\ : InMux
    port map (
            O => \N__77235\,
            I => \N__77048\
        );

    \I__19379\ : InMux
    port map (
            O => \N__77234\,
            I => \N__77048\
        );

    \I__19378\ : Span4Mux_h
    port map (
            O => \N__77231\,
            I => \N__77039\
        );

    \I__19377\ : LocalMux
    port map (
            O => \N__77222\,
            I => \N__77039\
        );

    \I__19376\ : Span4Mux_v
    port map (
            O => \N__77219\,
            I => \N__77039\
        );

    \I__19375\ : LocalMux
    port map (
            O => \N__77214\,
            I => \N__77039\
        );

    \I__19374\ : LocalMux
    port map (
            O => \N__77205\,
            I => \N__77034\
        );

    \I__19373\ : Span4Mux_v
    port map (
            O => \N__77202\,
            I => \N__77034\
        );

    \I__19372\ : InMux
    port map (
            O => \N__77201\,
            I => \N__77027\
        );

    \I__19371\ : InMux
    port map (
            O => \N__77200\,
            I => \N__77027\
        );

    \I__19370\ : InMux
    port map (
            O => \N__77199\,
            I => \N__77027\
        );

    \I__19369\ : InMux
    port map (
            O => \N__77198\,
            I => \N__77020\
        );

    \I__19368\ : InMux
    port map (
            O => \N__77197\,
            I => \N__77020\
        );

    \I__19367\ : InMux
    port map (
            O => \N__77196\,
            I => \N__77020\
        );

    \I__19366\ : LocalMux
    port map (
            O => \N__77193\,
            I => \N__77017\
        );

    \I__19365\ : InMux
    port map (
            O => \N__77192\,
            I => \N__77010\
        );

    \I__19364\ : InMux
    port map (
            O => \N__77191\,
            I => \N__77010\
        );

    \I__19363\ : InMux
    port map (
            O => \N__77190\,
            I => \N__77010\
        );

    \I__19362\ : InMux
    port map (
            O => \N__77189\,
            I => \N__77003\
        );

    \I__19361\ : InMux
    port map (
            O => \N__77188\,
            I => \N__77003\
        );

    \I__19360\ : InMux
    port map (
            O => \N__77187\,
            I => \N__77003\
        );

    \I__19359\ : InMux
    port map (
            O => \N__77186\,
            I => \N__76998\
        );

    \I__19358\ : InMux
    port map (
            O => \N__77185\,
            I => \N__76998\
        );

    \I__19357\ : InMux
    port map (
            O => \N__77184\,
            I => \N__76995\
        );

    \I__19356\ : InMux
    port map (
            O => \N__77183\,
            I => \N__76988\
        );

    \I__19355\ : InMux
    port map (
            O => \N__77182\,
            I => \N__76988\
        );

    \I__19354\ : InMux
    port map (
            O => \N__77181\,
            I => \N__76988\
        );

    \I__19353\ : LocalMux
    port map (
            O => \N__77176\,
            I => \N__76985\
        );

    \I__19352\ : InMux
    port map (
            O => \N__77175\,
            I => \N__76982\
        );

    \I__19351\ : InMux
    port map (
            O => \N__77174\,
            I => \N__76979\
        );

    \I__19350\ : InMux
    port map (
            O => \N__77173\,
            I => \N__76970\
        );

    \I__19349\ : InMux
    port map (
            O => \N__77172\,
            I => \N__76970\
        );

    \I__19348\ : InMux
    port map (
            O => \N__77171\,
            I => \N__76970\
        );

    \I__19347\ : LocalMux
    port map (
            O => \N__77166\,
            I => \N__76967\
        );

    \I__19346\ : InMux
    port map (
            O => \N__77165\,
            I => \N__76960\
        );

    \I__19345\ : InMux
    port map (
            O => \N__77164\,
            I => \N__76960\
        );

    \I__19344\ : Span4Mux_v
    port map (
            O => \N__77161\,
            I => \N__76957\
        );

    \I__19343\ : LocalMux
    port map (
            O => \N__77152\,
            I => \N__76954\
        );

    \I__19342\ : InMux
    port map (
            O => \N__77151\,
            I => \N__76947\
        );

    \I__19341\ : InMux
    port map (
            O => \N__77150\,
            I => \N__76947\
        );

    \I__19340\ : InMux
    port map (
            O => \N__77149\,
            I => \N__76947\
        );

    \I__19339\ : InMux
    port map (
            O => \N__77148\,
            I => \N__76938\
        );

    \I__19338\ : InMux
    port map (
            O => \N__77147\,
            I => \N__76938\
        );

    \I__19337\ : InMux
    port map (
            O => \N__77146\,
            I => \N__76938\
        );

    \I__19336\ : InMux
    port map (
            O => \N__77145\,
            I => \N__76938\
        );

    \I__19335\ : InMux
    port map (
            O => \N__77144\,
            I => \N__76914\
        );

    \I__19334\ : InMux
    port map (
            O => \N__77143\,
            I => \N__76914\
        );

    \I__19333\ : InMux
    port map (
            O => \N__77142\,
            I => \N__76914\
        );

    \I__19332\ : InMux
    port map (
            O => \N__77141\,
            I => \N__76914\
        );

    \I__19331\ : InMux
    port map (
            O => \N__77140\,
            I => \N__76914\
        );

    \I__19330\ : Span4Mux_h
    port map (
            O => \N__77137\,
            I => \N__76904\
        );

    \I__19329\ : Span4Mux_v
    port map (
            O => \N__77132\,
            I => \N__76904\
        );

    \I__19328\ : Span4Mux_h
    port map (
            O => \N__77129\,
            I => \N__76899\
        );

    \I__19327\ : LocalMux
    port map (
            O => \N__77126\,
            I => \N__76899\
        );

    \I__19326\ : InMux
    port map (
            O => \N__77125\,
            I => \N__76890\
        );

    \I__19325\ : InMux
    port map (
            O => \N__77124\,
            I => \N__76890\
        );

    \I__19324\ : InMux
    port map (
            O => \N__77123\,
            I => \N__76890\
        );

    \I__19323\ : InMux
    port map (
            O => \N__77122\,
            I => \N__76890\
        );

    \I__19322\ : InMux
    port map (
            O => \N__77121\,
            I => \N__76879\
        );

    \I__19321\ : InMux
    port map (
            O => \N__77120\,
            I => \N__76879\
        );

    \I__19320\ : InMux
    port map (
            O => \N__77119\,
            I => \N__76879\
        );

    \I__19319\ : InMux
    port map (
            O => \N__77118\,
            I => \N__76879\
        );

    \I__19318\ : InMux
    port map (
            O => \N__77117\,
            I => \N__76879\
        );

    \I__19317\ : InMux
    port map (
            O => \N__77116\,
            I => \N__76872\
        );

    \I__19316\ : InMux
    port map (
            O => \N__77115\,
            I => \N__76872\
        );

    \I__19315\ : InMux
    port map (
            O => \N__77114\,
            I => \N__76872\
        );

    \I__19314\ : LocalMux
    port map (
            O => \N__77109\,
            I => \N__76865\
        );

    \I__19313\ : LocalMux
    port map (
            O => \N__77100\,
            I => \N__76865\
        );

    \I__19312\ : LocalMux
    port map (
            O => \N__77093\,
            I => \N__76865\
        );

    \I__19311\ : LocalMux
    port map (
            O => \N__77088\,
            I => \N__76858\
        );

    \I__19310\ : LocalMux
    port map (
            O => \N__77081\,
            I => \N__76858\
        );

    \I__19309\ : LocalMux
    port map (
            O => \N__77074\,
            I => \N__76858\
        );

    \I__19308\ : InMux
    port map (
            O => \N__77073\,
            I => \N__76851\
        );

    \I__19307\ : InMux
    port map (
            O => \N__77072\,
            I => \N__76851\
        );

    \I__19306\ : InMux
    port map (
            O => \N__77071\,
            I => \N__76851\
        );

    \I__19305\ : InMux
    port map (
            O => \N__77070\,
            I => \N__76838\
        );

    \I__19304\ : InMux
    port map (
            O => \N__77069\,
            I => \N__76838\
        );

    \I__19303\ : InMux
    port map (
            O => \N__77068\,
            I => \N__76838\
        );

    \I__19302\ : InMux
    port map (
            O => \N__77067\,
            I => \N__76838\
        );

    \I__19301\ : InMux
    port map (
            O => \N__77066\,
            I => \N__76838\
        );

    \I__19300\ : InMux
    port map (
            O => \N__77065\,
            I => \N__76838\
        );

    \I__19299\ : LocalMux
    port map (
            O => \N__77062\,
            I => \N__76831\
        );

    \I__19298\ : LocalMux
    port map (
            O => \N__77055\,
            I => \N__76831\
        );

    \I__19297\ : LocalMux
    port map (
            O => \N__77048\,
            I => \N__76831\
        );

    \I__19296\ : Span4Mux_h
    port map (
            O => \N__77039\,
            I => \N__76822\
        );

    \I__19295\ : Span4Mux_h
    port map (
            O => \N__77034\,
            I => \N__76822\
        );

    \I__19294\ : LocalMux
    port map (
            O => \N__77027\,
            I => \N__76822\
        );

    \I__19293\ : LocalMux
    port map (
            O => \N__77020\,
            I => \N__76822\
        );

    \I__19292\ : Span4Mux_v
    port map (
            O => \N__77017\,
            I => \N__76811\
        );

    \I__19291\ : LocalMux
    port map (
            O => \N__77010\,
            I => \N__76811\
        );

    \I__19290\ : LocalMux
    port map (
            O => \N__77003\,
            I => \N__76811\
        );

    \I__19289\ : LocalMux
    port map (
            O => \N__76998\,
            I => \N__76811\
        );

    \I__19288\ : LocalMux
    port map (
            O => \N__76995\,
            I => \N__76811\
        );

    \I__19287\ : LocalMux
    port map (
            O => \N__76988\,
            I => \N__76802\
        );

    \I__19286\ : Span4Mux_v
    port map (
            O => \N__76985\,
            I => \N__76802\
        );

    \I__19285\ : LocalMux
    port map (
            O => \N__76982\,
            I => \N__76802\
        );

    \I__19284\ : LocalMux
    port map (
            O => \N__76979\,
            I => \N__76802\
        );

    \I__19283\ : InMux
    port map (
            O => \N__76978\,
            I => \N__76797\
        );

    \I__19282\ : InMux
    port map (
            O => \N__76977\,
            I => \N__76797\
        );

    \I__19281\ : LocalMux
    port map (
            O => \N__76970\,
            I => \N__76792\
        );

    \I__19280\ : Span12Mux_s10_v
    port map (
            O => \N__76967\,
            I => \N__76792\
        );

    \I__19279\ : InMux
    port map (
            O => \N__76966\,
            I => \N__76787\
        );

    \I__19278\ : InMux
    port map (
            O => \N__76965\,
            I => \N__76787\
        );

    \I__19277\ : LocalMux
    port map (
            O => \N__76960\,
            I => \N__76784\
        );

    \I__19276\ : Span4Mux_h
    port map (
            O => \N__76957\,
            I => \N__76775\
        );

    \I__19275\ : Span4Mux_v
    port map (
            O => \N__76954\,
            I => \N__76775\
        );

    \I__19274\ : LocalMux
    port map (
            O => \N__76947\,
            I => \N__76775\
        );

    \I__19273\ : LocalMux
    port map (
            O => \N__76938\,
            I => \N__76775\
        );

    \I__19272\ : InMux
    port map (
            O => \N__76937\,
            I => \N__76762\
        );

    \I__19271\ : InMux
    port map (
            O => \N__76936\,
            I => \N__76762\
        );

    \I__19270\ : InMux
    port map (
            O => \N__76935\,
            I => \N__76762\
        );

    \I__19269\ : InMux
    port map (
            O => \N__76934\,
            I => \N__76762\
        );

    \I__19268\ : InMux
    port map (
            O => \N__76933\,
            I => \N__76762\
        );

    \I__19267\ : InMux
    port map (
            O => \N__76932\,
            I => \N__76762\
        );

    \I__19266\ : InMux
    port map (
            O => \N__76931\,
            I => \N__76753\
        );

    \I__19265\ : InMux
    port map (
            O => \N__76930\,
            I => \N__76753\
        );

    \I__19264\ : InMux
    port map (
            O => \N__76929\,
            I => \N__76753\
        );

    \I__19263\ : InMux
    port map (
            O => \N__76928\,
            I => \N__76753\
        );

    \I__19262\ : InMux
    port map (
            O => \N__76927\,
            I => \N__76746\
        );

    \I__19261\ : InMux
    port map (
            O => \N__76926\,
            I => \N__76746\
        );

    \I__19260\ : InMux
    port map (
            O => \N__76925\,
            I => \N__76746\
        );

    \I__19259\ : LocalMux
    port map (
            O => \N__76914\,
            I => \N__76743\
        );

    \I__19258\ : InMux
    port map (
            O => \N__76913\,
            I => \N__76732\
        );

    \I__19257\ : InMux
    port map (
            O => \N__76912\,
            I => \N__76732\
        );

    \I__19256\ : InMux
    port map (
            O => \N__76911\,
            I => \N__76732\
        );

    \I__19255\ : InMux
    port map (
            O => \N__76910\,
            I => \N__76732\
        );

    \I__19254\ : InMux
    port map (
            O => \N__76909\,
            I => \N__76732\
        );

    \I__19253\ : Span4Mux_h
    port map (
            O => \N__76904\,
            I => \N__76723\
        );

    \I__19252\ : Span4Mux_h
    port map (
            O => \N__76899\,
            I => \N__76723\
        );

    \I__19251\ : LocalMux
    port map (
            O => \N__76890\,
            I => \N__76723\
        );

    \I__19250\ : LocalMux
    port map (
            O => \N__76879\,
            I => \N__76723\
        );

    \I__19249\ : LocalMux
    port map (
            O => \N__76872\,
            I => \N__76704\
        );

    \I__19248\ : Span4Mux_v
    port map (
            O => \N__76865\,
            I => \N__76704\
        );

    \I__19247\ : Span4Mux_v
    port map (
            O => \N__76858\,
            I => \N__76704\
        );

    \I__19246\ : LocalMux
    port map (
            O => \N__76851\,
            I => \N__76704\
        );

    \I__19245\ : LocalMux
    port map (
            O => \N__76838\,
            I => \N__76704\
        );

    \I__19244\ : Span4Mux_v
    port map (
            O => \N__76831\,
            I => \N__76704\
        );

    \I__19243\ : Span4Mux_v
    port map (
            O => \N__76822\,
            I => \N__76704\
        );

    \I__19242\ : Span4Mux_v
    port map (
            O => \N__76811\,
            I => \N__76704\
        );

    \I__19241\ : Span4Mux_h
    port map (
            O => \N__76802\,
            I => \N__76704\
        );

    \I__19240\ : LocalMux
    port map (
            O => \N__76797\,
            I => \progRomAddress_0\
        );

    \I__19239\ : Odrv12
    port map (
            O => \N__76792\,
            I => \progRomAddress_0\
        );

    \I__19238\ : LocalMux
    port map (
            O => \N__76787\,
            I => \progRomAddress_0\
        );

    \I__19237\ : Odrv4
    port map (
            O => \N__76784\,
            I => \progRomAddress_0\
        );

    \I__19236\ : Odrv4
    port map (
            O => \N__76775\,
            I => \progRomAddress_0\
        );

    \I__19235\ : LocalMux
    port map (
            O => \N__76762\,
            I => \progRomAddress_0\
        );

    \I__19234\ : LocalMux
    port map (
            O => \N__76753\,
            I => \progRomAddress_0\
        );

    \I__19233\ : LocalMux
    port map (
            O => \N__76746\,
            I => \progRomAddress_0\
        );

    \I__19232\ : Odrv4
    port map (
            O => \N__76743\,
            I => \progRomAddress_0\
        );

    \I__19231\ : LocalMux
    port map (
            O => \N__76732\,
            I => \progRomAddress_0\
        );

    \I__19230\ : Odrv4
    port map (
            O => \N__76723\,
            I => \progRomAddress_0\
        );

    \I__19229\ : Odrv4
    port map (
            O => \N__76704\,
            I => \progRomAddress_0\
        );

    \I__19228\ : InMux
    port map (
            O => \N__76679\,
            I => \N__76676\
        );

    \I__19227\ : LocalMux
    port map (
            O => \N__76676\,
            I => \N__76673\
        );

    \I__19226\ : Span4Mux_v
    port map (
            O => \N__76673\,
            I => \N__76670\
        );

    \I__19225\ : Span4Mux_h
    port map (
            O => \N__76670\,
            I => \N__76667\
        );

    \I__19224\ : Odrv4
    port map (
            O => \N__76667\,
            I => \PROM.ROMDATA.m338_bm\
        );

    \I__19223\ : CascadeMux
    port map (
            O => \N__76664\,
            I => \PROM.ROMDATA.m338_am_cascade_\
        );

    \I__19222\ : InMux
    port map (
            O => \N__76661\,
            I => \N__76658\
        );

    \I__19221\ : LocalMux
    port map (
            O => \N__76658\,
            I => \PROM.ROMDATA.m338_ns\
        );

    \I__19220\ : InMux
    port map (
            O => \N__76655\,
            I => \N__76652\
        );

    \I__19219\ : LocalMux
    port map (
            O => \N__76652\,
            I => \N__76649\
        );

    \I__19218\ : Span4Mux_h
    port map (
            O => \N__76649\,
            I => \N__76645\
        );

    \I__19217\ : InMux
    port map (
            O => \N__76648\,
            I => \N__76642\
        );

    \I__19216\ : Odrv4
    port map (
            O => \N__76645\,
            I => \PROM.ROMDATA.m246\
        );

    \I__19215\ : LocalMux
    port map (
            O => \N__76642\,
            I => \PROM.ROMDATA.m246\
        );

    \I__19214\ : InMux
    port map (
            O => \N__76637\,
            I => \N__76626\
        );

    \I__19213\ : InMux
    port map (
            O => \N__76636\,
            I => \N__76626\
        );

    \I__19212\ : InMux
    port map (
            O => \N__76635\,
            I => \N__76626\
        );

    \I__19211\ : CascadeMux
    port map (
            O => \N__76634\,
            I => \N__76620\
        );

    \I__19210\ : InMux
    port map (
            O => \N__76633\,
            I => \N__76613\
        );

    \I__19209\ : LocalMux
    port map (
            O => \N__76626\,
            I => \N__76610\
        );

    \I__19208\ : InMux
    port map (
            O => \N__76625\,
            I => \N__76597\
        );

    \I__19207\ : InMux
    port map (
            O => \N__76624\,
            I => \N__76594\
        );

    \I__19206\ : CascadeMux
    port map (
            O => \N__76623\,
            I => \N__76588\
        );

    \I__19205\ : InMux
    port map (
            O => \N__76620\,
            I => \N__76580\
        );

    \I__19204\ : CascadeMux
    port map (
            O => \N__76619\,
            I => \N__76576\
        );

    \I__19203\ : InMux
    port map (
            O => \N__76618\,
            I => \N__76566\
        );

    \I__19202\ : InMux
    port map (
            O => \N__76617\,
            I => \N__76563\
        );

    \I__19201\ : CascadeMux
    port map (
            O => \N__76616\,
            I => \N__76560\
        );

    \I__19200\ : LocalMux
    port map (
            O => \N__76613\,
            I => \N__76554\
        );

    \I__19199\ : Span4Mux_v
    port map (
            O => \N__76610\,
            I => \N__76554\
        );

    \I__19198\ : InMux
    port map (
            O => \N__76609\,
            I => \N__76551\
        );

    \I__19197\ : InMux
    port map (
            O => \N__76608\,
            I => \N__76546\
        );

    \I__19196\ : InMux
    port map (
            O => \N__76607\,
            I => \N__76546\
        );

    \I__19195\ : InMux
    port map (
            O => \N__76606\,
            I => \N__76541\
        );

    \I__19194\ : InMux
    port map (
            O => \N__76605\,
            I => \N__76541\
        );

    \I__19193\ : InMux
    port map (
            O => \N__76604\,
            I => \N__76536\
        );

    \I__19192\ : InMux
    port map (
            O => \N__76603\,
            I => \N__76536\
        );

    \I__19191\ : CascadeMux
    port map (
            O => \N__76602\,
            I => \N__76523\
        );

    \I__19190\ : CascadeMux
    port map (
            O => \N__76601\,
            I => \N__76519\
        );

    \I__19189\ : InMux
    port map (
            O => \N__76600\,
            I => \N__76516\
        );

    \I__19188\ : LocalMux
    port map (
            O => \N__76597\,
            I => \N__76513\
        );

    \I__19187\ : LocalMux
    port map (
            O => \N__76594\,
            I => \N__76510\
        );

    \I__19186\ : InMux
    port map (
            O => \N__76593\,
            I => \N__76507\
        );

    \I__19185\ : InMux
    port map (
            O => \N__76592\,
            I => \N__76504\
        );

    \I__19184\ : InMux
    port map (
            O => \N__76591\,
            I => \N__76501\
        );

    \I__19183\ : InMux
    port map (
            O => \N__76588\,
            I => \N__76493\
        );

    \I__19182\ : InMux
    port map (
            O => \N__76587\,
            I => \N__76493\
        );

    \I__19181\ : InMux
    port map (
            O => \N__76586\,
            I => \N__76486\
        );

    \I__19180\ : InMux
    port map (
            O => \N__76585\,
            I => \N__76486\
        );

    \I__19179\ : InMux
    port map (
            O => \N__76584\,
            I => \N__76486\
        );

    \I__19178\ : InMux
    port map (
            O => \N__76583\,
            I => \N__76476\
        );

    \I__19177\ : LocalMux
    port map (
            O => \N__76580\,
            I => \N__76467\
        );

    \I__19176\ : CascadeMux
    port map (
            O => \N__76579\,
            I => \N__76464\
        );

    \I__19175\ : InMux
    port map (
            O => \N__76576\,
            I => \N__76455\
        );

    \I__19174\ : InMux
    port map (
            O => \N__76575\,
            I => \N__76449\
        );

    \I__19173\ : InMux
    port map (
            O => \N__76574\,
            I => \N__76449\
        );

    \I__19172\ : InMux
    port map (
            O => \N__76573\,
            I => \N__76441\
        );

    \I__19171\ : InMux
    port map (
            O => \N__76572\,
            I => \N__76441\
        );

    \I__19170\ : InMux
    port map (
            O => \N__76571\,
            I => \N__76434\
        );

    \I__19169\ : InMux
    port map (
            O => \N__76570\,
            I => \N__76434\
        );

    \I__19168\ : InMux
    port map (
            O => \N__76569\,
            I => \N__76434\
        );

    \I__19167\ : LocalMux
    port map (
            O => \N__76566\,
            I => \N__76429\
        );

    \I__19166\ : LocalMux
    port map (
            O => \N__76563\,
            I => \N__76429\
        );

    \I__19165\ : InMux
    port map (
            O => \N__76560\,
            I => \N__76424\
        );

    \I__19164\ : InMux
    port map (
            O => \N__76559\,
            I => \N__76424\
        );

    \I__19163\ : Span4Mux_h
    port map (
            O => \N__76554\,
            I => \N__76421\
        );

    \I__19162\ : LocalMux
    port map (
            O => \N__76551\,
            I => \N__76414\
        );

    \I__19161\ : LocalMux
    port map (
            O => \N__76546\,
            I => \N__76414\
        );

    \I__19160\ : LocalMux
    port map (
            O => \N__76541\,
            I => \N__76414\
        );

    \I__19159\ : LocalMux
    port map (
            O => \N__76536\,
            I => \N__76411\
        );

    \I__19158\ : InMux
    port map (
            O => \N__76535\,
            I => \N__76406\
        );

    \I__19157\ : InMux
    port map (
            O => \N__76534\,
            I => \N__76406\
        );

    \I__19156\ : InMux
    port map (
            O => \N__76533\,
            I => \N__76396\
        );

    \I__19155\ : InMux
    port map (
            O => \N__76532\,
            I => \N__76396\
        );

    \I__19154\ : InMux
    port map (
            O => \N__76531\,
            I => \N__76396\
        );

    \I__19153\ : InMux
    port map (
            O => \N__76530\,
            I => \N__76391\
        );

    \I__19152\ : InMux
    port map (
            O => \N__76529\,
            I => \N__76391\
        );

    \I__19151\ : InMux
    port map (
            O => \N__76528\,
            I => \N__76388\
        );

    \I__19150\ : InMux
    port map (
            O => \N__76527\,
            I => \N__76381\
        );

    \I__19149\ : InMux
    port map (
            O => \N__76526\,
            I => \N__76381\
        );

    \I__19148\ : InMux
    port map (
            O => \N__76523\,
            I => \N__76381\
        );

    \I__19147\ : InMux
    port map (
            O => \N__76522\,
            I => \N__76378\
        );

    \I__19146\ : InMux
    port map (
            O => \N__76519\,
            I => \N__76375\
        );

    \I__19145\ : LocalMux
    port map (
            O => \N__76516\,
            I => \N__76369\
        );

    \I__19144\ : Span4Mux_h
    port map (
            O => \N__76513\,
            I => \N__76362\
        );

    \I__19143\ : Span4Mux_v
    port map (
            O => \N__76510\,
            I => \N__76362\
        );

    \I__19142\ : LocalMux
    port map (
            O => \N__76507\,
            I => \N__76362\
        );

    \I__19141\ : LocalMux
    port map (
            O => \N__76504\,
            I => \N__76357\
        );

    \I__19140\ : LocalMux
    port map (
            O => \N__76501\,
            I => \N__76357\
        );

    \I__19139\ : InMux
    port map (
            O => \N__76500\,
            I => \N__76354\
        );

    \I__19138\ : InMux
    port map (
            O => \N__76499\,
            I => \N__76351\
        );

    \I__19137\ : CascadeMux
    port map (
            O => \N__76498\,
            I => \N__76346\
        );

    \I__19136\ : LocalMux
    port map (
            O => \N__76493\,
            I => \N__76341\
        );

    \I__19135\ : LocalMux
    port map (
            O => \N__76486\,
            I => \N__76341\
        );

    \I__19134\ : InMux
    port map (
            O => \N__76485\,
            I => \N__76336\
        );

    \I__19133\ : InMux
    port map (
            O => \N__76484\,
            I => \N__76336\
        );

    \I__19132\ : InMux
    port map (
            O => \N__76483\,
            I => \N__76331\
        );

    \I__19131\ : InMux
    port map (
            O => \N__76482\,
            I => \N__76331\
        );

    \I__19130\ : InMux
    port map (
            O => \N__76481\,
            I => \N__76326\
        );

    \I__19129\ : InMux
    port map (
            O => \N__76480\,
            I => \N__76326\
        );

    \I__19128\ : InMux
    port map (
            O => \N__76479\,
            I => \N__76323\
        );

    \I__19127\ : LocalMux
    port map (
            O => \N__76476\,
            I => \N__76318\
        );

    \I__19126\ : InMux
    port map (
            O => \N__76475\,
            I => \N__76313\
        );

    \I__19125\ : InMux
    port map (
            O => \N__76474\,
            I => \N__76313\
        );

    \I__19124\ : InMux
    port map (
            O => \N__76473\,
            I => \N__76310\
        );

    \I__19123\ : InMux
    port map (
            O => \N__76472\,
            I => \N__76305\
        );

    \I__19122\ : InMux
    port map (
            O => \N__76471\,
            I => \N__76305\
        );

    \I__19121\ : InMux
    port map (
            O => \N__76470\,
            I => \N__76302\
        );

    \I__19120\ : Span4Mux_h
    port map (
            O => \N__76467\,
            I => \N__76299\
        );

    \I__19119\ : InMux
    port map (
            O => \N__76464\,
            I => \N__76294\
        );

    \I__19118\ : InMux
    port map (
            O => \N__76463\,
            I => \N__76294\
        );

    \I__19117\ : CascadeMux
    port map (
            O => \N__76462\,
            I => \N__76288\
        );

    \I__19116\ : InMux
    port map (
            O => \N__76461\,
            I => \N__76277\
        );

    \I__19115\ : InMux
    port map (
            O => \N__76460\,
            I => \N__76277\
        );

    \I__19114\ : InMux
    port map (
            O => \N__76459\,
            I => \N__76277\
        );

    \I__19113\ : InMux
    port map (
            O => \N__76458\,
            I => \N__76277\
        );

    \I__19112\ : LocalMux
    port map (
            O => \N__76455\,
            I => \N__76274\
        );

    \I__19111\ : CascadeMux
    port map (
            O => \N__76454\,
            I => \N__76265\
        );

    \I__19110\ : LocalMux
    port map (
            O => \N__76449\,
            I => \N__76258\
        );

    \I__19109\ : InMux
    port map (
            O => \N__76448\,
            I => \N__76251\
        );

    \I__19108\ : InMux
    port map (
            O => \N__76447\,
            I => \N__76251\
        );

    \I__19107\ : InMux
    port map (
            O => \N__76446\,
            I => \N__76251\
        );

    \I__19106\ : LocalMux
    port map (
            O => \N__76441\,
            I => \N__76248\
        );

    \I__19105\ : LocalMux
    port map (
            O => \N__76434\,
            I => \N__76241\
        );

    \I__19104\ : Span4Mux_v
    port map (
            O => \N__76429\,
            I => \N__76241\
        );

    \I__19103\ : LocalMux
    port map (
            O => \N__76424\,
            I => \N__76241\
        );

    \I__19102\ : Span4Mux_h
    port map (
            O => \N__76421\,
            I => \N__76232\
        );

    \I__19101\ : Span4Mux_v
    port map (
            O => \N__76414\,
            I => \N__76232\
        );

    \I__19100\ : Span4Mux_v
    port map (
            O => \N__76411\,
            I => \N__76232\
        );

    \I__19099\ : LocalMux
    port map (
            O => \N__76406\,
            I => \N__76232\
        );

    \I__19098\ : InMux
    port map (
            O => \N__76405\,
            I => \N__76225\
        );

    \I__19097\ : InMux
    port map (
            O => \N__76404\,
            I => \N__76225\
        );

    \I__19096\ : InMux
    port map (
            O => \N__76403\,
            I => \N__76225\
        );

    \I__19095\ : LocalMux
    port map (
            O => \N__76396\,
            I => \N__76222\
        );

    \I__19094\ : LocalMux
    port map (
            O => \N__76391\,
            I => \N__76215\
        );

    \I__19093\ : LocalMux
    port map (
            O => \N__76388\,
            I => \N__76215\
        );

    \I__19092\ : LocalMux
    port map (
            O => \N__76381\,
            I => \N__76215\
        );

    \I__19091\ : LocalMux
    port map (
            O => \N__76378\,
            I => \N__76210\
        );

    \I__19090\ : LocalMux
    port map (
            O => \N__76375\,
            I => \N__76210\
        );

    \I__19089\ : InMux
    port map (
            O => \N__76374\,
            I => \N__76203\
        );

    \I__19088\ : InMux
    port map (
            O => \N__76373\,
            I => \N__76203\
        );

    \I__19087\ : InMux
    port map (
            O => \N__76372\,
            I => \N__76203\
        );

    \I__19086\ : Span4Mux_v
    port map (
            O => \N__76369\,
            I => \N__76192\
        );

    \I__19085\ : Span4Mux_h
    port map (
            O => \N__76362\,
            I => \N__76192\
        );

    \I__19084\ : Span4Mux_v
    port map (
            O => \N__76357\,
            I => \N__76192\
        );

    \I__19083\ : LocalMux
    port map (
            O => \N__76354\,
            I => \N__76192\
        );

    \I__19082\ : LocalMux
    port map (
            O => \N__76351\,
            I => \N__76192\
        );

    \I__19081\ : InMux
    port map (
            O => \N__76350\,
            I => \N__76185\
        );

    \I__19080\ : InMux
    port map (
            O => \N__76349\,
            I => \N__76185\
        );

    \I__19079\ : InMux
    port map (
            O => \N__76346\,
            I => \N__76185\
        );

    \I__19078\ : Span4Mux_h
    port map (
            O => \N__76341\,
            I => \N__76174\
        );

    \I__19077\ : LocalMux
    port map (
            O => \N__76336\,
            I => \N__76174\
        );

    \I__19076\ : LocalMux
    port map (
            O => \N__76331\,
            I => \N__76174\
        );

    \I__19075\ : LocalMux
    port map (
            O => \N__76326\,
            I => \N__76174\
        );

    \I__19074\ : LocalMux
    port map (
            O => \N__76323\,
            I => \N__76174\
        );

    \I__19073\ : InMux
    port map (
            O => \N__76322\,
            I => \N__76168\
        );

    \I__19072\ : InMux
    port map (
            O => \N__76321\,
            I => \N__76168\
        );

    \I__19071\ : Span4Mux_h
    port map (
            O => \N__76318\,
            I => \N__76159\
        );

    \I__19070\ : LocalMux
    port map (
            O => \N__76313\,
            I => \N__76159\
        );

    \I__19069\ : LocalMux
    port map (
            O => \N__76310\,
            I => \N__76159\
        );

    \I__19068\ : LocalMux
    port map (
            O => \N__76305\,
            I => \N__76159\
        );

    \I__19067\ : LocalMux
    port map (
            O => \N__76302\,
            I => \N__76152\
        );

    \I__19066\ : Span4Mux_v
    port map (
            O => \N__76299\,
            I => \N__76152\
        );

    \I__19065\ : LocalMux
    port map (
            O => \N__76294\,
            I => \N__76152\
        );

    \I__19064\ : InMux
    port map (
            O => \N__76293\,
            I => \N__76145\
        );

    \I__19063\ : InMux
    port map (
            O => \N__76292\,
            I => \N__76145\
        );

    \I__19062\ : InMux
    port map (
            O => \N__76291\,
            I => \N__76145\
        );

    \I__19061\ : InMux
    port map (
            O => \N__76288\,
            I => \N__76142\
        );

    \I__19060\ : InMux
    port map (
            O => \N__76287\,
            I => \N__76139\
        );

    \I__19059\ : InMux
    port map (
            O => \N__76286\,
            I => \N__76136\
        );

    \I__19058\ : LocalMux
    port map (
            O => \N__76277\,
            I => \N__76131\
        );

    \I__19057\ : Span4Mux_h
    port map (
            O => \N__76274\,
            I => \N__76131\
        );

    \I__19056\ : InMux
    port map (
            O => \N__76273\,
            I => \N__76128\
        );

    \I__19055\ : InMux
    port map (
            O => \N__76272\,
            I => \N__76123\
        );

    \I__19054\ : InMux
    port map (
            O => \N__76271\,
            I => \N__76123\
        );

    \I__19053\ : InMux
    port map (
            O => \N__76270\,
            I => \N__76118\
        );

    \I__19052\ : InMux
    port map (
            O => \N__76269\,
            I => \N__76118\
        );

    \I__19051\ : InMux
    port map (
            O => \N__76268\,
            I => \N__76113\
        );

    \I__19050\ : InMux
    port map (
            O => \N__76265\,
            I => \N__76113\
        );

    \I__19049\ : InMux
    port map (
            O => \N__76264\,
            I => \N__76110\
        );

    \I__19048\ : InMux
    port map (
            O => \N__76263\,
            I => \N__76103\
        );

    \I__19047\ : InMux
    port map (
            O => \N__76262\,
            I => \N__76103\
        );

    \I__19046\ : InMux
    port map (
            O => \N__76261\,
            I => \N__76103\
        );

    \I__19045\ : Span4Mux_v
    port map (
            O => \N__76258\,
            I => \N__76098\
        );

    \I__19044\ : LocalMux
    port map (
            O => \N__76251\,
            I => \N__76098\
        );

    \I__19043\ : Span4Mux_v
    port map (
            O => \N__76248\,
            I => \N__76089\
        );

    \I__19042\ : Span4Mux_h
    port map (
            O => \N__76241\,
            I => \N__76089\
        );

    \I__19041\ : Span4Mux_h
    port map (
            O => \N__76232\,
            I => \N__76089\
        );

    \I__19040\ : LocalMux
    port map (
            O => \N__76225\,
            I => \N__76089\
        );

    \I__19039\ : Span4Mux_v
    port map (
            O => \N__76222\,
            I => \N__76074\
        );

    \I__19038\ : Span4Mux_v
    port map (
            O => \N__76215\,
            I => \N__76074\
        );

    \I__19037\ : Span4Mux_v
    port map (
            O => \N__76210\,
            I => \N__76074\
        );

    \I__19036\ : LocalMux
    port map (
            O => \N__76203\,
            I => \N__76074\
        );

    \I__19035\ : Span4Mux_h
    port map (
            O => \N__76192\,
            I => \N__76074\
        );

    \I__19034\ : LocalMux
    port map (
            O => \N__76185\,
            I => \N__76074\
        );

    \I__19033\ : Span4Mux_v
    port map (
            O => \N__76174\,
            I => \N__76074\
        );

    \I__19032\ : InMux
    port map (
            O => \N__76173\,
            I => \N__76071\
        );

    \I__19031\ : LocalMux
    port map (
            O => \N__76168\,
            I => \N__76062\
        );

    \I__19030\ : Span4Mux_v
    port map (
            O => \N__76159\,
            I => \N__76062\
        );

    \I__19029\ : Span4Mux_h
    port map (
            O => \N__76152\,
            I => \N__76062\
        );

    \I__19028\ : LocalMux
    port map (
            O => \N__76145\,
            I => \N__76062\
        );

    \I__19027\ : LocalMux
    port map (
            O => \N__76142\,
            I => \N__76059\
        );

    \I__19026\ : LocalMux
    port map (
            O => \N__76139\,
            I => \progRomAddress_4\
        );

    \I__19025\ : LocalMux
    port map (
            O => \N__76136\,
            I => \progRomAddress_4\
        );

    \I__19024\ : Odrv4
    port map (
            O => \N__76131\,
            I => \progRomAddress_4\
        );

    \I__19023\ : LocalMux
    port map (
            O => \N__76128\,
            I => \progRomAddress_4\
        );

    \I__19022\ : LocalMux
    port map (
            O => \N__76123\,
            I => \progRomAddress_4\
        );

    \I__19021\ : LocalMux
    port map (
            O => \N__76118\,
            I => \progRomAddress_4\
        );

    \I__19020\ : LocalMux
    port map (
            O => \N__76113\,
            I => \progRomAddress_4\
        );

    \I__19019\ : LocalMux
    port map (
            O => \N__76110\,
            I => \progRomAddress_4\
        );

    \I__19018\ : LocalMux
    port map (
            O => \N__76103\,
            I => \progRomAddress_4\
        );

    \I__19017\ : Odrv4
    port map (
            O => \N__76098\,
            I => \progRomAddress_4\
        );

    \I__19016\ : Odrv4
    port map (
            O => \N__76089\,
            I => \progRomAddress_4\
        );

    \I__19015\ : Odrv4
    port map (
            O => \N__76074\,
            I => \progRomAddress_4\
        );

    \I__19014\ : LocalMux
    port map (
            O => \N__76071\,
            I => \progRomAddress_4\
        );

    \I__19013\ : Odrv4
    port map (
            O => \N__76062\,
            I => \progRomAddress_4\
        );

    \I__19012\ : Odrv12
    port map (
            O => \N__76059\,
            I => \progRomAddress_4\
        );

    \I__19011\ : CascadeMux
    port map (
            O => \N__76028\,
            I => \N__76025\
        );

    \I__19010\ : InMux
    port map (
            O => \N__76025\,
            I => \N__76022\
        );

    \I__19009\ : LocalMux
    port map (
            O => \N__76022\,
            I => \N__76019\
        );

    \I__19008\ : Odrv4
    port map (
            O => \N__76019\,
            I => \PROM.ROMDATA.m341_ns_1\
        );

    \I__19007\ : CascadeMux
    port map (
            O => \N__76016\,
            I => \N__76012\
        );

    \I__19006\ : InMux
    port map (
            O => \N__76015\,
            I => \N__76005\
        );

    \I__19005\ : InMux
    port map (
            O => \N__76012\,
            I => \N__75997\
        );

    \I__19004\ : InMux
    port map (
            O => \N__76011\,
            I => \N__75997\
        );

    \I__19003\ : CascadeMux
    port map (
            O => \N__76010\,
            I => \N__75987\
        );

    \I__19002\ : CascadeMux
    port map (
            O => \N__76009\,
            I => \N__75980\
        );

    \I__19001\ : CascadeMux
    port map (
            O => \N__76008\,
            I => \N__75977\
        );

    \I__19000\ : LocalMux
    port map (
            O => \N__76005\,
            I => \N__75974\
        );

    \I__18999\ : CascadeMux
    port map (
            O => \N__76004\,
            I => \N__75970\
        );

    \I__18998\ : CascadeMux
    port map (
            O => \N__76003\,
            I => \N__75956\
        );

    \I__18997\ : CascadeMux
    port map (
            O => \N__76002\,
            I => \N__75951\
        );

    \I__18996\ : LocalMux
    port map (
            O => \N__75997\,
            I => \N__75947\
        );

    \I__18995\ : InMux
    port map (
            O => \N__75996\,
            I => \N__75942\
        );

    \I__18994\ : InMux
    port map (
            O => \N__75995\,
            I => \N__75942\
        );

    \I__18993\ : CascadeMux
    port map (
            O => \N__75994\,
            I => \N__75935\
        );

    \I__18992\ : CascadeMux
    port map (
            O => \N__75993\,
            I => \N__75929\
        );

    \I__18991\ : CascadeMux
    port map (
            O => \N__75992\,
            I => \N__75926\
        );

    \I__18990\ : CascadeMux
    port map (
            O => \N__75991\,
            I => \N__75923\
        );

    \I__18989\ : CascadeMux
    port map (
            O => \N__75990\,
            I => \N__75920\
        );

    \I__18988\ : InMux
    port map (
            O => \N__75987\,
            I => \N__75896\
        );

    \I__18987\ : CascadeMux
    port map (
            O => \N__75986\,
            I => \N__75893\
        );

    \I__18986\ : InMux
    port map (
            O => \N__75985\,
            I => \N__75882\
        );

    \I__18985\ : CascadeMux
    port map (
            O => \N__75984\,
            I => \N__75876\
        );

    \I__18984\ : InMux
    port map (
            O => \N__75983\,
            I => \N__75871\
        );

    \I__18983\ : InMux
    port map (
            O => \N__75980\,
            I => \N__75871\
        );

    \I__18982\ : InMux
    port map (
            O => \N__75977\,
            I => \N__75868\
        );

    \I__18981\ : Span4Mux_v
    port map (
            O => \N__75974\,
            I => \N__75865\
        );

    \I__18980\ : InMux
    port map (
            O => \N__75973\,
            I => \N__75860\
        );

    \I__18979\ : InMux
    port map (
            O => \N__75970\,
            I => \N__75860\
        );

    \I__18978\ : InMux
    port map (
            O => \N__75969\,
            I => \N__75857\
        );

    \I__18977\ : CascadeMux
    port map (
            O => \N__75968\,
            I => \N__75853\
        );

    \I__18976\ : CascadeMux
    port map (
            O => \N__75967\,
            I => \N__75848\
        );

    \I__18975\ : CascadeMux
    port map (
            O => \N__75966\,
            I => \N__75843\
        );

    \I__18974\ : CascadeMux
    port map (
            O => \N__75965\,
            I => \N__75840\
        );

    \I__18973\ : CascadeMux
    port map (
            O => \N__75964\,
            I => \N__75836\
        );

    \I__18972\ : CascadeMux
    port map (
            O => \N__75963\,
            I => \N__75833\
        );

    \I__18971\ : CascadeMux
    port map (
            O => \N__75962\,
            I => \N__75825\
        );

    \I__18970\ : CascadeMux
    port map (
            O => \N__75961\,
            I => \N__75822\
        );

    \I__18969\ : CascadeMux
    port map (
            O => \N__75960\,
            I => \N__75818\
        );

    \I__18968\ : CascadeMux
    port map (
            O => \N__75959\,
            I => \N__75811\
        );

    \I__18967\ : InMux
    port map (
            O => \N__75956\,
            I => \N__75805\
        );

    \I__18966\ : CascadeMux
    port map (
            O => \N__75955\,
            I => \N__75801\
        );

    \I__18965\ : CascadeMux
    port map (
            O => \N__75954\,
            I => \N__75796\
        );

    \I__18964\ : InMux
    port map (
            O => \N__75951\,
            I => \N__75792\
        );

    \I__18963\ : CascadeMux
    port map (
            O => \N__75950\,
            I => \N__75786\
        );

    \I__18962\ : Span4Mux_h
    port map (
            O => \N__75947\,
            I => \N__75781\
        );

    \I__18961\ : LocalMux
    port map (
            O => \N__75942\,
            I => \N__75781\
        );

    \I__18960\ : InMux
    port map (
            O => \N__75941\,
            I => \N__75770\
        );

    \I__18959\ : InMux
    port map (
            O => \N__75940\,
            I => \N__75770\
        );

    \I__18958\ : InMux
    port map (
            O => \N__75939\,
            I => \N__75770\
        );

    \I__18957\ : InMux
    port map (
            O => \N__75938\,
            I => \N__75770\
        );

    \I__18956\ : InMux
    port map (
            O => \N__75935\,
            I => \N__75770\
        );

    \I__18955\ : InMux
    port map (
            O => \N__75934\,
            I => \N__75763\
        );

    \I__18954\ : InMux
    port map (
            O => \N__75933\,
            I => \N__75763\
        );

    \I__18953\ : InMux
    port map (
            O => \N__75932\,
            I => \N__75763\
        );

    \I__18952\ : InMux
    port map (
            O => \N__75929\,
            I => \N__75754\
        );

    \I__18951\ : InMux
    port map (
            O => \N__75926\,
            I => \N__75754\
        );

    \I__18950\ : InMux
    port map (
            O => \N__75923\,
            I => \N__75754\
        );

    \I__18949\ : InMux
    port map (
            O => \N__75920\,
            I => \N__75754\
        );

    \I__18948\ : CascadeMux
    port map (
            O => \N__75919\,
            I => \N__75751\
        );

    \I__18947\ : CascadeMux
    port map (
            O => \N__75918\,
            I => \N__75747\
        );

    \I__18946\ : CascadeMux
    port map (
            O => \N__75917\,
            I => \N__75743\
        );

    \I__18945\ : CascadeMux
    port map (
            O => \N__75916\,
            I => \N__75740\
        );

    \I__18944\ : CascadeMux
    port map (
            O => \N__75915\,
            I => \N__75737\
        );

    \I__18943\ : CascadeMux
    port map (
            O => \N__75914\,
            I => \N__75733\
        );

    \I__18942\ : CascadeMux
    port map (
            O => \N__75913\,
            I => \N__75730\
        );

    \I__18941\ : CascadeMux
    port map (
            O => \N__75912\,
            I => \N__75727\
        );

    \I__18940\ : CascadeMux
    port map (
            O => \N__75911\,
            I => \N__75722\
        );

    \I__18939\ : CascadeMux
    port map (
            O => \N__75910\,
            I => \N__75715\
        );

    \I__18938\ : CascadeMux
    port map (
            O => \N__75909\,
            I => \N__75712\
        );

    \I__18937\ : InMux
    port map (
            O => \N__75908\,
            I => \N__75705\
        );

    \I__18936\ : InMux
    port map (
            O => \N__75907\,
            I => \N__75702\
        );

    \I__18935\ : InMux
    port map (
            O => \N__75906\,
            I => \N__75695\
        );

    \I__18934\ : InMux
    port map (
            O => \N__75905\,
            I => \N__75695\
        );

    \I__18933\ : InMux
    port map (
            O => \N__75904\,
            I => \N__75695\
        );

    \I__18932\ : CascadeMux
    port map (
            O => \N__75903\,
            I => \N__75692\
        );

    \I__18931\ : CascadeMux
    port map (
            O => \N__75902\,
            I => \N__75689\
        );

    \I__18930\ : CascadeMux
    port map (
            O => \N__75901\,
            I => \N__75685\
        );

    \I__18929\ : CascadeMux
    port map (
            O => \N__75900\,
            I => \N__75681\
        );

    \I__18928\ : CascadeMux
    port map (
            O => \N__75899\,
            I => \N__75677\
        );

    \I__18927\ : LocalMux
    port map (
            O => \N__75896\,
            I => \N__75673\
        );

    \I__18926\ : InMux
    port map (
            O => \N__75893\,
            I => \N__75665\
        );

    \I__18925\ : InMux
    port map (
            O => \N__75892\,
            I => \N__75660\
        );

    \I__18924\ : InMux
    port map (
            O => \N__75891\,
            I => \N__75660\
        );

    \I__18923\ : CascadeMux
    port map (
            O => \N__75890\,
            I => \N__75656\
        );

    \I__18922\ : CascadeMux
    port map (
            O => \N__75889\,
            I => \N__75650\
        );

    \I__18921\ : CascadeMux
    port map (
            O => \N__75888\,
            I => \N__75647\
        );

    \I__18920\ : CascadeMux
    port map (
            O => \N__75887\,
            I => \N__75642\
        );

    \I__18919\ : CascadeMux
    port map (
            O => \N__75886\,
            I => \N__75639\
        );

    \I__18918\ : CascadeMux
    port map (
            O => \N__75885\,
            I => \N__75632\
        );

    \I__18917\ : LocalMux
    port map (
            O => \N__75882\,
            I => \N__75627\
        );

    \I__18916\ : InMux
    port map (
            O => \N__75881\,
            I => \N__75620\
        );

    \I__18915\ : InMux
    port map (
            O => \N__75880\,
            I => \N__75620\
        );

    \I__18914\ : InMux
    port map (
            O => \N__75879\,
            I => \N__75620\
        );

    \I__18913\ : InMux
    port map (
            O => \N__75876\,
            I => \N__75616\
        );

    \I__18912\ : LocalMux
    port map (
            O => \N__75871\,
            I => \N__75606\
        );

    \I__18911\ : LocalMux
    port map (
            O => \N__75868\,
            I => \N__75606\
        );

    \I__18910\ : Span4Mux_h
    port map (
            O => \N__75865\,
            I => \N__75599\
        );

    \I__18909\ : LocalMux
    port map (
            O => \N__75860\,
            I => \N__75599\
        );

    \I__18908\ : LocalMux
    port map (
            O => \N__75857\,
            I => \N__75599\
        );

    \I__18907\ : InMux
    port map (
            O => \N__75856\,
            I => \N__75594\
        );

    \I__18906\ : InMux
    port map (
            O => \N__75853\,
            I => \N__75587\
        );

    \I__18905\ : InMux
    port map (
            O => \N__75852\,
            I => \N__75587\
        );

    \I__18904\ : InMux
    port map (
            O => \N__75851\,
            I => \N__75587\
        );

    \I__18903\ : InMux
    port map (
            O => \N__75848\,
            I => \N__75580\
        );

    \I__18902\ : InMux
    port map (
            O => \N__75847\,
            I => \N__75580\
        );

    \I__18901\ : InMux
    port map (
            O => \N__75846\,
            I => \N__75580\
        );

    \I__18900\ : InMux
    port map (
            O => \N__75843\,
            I => \N__75577\
        );

    \I__18899\ : InMux
    port map (
            O => \N__75840\,
            I => \N__75570\
        );

    \I__18898\ : InMux
    port map (
            O => \N__75839\,
            I => \N__75570\
        );

    \I__18897\ : InMux
    port map (
            O => \N__75836\,
            I => \N__75570\
        );

    \I__18896\ : InMux
    port map (
            O => \N__75833\,
            I => \N__75561\
        );

    \I__18895\ : InMux
    port map (
            O => \N__75832\,
            I => \N__75561\
        );

    \I__18894\ : InMux
    port map (
            O => \N__75831\,
            I => \N__75561\
        );

    \I__18893\ : InMux
    port map (
            O => \N__75830\,
            I => \N__75561\
        );

    \I__18892\ : InMux
    port map (
            O => \N__75829\,
            I => \N__75556\
        );

    \I__18891\ : InMux
    port map (
            O => \N__75828\,
            I => \N__75556\
        );

    \I__18890\ : InMux
    port map (
            O => \N__75825\,
            I => \N__75551\
        );

    \I__18889\ : InMux
    port map (
            O => \N__75822\,
            I => \N__75551\
        );

    \I__18888\ : InMux
    port map (
            O => \N__75821\,
            I => \N__75546\
        );

    \I__18887\ : InMux
    port map (
            O => \N__75818\,
            I => \N__75546\
        );

    \I__18886\ : InMux
    port map (
            O => \N__75817\,
            I => \N__75541\
        );

    \I__18885\ : InMux
    port map (
            O => \N__75816\,
            I => \N__75541\
        );

    \I__18884\ : InMux
    port map (
            O => \N__75815\,
            I => \N__75535\
        );

    \I__18883\ : CascadeMux
    port map (
            O => \N__75814\,
            I => \N__75530\
        );

    \I__18882\ : InMux
    port map (
            O => \N__75811\,
            I => \N__75521\
        );

    \I__18881\ : InMux
    port map (
            O => \N__75810\,
            I => \N__75521\
        );

    \I__18880\ : InMux
    port map (
            O => \N__75809\,
            I => \N__75516\
        );

    \I__18879\ : InMux
    port map (
            O => \N__75808\,
            I => \N__75516\
        );

    \I__18878\ : LocalMux
    port map (
            O => \N__75805\,
            I => \N__75513\
        );

    \I__18877\ : InMux
    port map (
            O => \N__75804\,
            I => \N__75502\
        );

    \I__18876\ : InMux
    port map (
            O => \N__75801\,
            I => \N__75502\
        );

    \I__18875\ : InMux
    port map (
            O => \N__75800\,
            I => \N__75502\
        );

    \I__18874\ : InMux
    port map (
            O => \N__75799\,
            I => \N__75502\
        );

    \I__18873\ : InMux
    port map (
            O => \N__75796\,
            I => \N__75502\
        );

    \I__18872\ : CascadeMux
    port map (
            O => \N__75795\,
            I => \N__75496\
        );

    \I__18871\ : LocalMux
    port map (
            O => \N__75792\,
            I => \N__75493\
        );

    \I__18870\ : InMux
    port map (
            O => \N__75791\,
            I => \N__75490\
        );

    \I__18869\ : InMux
    port map (
            O => \N__75790\,
            I => \N__75483\
        );

    \I__18868\ : InMux
    port map (
            O => \N__75789\,
            I => \N__75483\
        );

    \I__18867\ : InMux
    port map (
            O => \N__75786\,
            I => \N__75483\
        );

    \I__18866\ : Span4Mux_h
    port map (
            O => \N__75781\,
            I => \N__75474\
        );

    \I__18865\ : LocalMux
    port map (
            O => \N__75770\,
            I => \N__75474\
        );

    \I__18864\ : LocalMux
    port map (
            O => \N__75763\,
            I => \N__75474\
        );

    \I__18863\ : LocalMux
    port map (
            O => \N__75754\,
            I => \N__75474\
        );

    \I__18862\ : InMux
    port map (
            O => \N__75751\,
            I => \N__75467\
        );

    \I__18861\ : InMux
    port map (
            O => \N__75750\,
            I => \N__75467\
        );

    \I__18860\ : InMux
    port map (
            O => \N__75747\,
            I => \N__75467\
        );

    \I__18859\ : InMux
    port map (
            O => \N__75746\,
            I => \N__75460\
        );

    \I__18858\ : InMux
    port map (
            O => \N__75743\,
            I => \N__75460\
        );

    \I__18857\ : InMux
    port map (
            O => \N__75740\,
            I => \N__75460\
        );

    \I__18856\ : InMux
    port map (
            O => \N__75737\,
            I => \N__75453\
        );

    \I__18855\ : InMux
    port map (
            O => \N__75736\,
            I => \N__75453\
        );

    \I__18854\ : InMux
    port map (
            O => \N__75733\,
            I => \N__75453\
        );

    \I__18853\ : InMux
    port map (
            O => \N__75730\,
            I => \N__75446\
        );

    \I__18852\ : InMux
    port map (
            O => \N__75727\,
            I => \N__75446\
        );

    \I__18851\ : InMux
    port map (
            O => \N__75726\,
            I => \N__75446\
        );

    \I__18850\ : InMux
    port map (
            O => \N__75725\,
            I => \N__75439\
        );

    \I__18849\ : InMux
    port map (
            O => \N__75722\,
            I => \N__75439\
        );

    \I__18848\ : InMux
    port map (
            O => \N__75721\,
            I => \N__75439\
        );

    \I__18847\ : InMux
    port map (
            O => \N__75720\,
            I => \N__75430\
        );

    \I__18846\ : InMux
    port map (
            O => \N__75719\,
            I => \N__75430\
        );

    \I__18845\ : InMux
    port map (
            O => \N__75718\,
            I => \N__75430\
        );

    \I__18844\ : InMux
    port map (
            O => \N__75715\,
            I => \N__75430\
        );

    \I__18843\ : InMux
    port map (
            O => \N__75712\,
            I => \N__75425\
        );

    \I__18842\ : InMux
    port map (
            O => \N__75711\,
            I => \N__75425\
        );

    \I__18841\ : CascadeMux
    port map (
            O => \N__75710\,
            I => \N__75419\
        );

    \I__18840\ : CascadeMux
    port map (
            O => \N__75709\,
            I => \N__75416\
        );

    \I__18839\ : InMux
    port map (
            O => \N__75708\,
            I => \N__75413\
        );

    \I__18838\ : LocalMux
    port map (
            O => \N__75705\,
            I => \N__75410\
        );

    \I__18837\ : LocalMux
    port map (
            O => \N__75702\,
            I => \N__75407\
        );

    \I__18836\ : LocalMux
    port map (
            O => \N__75695\,
            I => \N__75404\
        );

    \I__18835\ : InMux
    port map (
            O => \N__75692\,
            I => \N__75401\
        );

    \I__18834\ : InMux
    port map (
            O => \N__75689\,
            I => \N__75394\
        );

    \I__18833\ : InMux
    port map (
            O => \N__75688\,
            I => \N__75394\
        );

    \I__18832\ : InMux
    port map (
            O => \N__75685\,
            I => \N__75394\
        );

    \I__18831\ : InMux
    port map (
            O => \N__75684\,
            I => \N__75385\
        );

    \I__18830\ : InMux
    port map (
            O => \N__75681\,
            I => \N__75385\
        );

    \I__18829\ : InMux
    port map (
            O => \N__75680\,
            I => \N__75385\
        );

    \I__18828\ : InMux
    port map (
            O => \N__75677\,
            I => \N__75385\
        );

    \I__18827\ : CascadeMux
    port map (
            O => \N__75676\,
            I => \N__75380\
        );

    \I__18826\ : Span4Mux_h
    port map (
            O => \N__75673\,
            I => \N__75377\
        );

    \I__18825\ : InMux
    port map (
            O => \N__75672\,
            I => \N__75366\
        );

    \I__18824\ : InMux
    port map (
            O => \N__75671\,
            I => \N__75366\
        );

    \I__18823\ : InMux
    port map (
            O => \N__75670\,
            I => \N__75366\
        );

    \I__18822\ : InMux
    port map (
            O => \N__75669\,
            I => \N__75366\
        );

    \I__18821\ : InMux
    port map (
            O => \N__75668\,
            I => \N__75366\
        );

    \I__18820\ : LocalMux
    port map (
            O => \N__75665\,
            I => \N__75361\
        );

    \I__18819\ : LocalMux
    port map (
            O => \N__75660\,
            I => \N__75361\
        );

    \I__18818\ : InMux
    port map (
            O => \N__75659\,
            I => \N__75348\
        );

    \I__18817\ : InMux
    port map (
            O => \N__75656\,
            I => \N__75348\
        );

    \I__18816\ : InMux
    port map (
            O => \N__75655\,
            I => \N__75348\
        );

    \I__18815\ : InMux
    port map (
            O => \N__75654\,
            I => \N__75348\
        );

    \I__18814\ : InMux
    port map (
            O => \N__75653\,
            I => \N__75348\
        );

    \I__18813\ : InMux
    port map (
            O => \N__75650\,
            I => \N__75348\
        );

    \I__18812\ : InMux
    port map (
            O => \N__75647\,
            I => \N__75339\
        );

    \I__18811\ : InMux
    port map (
            O => \N__75646\,
            I => \N__75339\
        );

    \I__18810\ : InMux
    port map (
            O => \N__75645\,
            I => \N__75339\
        );

    \I__18809\ : InMux
    port map (
            O => \N__75642\,
            I => \N__75339\
        );

    \I__18808\ : InMux
    port map (
            O => \N__75639\,
            I => \N__75336\
        );

    \I__18807\ : InMux
    port map (
            O => \N__75638\,
            I => \N__75329\
        );

    \I__18806\ : InMux
    port map (
            O => \N__75637\,
            I => \N__75329\
        );

    \I__18805\ : InMux
    port map (
            O => \N__75636\,
            I => \N__75329\
        );

    \I__18804\ : InMux
    port map (
            O => \N__75635\,
            I => \N__75320\
        );

    \I__18803\ : InMux
    port map (
            O => \N__75632\,
            I => \N__75320\
        );

    \I__18802\ : InMux
    port map (
            O => \N__75631\,
            I => \N__75320\
        );

    \I__18801\ : InMux
    port map (
            O => \N__75630\,
            I => \N__75320\
        );

    \I__18800\ : Span4Mux_v
    port map (
            O => \N__75627\,
            I => \N__75317\
        );

    \I__18799\ : LocalMux
    port map (
            O => \N__75620\,
            I => \N__75314\
        );

    \I__18798\ : InMux
    port map (
            O => \N__75619\,
            I => \N__75311\
        );

    \I__18797\ : LocalMux
    port map (
            O => \N__75616\,
            I => \N__75308\
        );

    \I__18796\ : CascadeMux
    port map (
            O => \N__75615\,
            I => \N__75300\
        );

    \I__18795\ : CascadeMux
    port map (
            O => \N__75614\,
            I => \N__75296\
        );

    \I__18794\ : CascadeMux
    port map (
            O => \N__75613\,
            I => \N__75293\
        );

    \I__18793\ : CascadeMux
    port map (
            O => \N__75612\,
            I => \N__75288\
        );

    \I__18792\ : CascadeMux
    port map (
            O => \N__75611\,
            I => \N__75284\
        );

    \I__18791\ : Span4Mux_v
    port map (
            O => \N__75606\,
            I => \N__75280\
        );

    \I__18790\ : Span4Mux_v
    port map (
            O => \N__75599\,
            I => \N__75277\
        );

    \I__18789\ : InMux
    port map (
            O => \N__75598\,
            I => \N__75272\
        );

    \I__18788\ : InMux
    port map (
            O => \N__75597\,
            I => \N__75272\
        );

    \I__18787\ : LocalMux
    port map (
            O => \N__75594\,
            I => \N__75263\
        );

    \I__18786\ : LocalMux
    port map (
            O => \N__75587\,
            I => \N__75263\
        );

    \I__18785\ : LocalMux
    port map (
            O => \N__75580\,
            I => \N__75263\
        );

    \I__18784\ : LocalMux
    port map (
            O => \N__75577\,
            I => \N__75263\
        );

    \I__18783\ : LocalMux
    port map (
            O => \N__75570\,
            I => \N__75258\
        );

    \I__18782\ : LocalMux
    port map (
            O => \N__75561\,
            I => \N__75258\
        );

    \I__18781\ : LocalMux
    port map (
            O => \N__75556\,
            I => \N__75249\
        );

    \I__18780\ : LocalMux
    port map (
            O => \N__75551\,
            I => \N__75249\
        );

    \I__18779\ : LocalMux
    port map (
            O => \N__75546\,
            I => \N__75249\
        );

    \I__18778\ : LocalMux
    port map (
            O => \N__75541\,
            I => \N__75249\
        );

    \I__18777\ : CascadeMux
    port map (
            O => \N__75540\,
            I => \N__75244\
        );

    \I__18776\ : CascadeMux
    port map (
            O => \N__75539\,
            I => \N__75240\
        );

    \I__18775\ : CascadeMux
    port map (
            O => \N__75538\,
            I => \N__75237\
        );

    \I__18774\ : LocalMux
    port map (
            O => \N__75535\,
            I => \N__75231\
        );

    \I__18773\ : InMux
    port map (
            O => \N__75534\,
            I => \N__75224\
        );

    \I__18772\ : InMux
    port map (
            O => \N__75533\,
            I => \N__75224\
        );

    \I__18771\ : InMux
    port map (
            O => \N__75530\,
            I => \N__75224\
        );

    \I__18770\ : InMux
    port map (
            O => \N__75529\,
            I => \N__75215\
        );

    \I__18769\ : InMux
    port map (
            O => \N__75528\,
            I => \N__75215\
        );

    \I__18768\ : InMux
    port map (
            O => \N__75527\,
            I => \N__75215\
        );

    \I__18767\ : InMux
    port map (
            O => \N__75526\,
            I => \N__75215\
        );

    \I__18766\ : LocalMux
    port map (
            O => \N__75521\,
            I => \N__75212\
        );

    \I__18765\ : LocalMux
    port map (
            O => \N__75516\,
            I => \N__75205\
        );

    \I__18764\ : Span4Mux_v
    port map (
            O => \N__75513\,
            I => \N__75205\
        );

    \I__18763\ : LocalMux
    port map (
            O => \N__75502\,
            I => \N__75205\
        );

    \I__18762\ : InMux
    port map (
            O => \N__75501\,
            I => \N__75196\
        );

    \I__18761\ : InMux
    port map (
            O => \N__75500\,
            I => \N__75196\
        );

    \I__18760\ : InMux
    port map (
            O => \N__75499\,
            I => \N__75196\
        );

    \I__18759\ : InMux
    port map (
            O => \N__75496\,
            I => \N__75196\
        );

    \I__18758\ : Span4Mux_h
    port map (
            O => \N__75493\,
            I => \N__75179\
        );

    \I__18757\ : LocalMux
    port map (
            O => \N__75490\,
            I => \N__75179\
        );

    \I__18756\ : LocalMux
    port map (
            O => \N__75483\,
            I => \N__75179\
        );

    \I__18755\ : Span4Mux_v
    port map (
            O => \N__75474\,
            I => \N__75179\
        );

    \I__18754\ : LocalMux
    port map (
            O => \N__75467\,
            I => \N__75179\
        );

    \I__18753\ : LocalMux
    port map (
            O => \N__75460\,
            I => \N__75179\
        );

    \I__18752\ : LocalMux
    port map (
            O => \N__75453\,
            I => \N__75179\
        );

    \I__18751\ : LocalMux
    port map (
            O => \N__75446\,
            I => \N__75179\
        );

    \I__18750\ : LocalMux
    port map (
            O => \N__75439\,
            I => \N__75172\
        );

    \I__18749\ : LocalMux
    port map (
            O => \N__75430\,
            I => \N__75172\
        );

    \I__18748\ : LocalMux
    port map (
            O => \N__75425\,
            I => \N__75172\
        );

    \I__18747\ : InMux
    port map (
            O => \N__75424\,
            I => \N__75161\
        );

    \I__18746\ : InMux
    port map (
            O => \N__75423\,
            I => \N__75161\
        );

    \I__18745\ : InMux
    port map (
            O => \N__75422\,
            I => \N__75161\
        );

    \I__18744\ : InMux
    port map (
            O => \N__75419\,
            I => \N__75161\
        );

    \I__18743\ : InMux
    port map (
            O => \N__75416\,
            I => \N__75161\
        );

    \I__18742\ : LocalMux
    port map (
            O => \N__75413\,
            I => \N__75158\
        );

    \I__18741\ : Span4Mux_h
    port map (
            O => \N__75410\,
            I => \N__75151\
        );

    \I__18740\ : Span4Mux_v
    port map (
            O => \N__75407\,
            I => \N__75151\
        );

    \I__18739\ : Span4Mux_h
    port map (
            O => \N__75404\,
            I => \N__75151\
        );

    \I__18738\ : LocalMux
    port map (
            O => \N__75401\,
            I => \N__75144\
        );

    \I__18737\ : LocalMux
    port map (
            O => \N__75394\,
            I => \N__75144\
        );

    \I__18736\ : LocalMux
    port map (
            O => \N__75385\,
            I => \N__75144\
        );

    \I__18735\ : InMux
    port map (
            O => \N__75384\,
            I => \N__75137\
        );

    \I__18734\ : InMux
    port map (
            O => \N__75383\,
            I => \N__75137\
        );

    \I__18733\ : InMux
    port map (
            O => \N__75380\,
            I => \N__75137\
        );

    \I__18732\ : Span4Mux_v
    port map (
            O => \N__75377\,
            I => \N__75126\
        );

    \I__18731\ : LocalMux
    port map (
            O => \N__75366\,
            I => \N__75126\
        );

    \I__18730\ : Span4Mux_h
    port map (
            O => \N__75361\,
            I => \N__75126\
        );

    \I__18729\ : LocalMux
    port map (
            O => \N__75348\,
            I => \N__75126\
        );

    \I__18728\ : LocalMux
    port map (
            O => \N__75339\,
            I => \N__75126\
        );

    \I__18727\ : LocalMux
    port map (
            O => \N__75336\,
            I => \N__75123\
        );

    \I__18726\ : LocalMux
    port map (
            O => \N__75329\,
            I => \N__75118\
        );

    \I__18725\ : LocalMux
    port map (
            O => \N__75320\,
            I => \N__75118\
        );

    \I__18724\ : Span4Mux_h
    port map (
            O => \N__75317\,
            I => \N__75109\
        );

    \I__18723\ : Span4Mux_v
    port map (
            O => \N__75314\,
            I => \N__75109\
        );

    \I__18722\ : LocalMux
    port map (
            O => \N__75311\,
            I => \N__75109\
        );

    \I__18721\ : Span4Mux_v
    port map (
            O => \N__75308\,
            I => \N__75109\
        );

    \I__18720\ : InMux
    port map (
            O => \N__75307\,
            I => \N__75106\
        );

    \I__18719\ : InMux
    port map (
            O => \N__75306\,
            I => \N__75101\
        );

    \I__18718\ : InMux
    port map (
            O => \N__75305\,
            I => \N__75101\
        );

    \I__18717\ : InMux
    port map (
            O => \N__75304\,
            I => \N__75090\
        );

    \I__18716\ : InMux
    port map (
            O => \N__75303\,
            I => \N__75090\
        );

    \I__18715\ : InMux
    port map (
            O => \N__75300\,
            I => \N__75090\
        );

    \I__18714\ : InMux
    port map (
            O => \N__75299\,
            I => \N__75090\
        );

    \I__18713\ : InMux
    port map (
            O => \N__75296\,
            I => \N__75090\
        );

    \I__18712\ : InMux
    port map (
            O => \N__75293\,
            I => \N__75083\
        );

    \I__18711\ : InMux
    port map (
            O => \N__75292\,
            I => \N__75083\
        );

    \I__18710\ : InMux
    port map (
            O => \N__75291\,
            I => \N__75083\
        );

    \I__18709\ : InMux
    port map (
            O => \N__75288\,
            I => \N__75074\
        );

    \I__18708\ : InMux
    port map (
            O => \N__75287\,
            I => \N__75074\
        );

    \I__18707\ : InMux
    port map (
            O => \N__75284\,
            I => \N__75074\
        );

    \I__18706\ : InMux
    port map (
            O => \N__75283\,
            I => \N__75074\
        );

    \I__18705\ : Span4Mux_h
    port map (
            O => \N__75280\,
            I => \N__75061\
        );

    \I__18704\ : Span4Mux_h
    port map (
            O => \N__75277\,
            I => \N__75061\
        );

    \I__18703\ : LocalMux
    port map (
            O => \N__75272\,
            I => \N__75061\
        );

    \I__18702\ : Span4Mux_v
    port map (
            O => \N__75263\,
            I => \N__75061\
        );

    \I__18701\ : Span4Mux_v
    port map (
            O => \N__75258\,
            I => \N__75061\
        );

    \I__18700\ : Span4Mux_v
    port map (
            O => \N__75249\,
            I => \N__75061\
        );

    \I__18699\ : InMux
    port map (
            O => \N__75248\,
            I => \N__75050\
        );

    \I__18698\ : InMux
    port map (
            O => \N__75247\,
            I => \N__75050\
        );

    \I__18697\ : InMux
    port map (
            O => \N__75244\,
            I => \N__75050\
        );

    \I__18696\ : InMux
    port map (
            O => \N__75243\,
            I => \N__75050\
        );

    \I__18695\ : InMux
    port map (
            O => \N__75240\,
            I => \N__75050\
        );

    \I__18694\ : InMux
    port map (
            O => \N__75237\,
            I => \N__75041\
        );

    \I__18693\ : InMux
    port map (
            O => \N__75236\,
            I => \N__75041\
        );

    \I__18692\ : InMux
    port map (
            O => \N__75235\,
            I => \N__75041\
        );

    \I__18691\ : InMux
    port map (
            O => \N__75234\,
            I => \N__75041\
        );

    \I__18690\ : Span4Mux_h
    port map (
            O => \N__75231\,
            I => \N__75034\
        );

    \I__18689\ : LocalMux
    port map (
            O => \N__75224\,
            I => \N__75034\
        );

    \I__18688\ : LocalMux
    port map (
            O => \N__75215\,
            I => \N__75034\
        );

    \I__18687\ : Span4Mux_h
    port map (
            O => \N__75212\,
            I => \N__75021\
        );

    \I__18686\ : Span4Mux_v
    port map (
            O => \N__75205\,
            I => \N__75021\
        );

    \I__18685\ : LocalMux
    port map (
            O => \N__75196\,
            I => \N__75021\
        );

    \I__18684\ : Span4Mux_v
    port map (
            O => \N__75179\,
            I => \N__75021\
        );

    \I__18683\ : Span4Mux_v
    port map (
            O => \N__75172\,
            I => \N__75021\
        );

    \I__18682\ : LocalMux
    port map (
            O => \N__75161\,
            I => \N__75021\
        );

    \I__18681\ : Span4Mux_h
    port map (
            O => \N__75158\,
            I => \N__75010\
        );

    \I__18680\ : Span4Mux_h
    port map (
            O => \N__75151\,
            I => \N__75010\
        );

    \I__18679\ : Span4Mux_h
    port map (
            O => \N__75144\,
            I => \N__75010\
        );

    \I__18678\ : LocalMux
    port map (
            O => \N__75137\,
            I => \N__75010\
        );

    \I__18677\ : Span4Mux_h
    port map (
            O => \N__75126\,
            I => \N__75010\
        );

    \I__18676\ : Span4Mux_h
    port map (
            O => \N__75123\,
            I => \N__75003\
        );

    \I__18675\ : Span4Mux_h
    port map (
            O => \N__75118\,
            I => \N__75003\
        );

    \I__18674\ : Span4Mux_h
    port map (
            O => \N__75109\,
            I => \N__75003\
        );

    \I__18673\ : LocalMux
    port map (
            O => \N__75106\,
            I => \progRomAddress_3\
        );

    \I__18672\ : LocalMux
    port map (
            O => \N__75101\,
            I => \progRomAddress_3\
        );

    \I__18671\ : LocalMux
    port map (
            O => \N__75090\,
            I => \progRomAddress_3\
        );

    \I__18670\ : LocalMux
    port map (
            O => \N__75083\,
            I => \progRomAddress_3\
        );

    \I__18669\ : LocalMux
    port map (
            O => \N__75074\,
            I => \progRomAddress_3\
        );

    \I__18668\ : Odrv4
    port map (
            O => \N__75061\,
            I => \progRomAddress_3\
        );

    \I__18667\ : LocalMux
    port map (
            O => \N__75050\,
            I => \progRomAddress_3\
        );

    \I__18666\ : LocalMux
    port map (
            O => \N__75041\,
            I => \progRomAddress_3\
        );

    \I__18665\ : Odrv4
    port map (
            O => \N__75034\,
            I => \progRomAddress_3\
        );

    \I__18664\ : Odrv4
    port map (
            O => \N__75021\,
            I => \progRomAddress_3\
        );

    \I__18663\ : Odrv4
    port map (
            O => \N__75010\,
            I => \progRomAddress_3\
        );

    \I__18662\ : Odrv4
    port map (
            O => \N__75003\,
            I => \progRomAddress_3\
        );

    \I__18661\ : InMux
    port map (
            O => \N__74978\,
            I => \N__74975\
        );

    \I__18660\ : LocalMux
    port map (
            O => \N__74975\,
            I => \PROM.ROMDATA.m341_ns\
        );

    \I__18659\ : InMux
    port map (
            O => \N__74972\,
            I => \N__74969\
        );

    \I__18658\ : LocalMux
    port map (
            O => \N__74969\,
            I => \N__74966\
        );

    \I__18657\ : Odrv4
    port map (
            O => \N__74966\,
            I => \PROM.ROMDATA.m347\
        );

    \I__18656\ : InMux
    port map (
            O => \N__74963\,
            I => \N__74959\
        );

    \I__18655\ : InMux
    port map (
            O => \N__74962\,
            I => \N__74956\
        );

    \I__18654\ : LocalMux
    port map (
            O => \N__74959\,
            I => \N__74953\
        );

    \I__18653\ : LocalMux
    port map (
            O => \N__74956\,
            I => \N__74950\
        );

    \I__18652\ : Odrv4
    port map (
            O => \N__74953\,
            I => \PROM.ROMDATA.m112\
        );

    \I__18651\ : Odrv4
    port map (
            O => \N__74950\,
            I => \PROM.ROMDATA.m112\
        );

    \I__18650\ : InMux
    port map (
            O => \N__74945\,
            I => \N__74942\
        );

    \I__18649\ : LocalMux
    port map (
            O => \N__74942\,
            I => \PROM.ROMDATA.m349_am\
        );

    \I__18648\ : CascadeMux
    port map (
            O => \N__74939\,
            I => \PROM.ROMDATA.m349_bm_cascade_\
        );

    \I__18647\ : InMux
    port map (
            O => \N__74936\,
            I => \N__74933\
        );

    \I__18646\ : LocalMux
    port map (
            O => \N__74933\,
            I => \PROM.ROMDATA.m349_ns\
        );

    \I__18645\ : CascadeMux
    port map (
            O => \N__74930\,
            I => \PROM.ROMDATA.m331_bm_cascade_\
        );

    \I__18644\ : InMux
    port map (
            O => \N__74927\,
            I => \N__74924\
        );

    \I__18643\ : LocalMux
    port map (
            O => \N__74924\,
            I => \N__74921\
        );

    \I__18642\ : Span4Mux_v
    port map (
            O => \N__74921\,
            I => \N__74918\
        );

    \I__18641\ : Odrv4
    port map (
            O => \N__74918\,
            I => \PROM.ROMDATA.m323_bm\
        );

    \I__18640\ : CascadeMux
    port map (
            O => \N__74915\,
            I => \PROM.ROMDATA.m323_am_cascade_\
        );

    \I__18639\ : InMux
    port map (
            O => \N__74912\,
            I => \N__74909\
        );

    \I__18638\ : LocalMux
    port map (
            O => \N__74909\,
            I => \N__74906\
        );

    \I__18637\ : Odrv12
    port map (
            O => \N__74906\,
            I => \PROM.ROMDATA.m323_ns\
        );

    \I__18636\ : CascadeMux
    port map (
            O => \N__74903\,
            I => \N__74899\
        );

    \I__18635\ : CascadeMux
    port map (
            O => \N__74902\,
            I => \N__74896\
        );

    \I__18634\ : InMux
    port map (
            O => \N__74899\,
            I => \N__74891\
        );

    \I__18633\ : InMux
    port map (
            O => \N__74896\,
            I => \N__74883\
        );

    \I__18632\ : InMux
    port map (
            O => \N__74895\,
            I => \N__74879\
        );

    \I__18631\ : CascadeMux
    port map (
            O => \N__74894\,
            I => \N__74876\
        );

    \I__18630\ : LocalMux
    port map (
            O => \N__74891\,
            I => \N__74873\
        );

    \I__18629\ : InMux
    port map (
            O => \N__74890\,
            I => \N__74870\
        );

    \I__18628\ : CascadeMux
    port map (
            O => \N__74889\,
            I => \N__74867\
        );

    \I__18627\ : CascadeMux
    port map (
            O => \N__74888\,
            I => \N__74864\
        );

    \I__18626\ : CascadeMux
    port map (
            O => \N__74887\,
            I => \N__74861\
        );

    \I__18625\ : CascadeMux
    port map (
            O => \N__74886\,
            I => \N__74857\
        );

    \I__18624\ : LocalMux
    port map (
            O => \N__74883\,
            I => \N__74850\
        );

    \I__18623\ : InMux
    port map (
            O => \N__74882\,
            I => \N__74847\
        );

    \I__18622\ : LocalMux
    port map (
            O => \N__74879\,
            I => \N__74844\
        );

    \I__18621\ : InMux
    port map (
            O => \N__74876\,
            I => \N__74841\
        );

    \I__18620\ : Span4Mux_v
    port map (
            O => \N__74873\,
            I => \N__74838\
        );

    \I__18619\ : LocalMux
    port map (
            O => \N__74870\,
            I => \N__74835\
        );

    \I__18618\ : InMux
    port map (
            O => \N__74867\,
            I => \N__74827\
        );

    \I__18617\ : InMux
    port map (
            O => \N__74864\,
            I => \N__74827\
        );

    \I__18616\ : InMux
    port map (
            O => \N__74861\,
            I => \N__74817\
        );

    \I__18615\ : InMux
    port map (
            O => \N__74860\,
            I => \N__74817\
        );

    \I__18614\ : InMux
    port map (
            O => \N__74857\,
            I => \N__74817\
        );

    \I__18613\ : InMux
    port map (
            O => \N__74856\,
            I => \N__74812\
        );

    \I__18612\ : InMux
    port map (
            O => \N__74855\,
            I => \N__74809\
        );

    \I__18611\ : InMux
    port map (
            O => \N__74854\,
            I => \N__74804\
        );

    \I__18610\ : InMux
    port map (
            O => \N__74853\,
            I => \N__74804\
        );

    \I__18609\ : Span4Mux_v
    port map (
            O => \N__74850\,
            I => \N__74801\
        );

    \I__18608\ : LocalMux
    port map (
            O => \N__74847\,
            I => \N__74798\
        );

    \I__18607\ : Span4Mux_h
    port map (
            O => \N__74844\,
            I => \N__74793\
        );

    \I__18606\ : LocalMux
    port map (
            O => \N__74841\,
            I => \N__74793\
        );

    \I__18605\ : Span4Mux_h
    port map (
            O => \N__74838\,
            I => \N__74788\
        );

    \I__18604\ : Span4Mux_h
    port map (
            O => \N__74835\,
            I => \N__74788\
        );

    \I__18603\ : InMux
    port map (
            O => \N__74834\,
            I => \N__74785\
        );

    \I__18602\ : InMux
    port map (
            O => \N__74833\,
            I => \N__74782\
        );

    \I__18601\ : CascadeMux
    port map (
            O => \N__74832\,
            I => \N__74779\
        );

    \I__18600\ : LocalMux
    port map (
            O => \N__74827\,
            I => \N__74775\
        );

    \I__18599\ : CascadeMux
    port map (
            O => \N__74826\,
            I => \N__74772\
        );

    \I__18598\ : CascadeMux
    port map (
            O => \N__74825\,
            I => \N__74768\
        );

    \I__18597\ : CascadeMux
    port map (
            O => \N__74824\,
            I => \N__74765\
        );

    \I__18596\ : LocalMux
    port map (
            O => \N__74817\,
            I => \N__74762\
        );

    \I__18595\ : CascadeMux
    port map (
            O => \N__74816\,
            I => \N__74759\
        );

    \I__18594\ : InMux
    port map (
            O => \N__74815\,
            I => \N__74756\
        );

    \I__18593\ : LocalMux
    port map (
            O => \N__74812\,
            I => \N__74753\
        );

    \I__18592\ : LocalMux
    port map (
            O => \N__74809\,
            I => \N__74750\
        );

    \I__18591\ : LocalMux
    port map (
            O => \N__74804\,
            I => \N__74739\
        );

    \I__18590\ : Span4Mux_h
    port map (
            O => \N__74801\,
            I => \N__74739\
        );

    \I__18589\ : Span4Mux_v
    port map (
            O => \N__74798\,
            I => \N__74739\
        );

    \I__18588\ : Span4Mux_v
    port map (
            O => \N__74793\,
            I => \N__74739\
        );

    \I__18587\ : Span4Mux_h
    port map (
            O => \N__74788\,
            I => \N__74739\
        );

    \I__18586\ : LocalMux
    port map (
            O => \N__74785\,
            I => \N__74736\
        );

    \I__18585\ : LocalMux
    port map (
            O => \N__74782\,
            I => \N__74733\
        );

    \I__18584\ : InMux
    port map (
            O => \N__74779\,
            I => \N__74730\
        );

    \I__18583\ : InMux
    port map (
            O => \N__74778\,
            I => \N__74727\
        );

    \I__18582\ : Span4Mux_v
    port map (
            O => \N__74775\,
            I => \N__74724\
        );

    \I__18581\ : InMux
    port map (
            O => \N__74772\,
            I => \N__74715\
        );

    \I__18580\ : InMux
    port map (
            O => \N__74771\,
            I => \N__74715\
        );

    \I__18579\ : InMux
    port map (
            O => \N__74768\,
            I => \N__74715\
        );

    \I__18578\ : InMux
    port map (
            O => \N__74765\,
            I => \N__74715\
        );

    \I__18577\ : Span4Mux_v
    port map (
            O => \N__74762\,
            I => \N__74712\
        );

    \I__18576\ : InMux
    port map (
            O => \N__74759\,
            I => \N__74709\
        );

    \I__18575\ : LocalMux
    port map (
            O => \N__74756\,
            I => \N__74706\
        );

    \I__18574\ : Span4Mux_h
    port map (
            O => \N__74753\,
            I => \N__74703\
        );

    \I__18573\ : Span4Mux_v
    port map (
            O => \N__74750\,
            I => \N__74700\
        );

    \I__18572\ : Span4Mux_h
    port map (
            O => \N__74739\,
            I => \N__74697\
        );

    \I__18571\ : Span4Mux_v
    port map (
            O => \N__74736\,
            I => \N__74694\
        );

    \I__18570\ : Span4Mux_v
    port map (
            O => \N__74733\,
            I => \N__74691\
        );

    \I__18569\ : LocalMux
    port map (
            O => \N__74730\,
            I => \N__74686\
        );

    \I__18568\ : LocalMux
    port map (
            O => \N__74727\,
            I => \N__74686\
        );

    \I__18567\ : Span4Mux_v
    port map (
            O => \N__74724\,
            I => \N__74683\
        );

    \I__18566\ : LocalMux
    port map (
            O => \N__74715\,
            I => \N__74674\
        );

    \I__18565\ : Sp12to4
    port map (
            O => \N__74712\,
            I => \N__74674\
        );

    \I__18564\ : LocalMux
    port map (
            O => \N__74709\,
            I => \N__74674\
        );

    \I__18563\ : Span4Mux_h
    port map (
            O => \N__74706\,
            I => \N__74671\
        );

    \I__18562\ : Span4Mux_v
    port map (
            O => \N__74703\,
            I => \N__74666\
        );

    \I__18561\ : Span4Mux_h
    port map (
            O => \N__74700\,
            I => \N__74666\
        );

    \I__18560\ : Span4Mux_v
    port map (
            O => \N__74697\,
            I => \N__74663\
        );

    \I__18559\ : Span4Mux_v
    port map (
            O => \N__74694\,
            I => \N__74658\
        );

    \I__18558\ : Span4Mux_h
    port map (
            O => \N__74691\,
            I => \N__74658\
        );

    \I__18557\ : Span4Mux_h
    port map (
            O => \N__74686\,
            I => \N__74655\
        );

    \I__18556\ : Span4Mux_h
    port map (
            O => \N__74683\,
            I => \N__74652\
        );

    \I__18555\ : InMux
    port map (
            O => \N__74682\,
            I => \N__74649\
        );

    \I__18554\ : InMux
    port map (
            O => \N__74681\,
            I => \N__74646\
        );

    \I__18553\ : Span12Mux_h
    port map (
            O => \N__74674\,
            I => \N__74643\
        );

    \I__18552\ : Span4Mux_h
    port map (
            O => \N__74671\,
            I => \N__74636\
        );

    \I__18551\ : Span4Mux_h
    port map (
            O => \N__74666\,
            I => \N__74636\
        );

    \I__18550\ : Span4Mux_v
    port map (
            O => \N__74663\,
            I => \N__74636\
        );

    \I__18549\ : Span4Mux_h
    port map (
            O => \N__74658\,
            I => \N__74629\
        );

    \I__18548\ : Span4Mux_v
    port map (
            O => \N__74655\,
            I => \N__74629\
        );

    \I__18547\ : Span4Mux_h
    port map (
            O => \N__74652\,
            I => \N__74629\
        );

    \I__18546\ : LocalMux
    port map (
            O => \N__74649\,
            I => \aluParams_1\
        );

    \I__18545\ : LocalMux
    port map (
            O => \N__74646\,
            I => \aluParams_1\
        );

    \I__18544\ : Odrv12
    port map (
            O => \N__74643\,
            I => \aluParams_1\
        );

    \I__18543\ : Odrv4
    port map (
            O => \N__74636\,
            I => \aluParams_1\
        );

    \I__18542\ : Odrv4
    port map (
            O => \N__74629\,
            I => \aluParams_1\
        );

    \I__18541\ : InMux
    port map (
            O => \N__74618\,
            I => \N__74615\
        );

    \I__18540\ : LocalMux
    port map (
            O => \N__74615\,
            I => \N__74612\
        );

    \I__18539\ : Odrv12
    port map (
            O => \N__74612\,
            I => \ALU.un14_log_0_0_15\
        );

    \I__18538\ : InMux
    port map (
            O => \N__74609\,
            I => \N__74604\
        );

    \I__18537\ : InMux
    port map (
            O => \N__74608\,
            I => \N__74600\
        );

    \I__18536\ : InMux
    port map (
            O => \N__74607\,
            I => \N__74597\
        );

    \I__18535\ : LocalMux
    port map (
            O => \N__74604\,
            I => \N__74593\
        );

    \I__18534\ : InMux
    port map (
            O => \N__74603\,
            I => \N__74590\
        );

    \I__18533\ : LocalMux
    port map (
            O => \N__74600\,
            I => \N__74587\
        );

    \I__18532\ : LocalMux
    port map (
            O => \N__74597\,
            I => \N__74584\
        );

    \I__18531\ : InMux
    port map (
            O => \N__74596\,
            I => \N__74581\
        );

    \I__18530\ : Span4Mux_h
    port map (
            O => \N__74593\,
            I => \N__74578\
        );

    \I__18529\ : LocalMux
    port map (
            O => \N__74590\,
            I => \N__74575\
        );

    \I__18528\ : Span12Mux_v
    port map (
            O => \N__74587\,
            I => \N__74572\
        );

    \I__18527\ : Span4Mux_v
    port map (
            O => \N__74584\,
            I => \N__74566\
        );

    \I__18526\ : LocalMux
    port map (
            O => \N__74581\,
            I => \N__74563\
        );

    \I__18525\ : Span4Mux_h
    port map (
            O => \N__74578\,
            I => \N__74560\
        );

    \I__18524\ : Span12Mux_s11_h
    port map (
            O => \N__74575\,
            I => \N__74555\
        );

    \I__18523\ : Span12Mux_h
    port map (
            O => \N__74572\,
            I => \N__74555\
        );

    \I__18522\ : InMux
    port map (
            O => \N__74571\,
            I => \N__74548\
        );

    \I__18521\ : InMux
    port map (
            O => \N__74570\,
            I => \N__74548\
        );

    \I__18520\ : InMux
    port map (
            O => \N__74569\,
            I => \N__74548\
        );

    \I__18519\ : Span4Mux_v
    port map (
            O => \N__74566\,
            I => \N__74545\
        );

    \I__18518\ : Span4Mux_h
    port map (
            O => \N__74563\,
            I => \N__74542\
        );

    \I__18517\ : Span4Mux_h
    port map (
            O => \N__74560\,
            I => \N__74539\
        );

    \I__18516\ : Odrv12
    port map (
            O => \N__74555\,
            I => \ALU.status_19_14\
        );

    \I__18515\ : LocalMux
    port map (
            O => \N__74548\,
            I => \ALU.status_19_14\
        );

    \I__18514\ : Odrv4
    port map (
            O => \N__74545\,
            I => \ALU.status_19_14\
        );

    \I__18513\ : Odrv4
    port map (
            O => \N__74542\,
            I => \ALU.status_19_14\
        );

    \I__18512\ : Odrv4
    port map (
            O => \N__74539\,
            I => \ALU.status_19_14\
        );

    \I__18511\ : InMux
    port map (
            O => \N__74528\,
            I => \N__74525\
        );

    \I__18510\ : LocalMux
    port map (
            O => \N__74525\,
            I => \N__74521\
        );

    \I__18509\ : InMux
    port map (
            O => \N__74524\,
            I => \N__74518\
        );

    \I__18508\ : Span4Mux_h
    port map (
            O => \N__74521\,
            I => \N__74515\
        );

    \I__18507\ : LocalMux
    port map (
            O => \N__74518\,
            I => \N__74512\
        );

    \I__18506\ : Odrv4
    port map (
            O => \N__74515\,
            I => \ALU.N_586\
        );

    \I__18505\ : Odrv12
    port map (
            O => \N__74512\,
            I => \ALU.N_586\
        );

    \I__18504\ : InMux
    port map (
            O => \N__74507\,
            I => \N__74504\
        );

    \I__18503\ : LocalMux
    port map (
            O => \N__74504\,
            I => \PROM.ROMDATA.m331_am\
        );

    \I__18502\ : InMux
    port map (
            O => \N__74501\,
            I => \N__74498\
        );

    \I__18501\ : LocalMux
    port map (
            O => \N__74498\,
            I => \PROM.ROMDATA.m357_bm\
        );

    \I__18500\ : CascadeMux
    port map (
            O => \N__74495\,
            I => \PROM.ROMDATA.m357_am_cascade_\
        );

    \I__18499\ : InMux
    port map (
            O => \N__74492\,
            I => \N__74484\
        );

    \I__18498\ : InMux
    port map (
            O => \N__74491\,
            I => \N__74481\
        );

    \I__18497\ : InMux
    port map (
            O => \N__74490\,
            I => \N__74477\
        );

    \I__18496\ : InMux
    port map (
            O => \N__74489\,
            I => \N__74474\
        );

    \I__18495\ : InMux
    port map (
            O => \N__74488\,
            I => \N__74471\
        );

    \I__18494\ : InMux
    port map (
            O => \N__74487\,
            I => \N__74468\
        );

    \I__18493\ : LocalMux
    port map (
            O => \N__74484\,
            I => \N__74465\
        );

    \I__18492\ : LocalMux
    port map (
            O => \N__74481\,
            I => \N__74462\
        );

    \I__18491\ : InMux
    port map (
            O => \N__74480\,
            I => \N__74459\
        );

    \I__18490\ : LocalMux
    port map (
            O => \N__74477\,
            I => \N__74454\
        );

    \I__18489\ : LocalMux
    port map (
            O => \N__74474\,
            I => \N__74454\
        );

    \I__18488\ : LocalMux
    port map (
            O => \N__74471\,
            I => \N__74451\
        );

    \I__18487\ : LocalMux
    port map (
            O => \N__74468\,
            I => \N__74448\
        );

    \I__18486\ : Span4Mux_v
    port map (
            O => \N__74465\,
            I => \N__74444\
        );

    \I__18485\ : Span4Mux_v
    port map (
            O => \N__74462\,
            I => \N__74439\
        );

    \I__18484\ : LocalMux
    port map (
            O => \N__74459\,
            I => \N__74439\
        );

    \I__18483\ : Span4Mux_v
    port map (
            O => \N__74454\,
            I => \N__74434\
        );

    \I__18482\ : Span4Mux_v
    port map (
            O => \N__74451\,
            I => \N__74434\
        );

    \I__18481\ : Span4Mux_v
    port map (
            O => \N__74448\,
            I => \N__74431\
        );

    \I__18480\ : InMux
    port map (
            O => \N__74447\,
            I => \N__74428\
        );

    \I__18479\ : Span4Mux_v
    port map (
            O => \N__74444\,
            I => \N__74423\
        );

    \I__18478\ : Span4Mux_h
    port map (
            O => \N__74439\,
            I => \N__74423\
        );

    \I__18477\ : Span4Mux_h
    port map (
            O => \N__74434\,
            I => \N__74416\
        );

    \I__18476\ : Span4Mux_h
    port map (
            O => \N__74431\,
            I => \N__74416\
        );

    \I__18475\ : LocalMux
    port map (
            O => \N__74428\,
            I => \N__74416\
        );

    \I__18474\ : Odrv4
    port map (
            O => \N__74423\,
            I => \PROM.ROMDATA.m178\
        );

    \I__18473\ : Odrv4
    port map (
            O => \N__74416\,
            I => \PROM.ROMDATA.m178\
        );

    \I__18472\ : CascadeMux
    port map (
            O => \N__74411\,
            I => \N__74407\
        );

    \I__18471\ : InMux
    port map (
            O => \N__74410\,
            I => \N__74403\
        );

    \I__18470\ : InMux
    port map (
            O => \N__74407\,
            I => \N__74400\
        );

    \I__18469\ : InMux
    port map (
            O => \N__74406\,
            I => \N__74397\
        );

    \I__18468\ : LocalMux
    port map (
            O => \N__74403\,
            I => \N__74394\
        );

    \I__18467\ : LocalMux
    port map (
            O => \N__74400\,
            I => \N__74391\
        );

    \I__18466\ : LocalMux
    port map (
            O => \N__74397\,
            I => \N__74386\
        );

    \I__18465\ : Span12Mux_h
    port map (
            O => \N__74394\,
            I => \N__74386\
        );

    \I__18464\ : Span4Mux_v
    port map (
            O => \N__74391\,
            I => \N__74383\
        );

    \I__18463\ : Odrv12
    port map (
            O => \N__74386\,
            I => \PROM.ROMDATA.m287\
        );

    \I__18462\ : Odrv4
    port map (
            O => \N__74383\,
            I => \PROM.ROMDATA.m287\
        );

    \I__18461\ : InMux
    port map (
            O => \N__74378\,
            I => \N__74375\
        );

    \I__18460\ : LocalMux
    port map (
            O => \N__74375\,
            I => \N__74372\
        );

    \I__18459\ : Span4Mux_h
    port map (
            O => \N__74372\,
            I => \N__74369\
        );

    \I__18458\ : Span4Mux_h
    port map (
            O => \N__74369\,
            I => \N__74366\
        );

    \I__18457\ : Odrv4
    port map (
            O => \N__74366\,
            I => \PROM.ROMDATA.m294_ns\
        );

    \I__18456\ : CascadeMux
    port map (
            O => \N__74363\,
            I => \PROM.ROMDATA.m290_cascade_\
        );

    \I__18455\ : CascadeMux
    port map (
            O => \N__74360\,
            I => \N__74357\
        );

    \I__18454\ : InMux
    port map (
            O => \N__74357\,
            I => \N__74354\
        );

    \I__18453\ : LocalMux
    port map (
            O => \N__74354\,
            I => \N__74351\
        );

    \I__18452\ : Odrv4
    port map (
            O => \N__74351\,
            I => \PROM.ROMDATA.m303_ns_1\
        );

    \I__18451\ : InMux
    port map (
            O => \N__74348\,
            I => \N__74345\
        );

    \I__18450\ : LocalMux
    port map (
            O => \N__74345\,
            I => \N__74342\
        );

    \I__18449\ : Odrv4
    port map (
            O => \N__74342\,
            I => \PROM.ROMDATA.m361_ns\
        );

    \I__18448\ : CascadeMux
    port map (
            O => \N__74339\,
            I => \N__74336\
        );

    \I__18447\ : InMux
    port map (
            O => \N__74336\,
            I => \N__74333\
        );

    \I__18446\ : LocalMux
    port map (
            O => \N__74333\,
            I => \PROM.ROMDATA.m357_ns\
        );

    \I__18445\ : InMux
    port map (
            O => \N__74330\,
            I => \N__74324\
        );

    \I__18444\ : InMux
    port map (
            O => \N__74329\,
            I => \N__74324\
        );

    \I__18443\ : LocalMux
    port map (
            O => \N__74324\,
            I => \N__74321\
        );

    \I__18442\ : Sp12to4
    port map (
            O => \N__74321\,
            I => \N__74318\
        );

    \I__18441\ : Span12Mux_h
    port map (
            O => \N__74318\,
            I => \N__74315\
        );

    \I__18440\ : Odrv12
    port map (
            O => \N__74315\,
            I => \PROM.ROMDATA.m363_ns\
        );

    \I__18439\ : CascadeMux
    port map (
            O => \N__74312\,
            I => \PROM.ROMDATA.m353_am_cascade_\
        );

    \I__18438\ : InMux
    port map (
            O => \N__74309\,
            I => \N__74306\
        );

    \I__18437\ : LocalMux
    port map (
            O => \N__74306\,
            I => \N__74303\
        );

    \I__18436\ : Span4Mux_v
    port map (
            O => \N__74303\,
            I => \N__74300\
        );

    \I__18435\ : Span4Mux_h
    port map (
            O => \N__74300\,
            I => \N__74297\
        );

    \I__18434\ : Odrv4
    port map (
            O => \N__74297\,
            I => \PROM.ROMDATA.m353_bm\
        );

    \I__18433\ : CascadeMux
    port map (
            O => \N__74294\,
            I => \PROM.ROMDATA.m353_ns_cascade_\
        );

    \I__18432\ : InMux
    port map (
            O => \N__74291\,
            I => \N__74288\
        );

    \I__18431\ : LocalMux
    port map (
            O => \N__74288\,
            I => \PROM.ROMDATA.m363_ns_1\
        );

    \I__18430\ : CascadeMux
    port map (
            O => \N__74285\,
            I => \N__74282\
        );

    \I__18429\ : InMux
    port map (
            O => \N__74282\,
            I => \N__74279\
        );

    \I__18428\ : LocalMux
    port map (
            O => \N__74279\,
            I => \N__74276\
        );

    \I__18427\ : Span4Mux_v
    port map (
            O => \N__74276\,
            I => \N__74273\
        );

    \I__18426\ : Odrv4
    port map (
            O => \N__74273\,
            I => \PROM.ROMDATA.m373\
        );

    \I__18425\ : InMux
    port map (
            O => \N__74270\,
            I => \N__74267\
        );

    \I__18424\ : LocalMux
    port map (
            O => \N__74267\,
            I => \N__74264\
        );

    \I__18423\ : Span4Mux_v
    port map (
            O => \N__74264\,
            I => \N__74261\
        );

    \I__18422\ : Odrv4
    port map (
            O => \N__74261\,
            I => \PROM.ROMDATA.m298_ns\
        );

    \I__18421\ : InMux
    port map (
            O => \N__74258\,
            I => \N__74255\
        );

    \I__18420\ : LocalMux
    port map (
            O => \N__74255\,
            I => \N__74252\
        );

    \I__18419\ : Span4Mux_h
    port map (
            O => \N__74252\,
            I => \N__74249\
        );

    \I__18418\ : Odrv4
    port map (
            O => \N__74249\,
            I => \PROM.ROMDATA.m303_ns\
        );

    \I__18417\ : InMux
    port map (
            O => \N__74246\,
            I => \N__74243\
        );

    \I__18416\ : LocalMux
    port map (
            O => \N__74243\,
            I => \N__74240\
        );

    \I__18415\ : Span4Mux_v
    port map (
            O => \N__74240\,
            I => \N__74236\
        );

    \I__18414\ : InMux
    port map (
            O => \N__74239\,
            I => \N__74233\
        );

    \I__18413\ : Span4Mux_h
    port map (
            O => \N__74236\,
            I => \N__74230\
        );

    \I__18412\ : LocalMux
    port map (
            O => \N__74233\,
            I => \PROM.ROMDATA.m262\
        );

    \I__18411\ : Odrv4
    port map (
            O => \N__74230\,
            I => \PROM.ROMDATA.m262\
        );

    \I__18410\ : InMux
    port map (
            O => \N__74225\,
            I => \N__74222\
        );

    \I__18409\ : LocalMux
    port map (
            O => \N__74222\,
            I => \N__74219\
        );

    \I__18408\ : Span4Mux_h
    port map (
            O => \N__74219\,
            I => \N__74216\
        );

    \I__18407\ : Odrv4
    port map (
            O => \N__74216\,
            I => \PROM.ROMDATA.m422_ns\
        );

    \I__18406\ : InMux
    port map (
            O => \N__74213\,
            I => \N__74207\
        );

    \I__18405\ : InMux
    port map (
            O => \N__74212\,
            I => \N__74207\
        );

    \I__18404\ : LocalMux
    port map (
            O => \N__74207\,
            I => \N__74204\
        );

    \I__18403\ : Span4Mux_h
    port map (
            O => \N__74204\,
            I => \N__74201\
        );

    \I__18402\ : Span4Mux_h
    port map (
            O => \N__74201\,
            I => \N__74198\
        );

    \I__18401\ : Span4Mux_h
    port map (
            O => \N__74198\,
            I => \N__74195\
        );

    \I__18400\ : Odrv4
    port map (
            O => \N__74195\,
            I => \PROM.ROMDATA.m424\
        );

    \I__18399\ : InMux
    port map (
            O => \N__74192\,
            I => \N__74189\
        );

    \I__18398\ : LocalMux
    port map (
            O => \N__74189\,
            I => \PROM.ROMDATA.m361_bm\
        );

    \I__18397\ : InMux
    port map (
            O => \N__74186\,
            I => \N__74182\
        );

    \I__18396\ : InMux
    port map (
            O => \N__74185\,
            I => \N__74179\
        );

    \I__18395\ : LocalMux
    port map (
            O => \N__74182\,
            I => \N__74176\
        );

    \I__18394\ : LocalMux
    port map (
            O => \N__74179\,
            I => \PROM.ROMDATA.m127\
        );

    \I__18393\ : Odrv12
    port map (
            O => \N__74176\,
            I => \PROM.ROMDATA.m127\
        );

    \I__18392\ : InMux
    port map (
            O => \N__74171\,
            I => \N__74168\
        );

    \I__18391\ : LocalMux
    port map (
            O => \N__74168\,
            I => \PROM.ROMDATA.m128\
        );

    \I__18390\ : CascadeMux
    port map (
            O => \N__74165\,
            I => \PROM.ROMDATA.m137_am_cascade_\
        );

    \I__18389\ : InMux
    port map (
            O => \N__74162\,
            I => \N__74159\
        );

    \I__18388\ : LocalMux
    port map (
            O => \N__74159\,
            I => \PROM.ROMDATA.m137_bm\
        );

    \I__18387\ : InMux
    port map (
            O => \N__74156\,
            I => \N__74153\
        );

    \I__18386\ : LocalMux
    port map (
            O => \N__74153\,
            I => \PROM.ROMDATA.m147_am\
        );

    \I__18385\ : InMux
    port map (
            O => \N__74150\,
            I => \N__74147\
        );

    \I__18384\ : LocalMux
    port map (
            O => \N__74147\,
            I => \N__74144\
        );

    \I__18383\ : Odrv4
    port map (
            O => \N__74144\,
            I => \PROM.ROMDATA.m147_bm\
        );

    \I__18382\ : CascadeMux
    port map (
            O => \N__74141\,
            I => \PROM.ROMDATA.m148_ns_1_cascade_\
        );

    \I__18381\ : InMux
    port map (
            O => \N__74138\,
            I => \N__74135\
        );

    \I__18380\ : LocalMux
    port map (
            O => \N__74135\,
            I => \N__74132\
        );

    \I__18379\ : Odrv12
    port map (
            O => \N__74132\,
            I => \PROM.ROMDATA.m148_ns\
        );

    \I__18378\ : InMux
    port map (
            O => \N__74129\,
            I => \N__74126\
        );

    \I__18377\ : LocalMux
    port map (
            O => \N__74126\,
            I => \N__74122\
        );

    \I__18376\ : InMux
    port map (
            O => \N__74125\,
            I => \N__74119\
        );

    \I__18375\ : Span4Mux_v
    port map (
            O => \N__74122\,
            I => \N__74116\
        );

    \I__18374\ : LocalMux
    port map (
            O => \N__74119\,
            I => \N__74111\
        );

    \I__18373\ : Span4Mux_h
    port map (
            O => \N__74116\,
            I => \N__74111\
        );

    \I__18372\ : Odrv4
    port map (
            O => \N__74111\,
            I => \PROM.ROMDATA.m292\
        );

    \I__18371\ : CascadeMux
    port map (
            O => \N__74108\,
            I => \N__74105\
        );

    \I__18370\ : InMux
    port map (
            O => \N__74105\,
            I => \N__74102\
        );

    \I__18369\ : LocalMux
    port map (
            O => \N__74102\,
            I => \N__74099\
        );

    \I__18368\ : Span12Mux_v
    port map (
            O => \N__74099\,
            I => \N__74096\
        );

    \I__18367\ : Odrv12
    port map (
            O => \N__74096\,
            I => \PROM.ROMDATA.m299\
        );

    \I__18366\ : InMux
    port map (
            O => \N__74093\,
            I => \N__74090\
        );

    \I__18365\ : LocalMux
    port map (
            O => \N__74090\,
            I => \PROM.ROMDATA.m301\
        );

    \I__18364\ : InMux
    port map (
            O => \N__74087\,
            I => \N__74084\
        );

    \I__18363\ : LocalMux
    port map (
            O => \N__74084\,
            I => \N__74081\
        );

    \I__18362\ : Span4Mux_v
    port map (
            O => \N__74081\,
            I => \N__74078\
        );

    \I__18361\ : Span4Mux_h
    port map (
            O => \N__74078\,
            I => \N__74075\
        );

    \I__18360\ : Odrv4
    port map (
            O => \N__74075\,
            I => \PROM.ROMDATA.m488_ns_1\
        );

    \I__18359\ : InMux
    port map (
            O => \N__74072\,
            I => \N__74062\
        );

    \I__18358\ : InMux
    port map (
            O => \N__74071\,
            I => \N__74058\
        );

    \I__18357\ : InMux
    port map (
            O => \N__74070\,
            I => \N__74053\
        );

    \I__18356\ : InMux
    port map (
            O => \N__74069\,
            I => \N__74053\
        );

    \I__18355\ : InMux
    port map (
            O => \N__74068\,
            I => \N__74050\
        );

    \I__18354\ : InMux
    port map (
            O => \N__74067\,
            I => \N__74045\
        );

    \I__18353\ : InMux
    port map (
            O => \N__74066\,
            I => \N__74045\
        );

    \I__18352\ : InMux
    port map (
            O => \N__74065\,
            I => \N__74042\
        );

    \I__18351\ : LocalMux
    port map (
            O => \N__74062\,
            I => \N__74039\
        );

    \I__18350\ : InMux
    port map (
            O => \N__74061\,
            I => \N__74034\
        );

    \I__18349\ : LocalMux
    port map (
            O => \N__74058\,
            I => \N__74031\
        );

    \I__18348\ : LocalMux
    port map (
            O => \N__74053\,
            I => \N__74024\
        );

    \I__18347\ : LocalMux
    port map (
            O => \N__74050\,
            I => \N__74024\
        );

    \I__18346\ : LocalMux
    port map (
            O => \N__74045\,
            I => \N__74024\
        );

    \I__18345\ : LocalMux
    port map (
            O => \N__74042\,
            I => \N__74020\
        );

    \I__18344\ : Span4Mux_v
    port map (
            O => \N__74039\,
            I => \N__74017\
        );

    \I__18343\ : InMux
    port map (
            O => \N__74038\,
            I => \N__74012\
        );

    \I__18342\ : InMux
    port map (
            O => \N__74037\,
            I => \N__74012\
        );

    \I__18341\ : LocalMux
    port map (
            O => \N__74034\,
            I => \N__74008\
        );

    \I__18340\ : Span4Mux_v
    port map (
            O => \N__74031\,
            I => \N__74004\
        );

    \I__18339\ : Span4Mux_v
    port map (
            O => \N__74024\,
            I => \N__74001\
        );

    \I__18338\ : InMux
    port map (
            O => \N__74023\,
            I => \N__73998\
        );

    \I__18337\ : Span4Mux_v
    port map (
            O => \N__74020\,
            I => \N__73994\
        );

    \I__18336\ : Span4Mux_h
    port map (
            O => \N__74017\,
            I => \N__73989\
        );

    \I__18335\ : LocalMux
    port map (
            O => \N__74012\,
            I => \N__73989\
        );

    \I__18334\ : InMux
    port map (
            O => \N__74011\,
            I => \N__73986\
        );

    \I__18333\ : Span4Mux_v
    port map (
            O => \N__74008\,
            I => \N__73983\
        );

    \I__18332\ : InMux
    port map (
            O => \N__74007\,
            I => \N__73980\
        );

    \I__18331\ : Span4Mux_h
    port map (
            O => \N__74004\,
            I => \N__73977\
        );

    \I__18330\ : Span4Mux_h
    port map (
            O => \N__74001\,
            I => \N__73972\
        );

    \I__18329\ : LocalMux
    port map (
            O => \N__73998\,
            I => \N__73972\
        );

    \I__18328\ : InMux
    port map (
            O => \N__73997\,
            I => \N__73969\
        );

    \I__18327\ : Span4Mux_h
    port map (
            O => \N__73994\,
            I => \N__73964\
        );

    \I__18326\ : Span4Mux_h
    port map (
            O => \N__73989\,
            I => \N__73964\
        );

    \I__18325\ : LocalMux
    port map (
            O => \N__73986\,
            I => \N__73959\
        );

    \I__18324\ : Span4Mux_h
    port map (
            O => \N__73983\,
            I => \N__73959\
        );

    \I__18323\ : LocalMux
    port map (
            O => \N__73980\,
            I => m125_e
        );

    \I__18322\ : Odrv4
    port map (
            O => \N__73977\,
            I => m125_e
        );

    \I__18321\ : Odrv4
    port map (
            O => \N__73972\,
            I => m125_e
        );

    \I__18320\ : LocalMux
    port map (
            O => \N__73969\,
            I => m125_e
        );

    \I__18319\ : Odrv4
    port map (
            O => \N__73964\,
            I => m125_e
        );

    \I__18318\ : Odrv4
    port map (
            O => \N__73959\,
            I => m125_e
        );

    \I__18317\ : CascadeMux
    port map (
            O => \N__73946\,
            I => \N__73942\
        );

    \I__18316\ : InMux
    port map (
            O => \N__73945\,
            I => \N__73937\
        );

    \I__18315\ : InMux
    port map (
            O => \N__73942\,
            I => \N__73937\
        );

    \I__18314\ : LocalMux
    port map (
            O => \N__73937\,
            I => \N__73934\
        );

    \I__18313\ : Span4Mux_v
    port map (
            O => \N__73934\,
            I => \N__73931\
        );

    \I__18312\ : Span4Mux_h
    port map (
            O => \N__73931\,
            I => \N__73928\
        );

    \I__18311\ : Span4Mux_h
    port map (
            O => \N__73928\,
            I => \N__73925\
        );

    \I__18310\ : Span4Mux_h
    port map (
            O => \N__73925\,
            I => \N__73922\
        );

    \I__18309\ : Odrv4
    port map (
            O => \N__73922\,
            I => \PROM.ROMDATA.N_570_mux\
        );

    \I__18308\ : CascadeMux
    port map (
            O => \N__73919\,
            I => \N__73915\
        );

    \I__18307\ : CascadeMux
    port map (
            O => \N__73918\,
            I => \N__73912\
        );

    \I__18306\ : InMux
    port map (
            O => \N__73915\,
            I => \N__73906\
        );

    \I__18305\ : InMux
    port map (
            O => \N__73912\,
            I => \N__73906\
        );

    \I__18304\ : CascadeMux
    port map (
            O => \N__73911\,
            I => \N__73902\
        );

    \I__18303\ : LocalMux
    port map (
            O => \N__73906\,
            I => \N__73899\
        );

    \I__18302\ : InMux
    port map (
            O => \N__73905\,
            I => \N__73896\
        );

    \I__18301\ : InMux
    port map (
            O => \N__73902\,
            I => \N__73893\
        );

    \I__18300\ : Span4Mux_v
    port map (
            O => \N__73899\,
            I => \N__73886\
        );

    \I__18299\ : LocalMux
    port map (
            O => \N__73896\,
            I => \N__73886\
        );

    \I__18298\ : LocalMux
    port map (
            O => \N__73893\,
            I => \N__73883\
        );

    \I__18297\ : CascadeMux
    port map (
            O => \N__73892\,
            I => \N__73880\
        );

    \I__18296\ : CascadeMux
    port map (
            O => \N__73891\,
            I => \N__73877\
        );

    \I__18295\ : Span4Mux_v
    port map (
            O => \N__73886\,
            I => \N__73874\
        );

    \I__18294\ : Span4Mux_h
    port map (
            O => \N__73883\,
            I => \N__73870\
        );

    \I__18293\ : InMux
    port map (
            O => \N__73880\,
            I => \N__73867\
        );

    \I__18292\ : InMux
    port map (
            O => \N__73877\,
            I => \N__73864\
        );

    \I__18291\ : Span4Mux_h
    port map (
            O => \N__73874\,
            I => \N__73861\
        );

    \I__18290\ : CascadeMux
    port map (
            O => \N__73873\,
            I => \N__73858\
        );

    \I__18289\ : Span4Mux_v
    port map (
            O => \N__73870\,
            I => \N__73852\
        );

    \I__18288\ : LocalMux
    port map (
            O => \N__73867\,
            I => \N__73852\
        );

    \I__18287\ : LocalMux
    port map (
            O => \N__73864\,
            I => \N__73849\
        );

    \I__18286\ : Span4Mux_h
    port map (
            O => \N__73861\,
            I => \N__73846\
        );

    \I__18285\ : InMux
    port map (
            O => \N__73858\,
            I => \N__73841\
        );

    \I__18284\ : InMux
    port map (
            O => \N__73857\,
            I => \N__73841\
        );

    \I__18283\ : Span4Mux_h
    port map (
            O => \N__73852\,
            I => \N__73838\
        );

    \I__18282\ : Odrv12
    port map (
            O => \N__73849\,
            I => \PROM.ROMDATA.m2\
        );

    \I__18281\ : Odrv4
    port map (
            O => \N__73846\,
            I => \PROM.ROMDATA.m2\
        );

    \I__18280\ : LocalMux
    port map (
            O => \N__73841\,
            I => \PROM.ROMDATA.m2\
        );

    \I__18279\ : Odrv4
    port map (
            O => \N__73838\,
            I => \PROM.ROMDATA.m2\
        );

    \I__18278\ : InMux
    port map (
            O => \N__73829\,
            I => \N__73826\
        );

    \I__18277\ : LocalMux
    port map (
            O => \N__73826\,
            I => \N__73823\
        );

    \I__18276\ : Odrv4
    port map (
            O => \N__73823\,
            I => \PROM.ROMDATA.m493_am\
        );

    \I__18275\ : InMux
    port map (
            O => \N__73820\,
            I => \N__73817\
        );

    \I__18274\ : LocalMux
    port map (
            O => \N__73817\,
            I => \N__73814\
        );

    \I__18273\ : Span4Mux_v
    port map (
            O => \N__73814\,
            I => \N__73805\
        );

    \I__18272\ : InMux
    port map (
            O => \N__73813\,
            I => \N__73800\
        );

    \I__18271\ : InMux
    port map (
            O => \N__73812\,
            I => \N__73800\
        );

    \I__18270\ : InMux
    port map (
            O => \N__73811\,
            I => \N__73797\
        );

    \I__18269\ : InMux
    port map (
            O => \N__73810\,
            I => \N__73794\
        );

    \I__18268\ : InMux
    port map (
            O => \N__73809\,
            I => \N__73791\
        );

    \I__18267\ : InMux
    port map (
            O => \N__73808\,
            I => \N__73788\
        );

    \I__18266\ : Span4Mux_h
    port map (
            O => \N__73805\,
            I => \N__73784\
        );

    \I__18265\ : LocalMux
    port map (
            O => \N__73800\,
            I => \N__73781\
        );

    \I__18264\ : LocalMux
    port map (
            O => \N__73797\,
            I => \N__73778\
        );

    \I__18263\ : LocalMux
    port map (
            O => \N__73794\,
            I => \N__73773\
        );

    \I__18262\ : LocalMux
    port map (
            O => \N__73791\,
            I => \N__73773\
        );

    \I__18261\ : LocalMux
    port map (
            O => \N__73788\,
            I => \N__73770\
        );

    \I__18260\ : InMux
    port map (
            O => \N__73787\,
            I => \N__73767\
        );

    \I__18259\ : Span4Mux_h
    port map (
            O => \N__73784\,
            I => \N__73761\
        );

    \I__18258\ : Span4Mux_v
    port map (
            O => \N__73781\,
            I => \N__73761\
        );

    \I__18257\ : Span4Mux_v
    port map (
            O => \N__73778\,
            I => \N__73752\
        );

    \I__18256\ : Span4Mux_v
    port map (
            O => \N__73773\,
            I => \N__73752\
        );

    \I__18255\ : Span4Mux_v
    port map (
            O => \N__73770\,
            I => \N__73752\
        );

    \I__18254\ : LocalMux
    port map (
            O => \N__73767\,
            I => \N__73752\
        );

    \I__18253\ : InMux
    port map (
            O => \N__73766\,
            I => \N__73749\
        );

    \I__18252\ : Odrv4
    port map (
            O => \N__73761\,
            I => \CONTROL_addrstack_reto_1\
        );

    \I__18251\ : Odrv4
    port map (
            O => \N__73752\,
            I => \CONTROL_addrstack_reto_1\
        );

    \I__18250\ : LocalMux
    port map (
            O => \N__73749\,
            I => \CONTROL_addrstack_reto_1\
        );

    \I__18249\ : CascadeMux
    port map (
            O => \N__73742\,
            I => \N__73737\
        );

    \I__18248\ : CascadeMux
    port map (
            O => \N__73741\,
            I => \N__73734\
        );

    \I__18247\ : CascadeMux
    port map (
            O => \N__73740\,
            I => \N__73731\
        );

    \I__18246\ : InMux
    port map (
            O => \N__73737\,
            I => \N__73725\
        );

    \I__18245\ : InMux
    port map (
            O => \N__73734\,
            I => \N__73722\
        );

    \I__18244\ : InMux
    port map (
            O => \N__73731\,
            I => \N__73716\
        );

    \I__18243\ : CascadeMux
    port map (
            O => \N__73730\,
            I => \N__73713\
        );

    \I__18242\ : InMux
    port map (
            O => \N__73729\,
            I => \N__73707\
        );

    \I__18241\ : InMux
    port map (
            O => \N__73728\,
            I => \N__73707\
        );

    \I__18240\ : LocalMux
    port map (
            O => \N__73725\,
            I => \N__73702\
        );

    \I__18239\ : LocalMux
    port map (
            O => \N__73722\,
            I => \N__73702\
        );

    \I__18238\ : InMux
    port map (
            O => \N__73721\,
            I => \N__73697\
        );

    \I__18237\ : InMux
    port map (
            O => \N__73720\,
            I => \N__73697\
        );

    \I__18236\ : CascadeMux
    port map (
            O => \N__73719\,
            I => \N__73694\
        );

    \I__18235\ : LocalMux
    port map (
            O => \N__73716\,
            I => \N__73691\
        );

    \I__18234\ : InMux
    port map (
            O => \N__73713\,
            I => \N__73688\
        );

    \I__18233\ : InMux
    port map (
            O => \N__73712\,
            I => \N__73683\
        );

    \I__18232\ : LocalMux
    port map (
            O => \N__73707\,
            I => \N__73680\
        );

    \I__18231\ : Span4Mux_v
    port map (
            O => \N__73702\,
            I => \N__73672\
        );

    \I__18230\ : LocalMux
    port map (
            O => \N__73697\,
            I => \N__73672\
        );

    \I__18229\ : InMux
    port map (
            O => \N__73694\,
            I => \N__73669\
        );

    \I__18228\ : Span4Mux_v
    port map (
            O => \N__73691\,
            I => \N__73665\
        );

    \I__18227\ : LocalMux
    port map (
            O => \N__73688\,
            I => \N__73662\
        );

    \I__18226\ : InMux
    port map (
            O => \N__73687\,
            I => \N__73658\
        );

    \I__18225\ : InMux
    port map (
            O => \N__73686\,
            I => \N__73655\
        );

    \I__18224\ : LocalMux
    port map (
            O => \N__73683\,
            I => \N__73652\
        );

    \I__18223\ : Span4Mux_v
    port map (
            O => \N__73680\,
            I => \N__73649\
        );

    \I__18222\ : InMux
    port map (
            O => \N__73679\,
            I => \N__73642\
        );

    \I__18221\ : InMux
    port map (
            O => \N__73678\,
            I => \N__73642\
        );

    \I__18220\ : InMux
    port map (
            O => \N__73677\,
            I => \N__73642\
        );

    \I__18219\ : Span4Mux_h
    port map (
            O => \N__73672\,
            I => \N__73637\
        );

    \I__18218\ : LocalMux
    port map (
            O => \N__73669\,
            I => \N__73637\
        );

    \I__18217\ : InMux
    port map (
            O => \N__73668\,
            I => \N__73633\
        );

    \I__18216\ : Span4Mux_h
    port map (
            O => \N__73665\,
            I => \N__73628\
        );

    \I__18215\ : Span4Mux_v
    port map (
            O => \N__73662\,
            I => \N__73628\
        );

    \I__18214\ : CascadeMux
    port map (
            O => \N__73661\,
            I => \N__73624\
        );

    \I__18213\ : LocalMux
    port map (
            O => \N__73658\,
            I => \N__73619\
        );

    \I__18212\ : LocalMux
    port map (
            O => \N__73655\,
            I => \N__73619\
        );

    \I__18211\ : Span4Mux_v
    port map (
            O => \N__73652\,
            I => \N__73614\
        );

    \I__18210\ : Span4Mux_h
    port map (
            O => \N__73649\,
            I => \N__73614\
        );

    \I__18209\ : LocalMux
    port map (
            O => \N__73642\,
            I => \N__73611\
        );

    \I__18208\ : Span4Mux_v
    port map (
            O => \N__73637\,
            I => \N__73608\
        );

    \I__18207\ : InMux
    port map (
            O => \N__73636\,
            I => \N__73605\
        );

    \I__18206\ : LocalMux
    port map (
            O => \N__73633\,
            I => \N__73600\
        );

    \I__18205\ : Sp12to4
    port map (
            O => \N__73628\,
            I => \N__73600\
        );

    \I__18204\ : InMux
    port map (
            O => \N__73627\,
            I => \N__73595\
        );

    \I__18203\ : InMux
    port map (
            O => \N__73624\,
            I => \N__73595\
        );

    \I__18202\ : Span4Mux_v
    port map (
            O => \N__73619\,
            I => \N__73588\
        );

    \I__18201\ : Span4Mux_h
    port map (
            O => \N__73614\,
            I => \N__73588\
        );

    \I__18200\ : Span4Mux_v
    port map (
            O => \N__73611\,
            I => \N__73588\
        );

    \I__18199\ : Span4Mux_h
    port map (
            O => \N__73608\,
            I => \N__73585\
        );

    \I__18198\ : LocalMux
    port map (
            O => \N__73605\,
            I => \CONTROL_programCounter11_reto\
        );

    \I__18197\ : Odrv12
    port map (
            O => \N__73600\,
            I => \CONTROL_programCounter11_reto\
        );

    \I__18196\ : LocalMux
    port map (
            O => \N__73595\,
            I => \CONTROL_programCounter11_reto\
        );

    \I__18195\ : Odrv4
    port map (
            O => \N__73588\,
            I => \CONTROL_programCounter11_reto\
        );

    \I__18194\ : Odrv4
    port map (
            O => \N__73585\,
            I => \CONTROL_programCounter11_reto\
        );

    \I__18193\ : InMux
    port map (
            O => \N__73574\,
            I => \N__73569\
        );

    \I__18192\ : CascadeMux
    port map (
            O => \N__73573\,
            I => \N__73566\
        );

    \I__18191\ : InMux
    port map (
            O => \N__73572\,
            I => \N__73562\
        );

    \I__18190\ : LocalMux
    port map (
            O => \N__73569\,
            I => \N__73559\
        );

    \I__18189\ : InMux
    port map (
            O => \N__73566\,
            I => \N__73554\
        );

    \I__18188\ : InMux
    port map (
            O => \N__73565\,
            I => \N__73554\
        );

    \I__18187\ : LocalMux
    port map (
            O => \N__73562\,
            I => \N__73549\
        );

    \I__18186\ : Span4Mux_v
    port map (
            O => \N__73559\,
            I => \N__73546\
        );

    \I__18185\ : LocalMux
    port map (
            O => \N__73554\,
            I => \N__73543\
        );

    \I__18184\ : InMux
    port map (
            O => \N__73553\,
            I => \N__73539\
        );

    \I__18183\ : InMux
    port map (
            O => \N__73552\,
            I => \N__73536\
        );

    \I__18182\ : Span4Mux_v
    port map (
            O => \N__73549\,
            I => \N__73533\
        );

    \I__18181\ : Sp12to4
    port map (
            O => \N__73546\,
            I => \N__73530\
        );

    \I__18180\ : Span4Mux_h
    port map (
            O => \N__73543\,
            I => \N__73527\
        );

    \I__18179\ : InMux
    port map (
            O => \N__73542\,
            I => \N__73524\
        );

    \I__18178\ : LocalMux
    port map (
            O => \N__73539\,
            I => \N__73519\
        );

    \I__18177\ : LocalMux
    port map (
            O => \N__73536\,
            I => \N__73519\
        );

    \I__18176\ : Span4Mux_h
    port map (
            O => \N__73533\,
            I => \N__73516\
        );

    \I__18175\ : Odrv12
    port map (
            O => \N__73530\,
            I => \N_416\
        );

    \I__18174\ : Odrv4
    port map (
            O => \N__73527\,
            I => \N_416\
        );

    \I__18173\ : LocalMux
    port map (
            O => \N__73524\,
            I => \N_416\
        );

    \I__18172\ : Odrv4
    port map (
            O => \N__73519\,
            I => \N_416\
        );

    \I__18171\ : Odrv4
    port map (
            O => \N__73516\,
            I => \N_416\
        );

    \I__18170\ : InMux
    port map (
            O => \N__73505\,
            I => \N__73498\
        );

    \I__18169\ : InMux
    port map (
            O => \N__73504\,
            I => \N__73498\
        );

    \I__18168\ : InMux
    port map (
            O => \N__73503\,
            I => \N__73495\
        );

    \I__18167\ : LocalMux
    port map (
            O => \N__73498\,
            I => \N__73492\
        );

    \I__18166\ : LocalMux
    port map (
            O => \N__73495\,
            I => \N__73488\
        );

    \I__18165\ : Span4Mux_h
    port map (
            O => \N__73492\,
            I => \N__73485\
        );

    \I__18164\ : InMux
    port map (
            O => \N__73491\,
            I => \N__73482\
        );

    \I__18163\ : Span4Mux_h
    port map (
            O => \N__73488\,
            I => \N__73475\
        );

    \I__18162\ : Span4Mux_h
    port map (
            O => \N__73485\,
            I => \N__73475\
        );

    \I__18161\ : LocalMux
    port map (
            O => \N__73482\,
            I => \N__73475\
        );

    \I__18160\ : Span4Mux_v
    port map (
            O => \N__73475\,
            I => \N__73472\
        );

    \I__18159\ : Odrv4
    port map (
            O => \N__73472\,
            I => \PROM.ROMDATA.m1\
        );

    \I__18158\ : CascadeMux
    port map (
            O => \N__73469\,
            I => \N__73466\
        );

    \I__18157\ : InMux
    port map (
            O => \N__73466\,
            I => \N__73463\
        );

    \I__18156\ : LocalMux
    port map (
            O => \N__73463\,
            I => \N__73460\
        );

    \I__18155\ : Span4Mux_h
    port map (
            O => \N__73460\,
            I => \N__73457\
        );

    \I__18154\ : Odrv4
    port map (
            O => \N__73457\,
            I => \PROM.ROMDATA.m493_bm\
        );

    \I__18153\ : InMux
    port map (
            O => \N__73454\,
            I => \N__73451\
        );

    \I__18152\ : LocalMux
    port map (
            O => \N__73451\,
            I => \PROM.ROMDATA.m361_am\
        );

    \I__18151\ : CascadeMux
    port map (
            O => \N__73448\,
            I => \N__73445\
        );

    \I__18150\ : InMux
    port map (
            O => \N__73445\,
            I => \N__73442\
        );

    \I__18149\ : LocalMux
    port map (
            O => \N__73442\,
            I => \N__73439\
        );

    \I__18148\ : Odrv4
    port map (
            O => \N__73439\,
            I => \PROM.ROMDATA.m211_ns_N_2L1\
        );

    \I__18147\ : CascadeMux
    port map (
            O => \N__73436\,
            I => \PROM.ROMDATA.m211_ns_cascade_\
        );

    \I__18146\ : InMux
    port map (
            O => \N__73433\,
            I => \N__73430\
        );

    \I__18145\ : LocalMux
    port map (
            O => \N__73430\,
            I => \N__73427\
        );

    \I__18144\ : Span4Mux_h
    port map (
            O => \N__73427\,
            I => \N__73424\
        );

    \I__18143\ : Span4Mux_h
    port map (
            O => \N__73424\,
            I => \N__73421\
        );

    \I__18142\ : Odrv4
    port map (
            O => \N__73421\,
            I => \PROM.ROMDATA.m221cf0_1\
        );

    \I__18141\ : InMux
    port map (
            O => \N__73418\,
            I => \N__73415\
        );

    \I__18140\ : LocalMux
    port map (
            O => \N__73415\,
            I => \PROM.ROMDATA.m211_ns\
        );

    \I__18139\ : CascadeMux
    port map (
            O => \N__73412\,
            I => \N__73409\
        );

    \I__18138\ : InMux
    port map (
            O => \N__73409\,
            I => \N__73406\
        );

    \I__18137\ : LocalMux
    port map (
            O => \N__73406\,
            I => \N__73403\
        );

    \I__18136\ : Span4Mux_v
    port map (
            O => \N__73403\,
            I => \N__73400\
        );

    \I__18135\ : Sp12to4
    port map (
            O => \N__73400\,
            I => \N__73397\
        );

    \I__18134\ : Odrv12
    port map (
            O => \N__73397\,
            I => \PROM.ROMDATA.m221cf1_1\
        );

    \I__18133\ : CascadeMux
    port map (
            O => \N__73394\,
            I => \N__73391\
        );

    \I__18132\ : InMux
    port map (
            O => \N__73391\,
            I => \N__73388\
        );

    \I__18131\ : LocalMux
    port map (
            O => \N__73388\,
            I => \N__73385\
        );

    \I__18130\ : Span4Mux_v
    port map (
            O => \N__73385\,
            I => \N__73382\
        );

    \I__18129\ : Span4Mux_h
    port map (
            O => \N__73382\,
            I => \N__73379\
        );

    \I__18128\ : Sp12to4
    port map (
            O => \N__73379\,
            I => \N__73376\
        );

    \I__18127\ : Odrv12
    port map (
            O => \N__73376\,
            I => \PROM.ROMDATA.m369\
        );

    \I__18126\ : CascadeMux
    port map (
            O => \N__73373\,
            I => \N__73370\
        );

    \I__18125\ : InMux
    port map (
            O => \N__73370\,
            I => \N__73367\
        );

    \I__18124\ : LocalMux
    port map (
            O => \N__73367\,
            I => \N__73364\
        );

    \I__18123\ : Span4Mux_h
    port map (
            O => \N__73364\,
            I => \N__73361\
        );

    \I__18122\ : Span4Mux_v
    port map (
            O => \N__73361\,
            I => \N__73358\
        );

    \I__18121\ : Odrv4
    port map (
            O => \N__73358\,
            I => \PROM.ROMDATA.m60\
        );

    \I__18120\ : InMux
    port map (
            O => \N__73355\,
            I => \N__73352\
        );

    \I__18119\ : LocalMux
    port map (
            O => \N__73352\,
            I => \N__73349\
        );

    \I__18118\ : Span4Mux_v
    port map (
            O => \N__73349\,
            I => \N__73345\
        );

    \I__18117\ : InMux
    port map (
            O => \N__73348\,
            I => \N__73342\
        );

    \I__18116\ : Span4Mux_h
    port map (
            O => \N__73345\,
            I => \N__73339\
        );

    \I__18115\ : LocalMux
    port map (
            O => \N__73342\,
            I => \N__73336\
        );

    \I__18114\ : Span4Mux_h
    port map (
            O => \N__73339\,
            I => \N__73333\
        );

    \I__18113\ : Span4Mux_v
    port map (
            O => \N__73336\,
            I => \N__73330\
        );

    \I__18112\ : Span4Mux_h
    port map (
            O => \N__73333\,
            I => \N__73327\
        );

    \I__18111\ : Span4Mux_h
    port map (
            O => \N__73330\,
            I => \N__73324\
        );

    \I__18110\ : Odrv4
    port map (
            O => \N__73327\,
            I => \CONTROL.programCounter_1_7\
        );

    \I__18109\ : Odrv4
    port map (
            O => \N__73324\,
            I => \CONTROL.programCounter_1_7\
        );

    \I__18108\ : InMux
    port map (
            O => \N__73319\,
            I => \N__73316\
        );

    \I__18107\ : LocalMux
    port map (
            O => \N__73316\,
            I => \N__73313\
        );

    \I__18106\ : Span4Mux_h
    port map (
            O => \N__73313\,
            I => \N__73310\
        );

    \I__18105\ : Span4Mux_h
    port map (
            O => \N__73310\,
            I => \N__73307\
        );

    \I__18104\ : Odrv4
    port map (
            O => \N__73307\,
            I => \CONTROL.programCounter_1_reto_7\
        );

    \I__18103\ : InMux
    port map (
            O => \N__73304\,
            I => \N__73299\
        );

    \I__18102\ : InMux
    port map (
            O => \N__73303\,
            I => \N__73294\
        );

    \I__18101\ : InMux
    port map (
            O => \N__73302\,
            I => \N__73294\
        );

    \I__18100\ : LocalMux
    port map (
            O => \N__73299\,
            I => \N__73287\
        );

    \I__18099\ : LocalMux
    port map (
            O => \N__73294\,
            I => \N__73283\
        );

    \I__18098\ : ClkMux
    port map (
            O => \N__73293\,
            I => \N__72833\
        );

    \I__18097\ : ClkMux
    port map (
            O => \N__73292\,
            I => \N__72833\
        );

    \I__18096\ : ClkMux
    port map (
            O => \N__73291\,
            I => \N__72833\
        );

    \I__18095\ : ClkMux
    port map (
            O => \N__73290\,
            I => \N__72833\
        );

    \I__18094\ : Glb2LocalMux
    port map (
            O => \N__73287\,
            I => \N__72833\
        );

    \I__18093\ : ClkMux
    port map (
            O => \N__73286\,
            I => \N__72833\
        );

    \I__18092\ : Glb2LocalMux
    port map (
            O => \N__73283\,
            I => \N__72833\
        );

    \I__18091\ : ClkMux
    port map (
            O => \N__73282\,
            I => \N__72833\
        );

    \I__18090\ : ClkMux
    port map (
            O => \N__73281\,
            I => \N__72833\
        );

    \I__18089\ : ClkMux
    port map (
            O => \N__73280\,
            I => \N__72833\
        );

    \I__18088\ : ClkMux
    port map (
            O => \N__73279\,
            I => \N__72833\
        );

    \I__18087\ : ClkMux
    port map (
            O => \N__73278\,
            I => \N__72833\
        );

    \I__18086\ : ClkMux
    port map (
            O => \N__73277\,
            I => \N__72833\
        );

    \I__18085\ : ClkMux
    port map (
            O => \N__73276\,
            I => \N__72833\
        );

    \I__18084\ : ClkMux
    port map (
            O => \N__73275\,
            I => \N__72833\
        );

    \I__18083\ : ClkMux
    port map (
            O => \N__73274\,
            I => \N__72833\
        );

    \I__18082\ : ClkMux
    port map (
            O => \N__73273\,
            I => \N__72833\
        );

    \I__18081\ : ClkMux
    port map (
            O => \N__73272\,
            I => \N__72833\
        );

    \I__18080\ : ClkMux
    port map (
            O => \N__73271\,
            I => \N__72833\
        );

    \I__18079\ : ClkMux
    port map (
            O => \N__73270\,
            I => \N__72833\
        );

    \I__18078\ : ClkMux
    port map (
            O => \N__73269\,
            I => \N__72833\
        );

    \I__18077\ : ClkMux
    port map (
            O => \N__73268\,
            I => \N__72833\
        );

    \I__18076\ : ClkMux
    port map (
            O => \N__73267\,
            I => \N__72833\
        );

    \I__18075\ : ClkMux
    port map (
            O => \N__73266\,
            I => \N__72833\
        );

    \I__18074\ : ClkMux
    port map (
            O => \N__73265\,
            I => \N__72833\
        );

    \I__18073\ : ClkMux
    port map (
            O => \N__73264\,
            I => \N__72833\
        );

    \I__18072\ : ClkMux
    port map (
            O => \N__73263\,
            I => \N__72833\
        );

    \I__18071\ : ClkMux
    port map (
            O => \N__73262\,
            I => \N__72833\
        );

    \I__18070\ : ClkMux
    port map (
            O => \N__73261\,
            I => \N__72833\
        );

    \I__18069\ : ClkMux
    port map (
            O => \N__73260\,
            I => \N__72833\
        );

    \I__18068\ : ClkMux
    port map (
            O => \N__73259\,
            I => \N__72833\
        );

    \I__18067\ : ClkMux
    port map (
            O => \N__73258\,
            I => \N__72833\
        );

    \I__18066\ : ClkMux
    port map (
            O => \N__73257\,
            I => \N__72833\
        );

    \I__18065\ : ClkMux
    port map (
            O => \N__73256\,
            I => \N__72833\
        );

    \I__18064\ : ClkMux
    port map (
            O => \N__73255\,
            I => \N__72833\
        );

    \I__18063\ : ClkMux
    port map (
            O => \N__73254\,
            I => \N__72833\
        );

    \I__18062\ : ClkMux
    port map (
            O => \N__73253\,
            I => \N__72833\
        );

    \I__18061\ : ClkMux
    port map (
            O => \N__73252\,
            I => \N__72833\
        );

    \I__18060\ : ClkMux
    port map (
            O => \N__73251\,
            I => \N__72833\
        );

    \I__18059\ : ClkMux
    port map (
            O => \N__73250\,
            I => \N__72833\
        );

    \I__18058\ : ClkMux
    port map (
            O => \N__73249\,
            I => \N__72833\
        );

    \I__18057\ : ClkMux
    port map (
            O => \N__73248\,
            I => \N__72833\
        );

    \I__18056\ : ClkMux
    port map (
            O => \N__73247\,
            I => \N__72833\
        );

    \I__18055\ : ClkMux
    port map (
            O => \N__73246\,
            I => \N__72833\
        );

    \I__18054\ : ClkMux
    port map (
            O => \N__73245\,
            I => \N__72833\
        );

    \I__18053\ : ClkMux
    port map (
            O => \N__73244\,
            I => \N__72833\
        );

    \I__18052\ : ClkMux
    port map (
            O => \N__73243\,
            I => \N__72833\
        );

    \I__18051\ : ClkMux
    port map (
            O => \N__73242\,
            I => \N__72833\
        );

    \I__18050\ : ClkMux
    port map (
            O => \N__73241\,
            I => \N__72833\
        );

    \I__18049\ : ClkMux
    port map (
            O => \N__73240\,
            I => \N__72833\
        );

    \I__18048\ : ClkMux
    port map (
            O => \N__73239\,
            I => \N__72833\
        );

    \I__18047\ : ClkMux
    port map (
            O => \N__73238\,
            I => \N__72833\
        );

    \I__18046\ : ClkMux
    port map (
            O => \N__73237\,
            I => \N__72833\
        );

    \I__18045\ : ClkMux
    port map (
            O => \N__73236\,
            I => \N__72833\
        );

    \I__18044\ : ClkMux
    port map (
            O => \N__73235\,
            I => \N__72833\
        );

    \I__18043\ : ClkMux
    port map (
            O => \N__73234\,
            I => \N__72833\
        );

    \I__18042\ : ClkMux
    port map (
            O => \N__73233\,
            I => \N__72833\
        );

    \I__18041\ : ClkMux
    port map (
            O => \N__73232\,
            I => \N__72833\
        );

    \I__18040\ : ClkMux
    port map (
            O => \N__73231\,
            I => \N__72833\
        );

    \I__18039\ : ClkMux
    port map (
            O => \N__73230\,
            I => \N__72833\
        );

    \I__18038\ : ClkMux
    port map (
            O => \N__73229\,
            I => \N__72833\
        );

    \I__18037\ : ClkMux
    port map (
            O => \N__73228\,
            I => \N__72833\
        );

    \I__18036\ : ClkMux
    port map (
            O => \N__73227\,
            I => \N__72833\
        );

    \I__18035\ : ClkMux
    port map (
            O => \N__73226\,
            I => \N__72833\
        );

    \I__18034\ : ClkMux
    port map (
            O => \N__73225\,
            I => \N__72833\
        );

    \I__18033\ : ClkMux
    port map (
            O => \N__73224\,
            I => \N__72833\
        );

    \I__18032\ : ClkMux
    port map (
            O => \N__73223\,
            I => \N__72833\
        );

    \I__18031\ : ClkMux
    port map (
            O => \N__73222\,
            I => \N__72833\
        );

    \I__18030\ : ClkMux
    port map (
            O => \N__73221\,
            I => \N__72833\
        );

    \I__18029\ : ClkMux
    port map (
            O => \N__73220\,
            I => \N__72833\
        );

    \I__18028\ : ClkMux
    port map (
            O => \N__73219\,
            I => \N__72833\
        );

    \I__18027\ : ClkMux
    port map (
            O => \N__73218\,
            I => \N__72833\
        );

    \I__18026\ : ClkMux
    port map (
            O => \N__73217\,
            I => \N__72833\
        );

    \I__18025\ : ClkMux
    port map (
            O => \N__73216\,
            I => \N__72833\
        );

    \I__18024\ : ClkMux
    port map (
            O => \N__73215\,
            I => \N__72833\
        );

    \I__18023\ : ClkMux
    port map (
            O => \N__73214\,
            I => \N__72833\
        );

    \I__18022\ : ClkMux
    port map (
            O => \N__73213\,
            I => \N__72833\
        );

    \I__18021\ : ClkMux
    port map (
            O => \N__73212\,
            I => \N__72833\
        );

    \I__18020\ : ClkMux
    port map (
            O => \N__73211\,
            I => \N__72833\
        );

    \I__18019\ : ClkMux
    port map (
            O => \N__73210\,
            I => \N__72833\
        );

    \I__18018\ : ClkMux
    port map (
            O => \N__73209\,
            I => \N__72833\
        );

    \I__18017\ : ClkMux
    port map (
            O => \N__73208\,
            I => \N__72833\
        );

    \I__18016\ : ClkMux
    port map (
            O => \N__73207\,
            I => \N__72833\
        );

    \I__18015\ : ClkMux
    port map (
            O => \N__73206\,
            I => \N__72833\
        );

    \I__18014\ : ClkMux
    port map (
            O => \N__73205\,
            I => \N__72833\
        );

    \I__18013\ : ClkMux
    port map (
            O => \N__73204\,
            I => \N__72833\
        );

    \I__18012\ : ClkMux
    port map (
            O => \N__73203\,
            I => \N__72833\
        );

    \I__18011\ : ClkMux
    port map (
            O => \N__73202\,
            I => \N__72833\
        );

    \I__18010\ : ClkMux
    port map (
            O => \N__73201\,
            I => \N__72833\
        );

    \I__18009\ : ClkMux
    port map (
            O => \N__73200\,
            I => \N__72833\
        );

    \I__18008\ : ClkMux
    port map (
            O => \N__73199\,
            I => \N__72833\
        );

    \I__18007\ : ClkMux
    port map (
            O => \N__73198\,
            I => \N__72833\
        );

    \I__18006\ : ClkMux
    port map (
            O => \N__73197\,
            I => \N__72833\
        );

    \I__18005\ : ClkMux
    port map (
            O => \N__73196\,
            I => \N__72833\
        );

    \I__18004\ : ClkMux
    port map (
            O => \N__73195\,
            I => \N__72833\
        );

    \I__18003\ : ClkMux
    port map (
            O => \N__73194\,
            I => \N__72833\
        );

    \I__18002\ : ClkMux
    port map (
            O => \N__73193\,
            I => \N__72833\
        );

    \I__18001\ : ClkMux
    port map (
            O => \N__73192\,
            I => \N__72833\
        );

    \I__18000\ : ClkMux
    port map (
            O => \N__73191\,
            I => \N__72833\
        );

    \I__17999\ : ClkMux
    port map (
            O => \N__73190\,
            I => \N__72833\
        );

    \I__17998\ : ClkMux
    port map (
            O => \N__73189\,
            I => \N__72833\
        );

    \I__17997\ : ClkMux
    port map (
            O => \N__73188\,
            I => \N__72833\
        );

    \I__17996\ : ClkMux
    port map (
            O => \N__73187\,
            I => \N__72833\
        );

    \I__17995\ : ClkMux
    port map (
            O => \N__73186\,
            I => \N__72833\
        );

    \I__17994\ : ClkMux
    port map (
            O => \N__73185\,
            I => \N__72833\
        );

    \I__17993\ : ClkMux
    port map (
            O => \N__73184\,
            I => \N__72833\
        );

    \I__17992\ : ClkMux
    port map (
            O => \N__73183\,
            I => \N__72833\
        );

    \I__17991\ : ClkMux
    port map (
            O => \N__73182\,
            I => \N__72833\
        );

    \I__17990\ : ClkMux
    port map (
            O => \N__73181\,
            I => \N__72833\
        );

    \I__17989\ : ClkMux
    port map (
            O => \N__73180\,
            I => \N__72833\
        );

    \I__17988\ : ClkMux
    port map (
            O => \N__73179\,
            I => \N__72833\
        );

    \I__17987\ : ClkMux
    port map (
            O => \N__73178\,
            I => \N__72833\
        );

    \I__17986\ : ClkMux
    port map (
            O => \N__73177\,
            I => \N__72833\
        );

    \I__17985\ : ClkMux
    port map (
            O => \N__73176\,
            I => \N__72833\
        );

    \I__17984\ : ClkMux
    port map (
            O => \N__73175\,
            I => \N__72833\
        );

    \I__17983\ : ClkMux
    port map (
            O => \N__73174\,
            I => \N__72833\
        );

    \I__17982\ : ClkMux
    port map (
            O => \N__73173\,
            I => \N__72833\
        );

    \I__17981\ : ClkMux
    port map (
            O => \N__73172\,
            I => \N__72833\
        );

    \I__17980\ : ClkMux
    port map (
            O => \N__73171\,
            I => \N__72833\
        );

    \I__17979\ : ClkMux
    port map (
            O => \N__73170\,
            I => \N__72833\
        );

    \I__17978\ : ClkMux
    port map (
            O => \N__73169\,
            I => \N__72833\
        );

    \I__17977\ : ClkMux
    port map (
            O => \N__73168\,
            I => \N__72833\
        );

    \I__17976\ : ClkMux
    port map (
            O => \N__73167\,
            I => \N__72833\
        );

    \I__17975\ : ClkMux
    port map (
            O => \N__73166\,
            I => \N__72833\
        );

    \I__17974\ : ClkMux
    port map (
            O => \N__73165\,
            I => \N__72833\
        );

    \I__17973\ : ClkMux
    port map (
            O => \N__73164\,
            I => \N__72833\
        );

    \I__17972\ : ClkMux
    port map (
            O => \N__73163\,
            I => \N__72833\
        );

    \I__17971\ : ClkMux
    port map (
            O => \N__73162\,
            I => \N__72833\
        );

    \I__17970\ : ClkMux
    port map (
            O => \N__73161\,
            I => \N__72833\
        );

    \I__17969\ : ClkMux
    port map (
            O => \N__73160\,
            I => \N__72833\
        );

    \I__17968\ : ClkMux
    port map (
            O => \N__73159\,
            I => \N__72833\
        );

    \I__17967\ : ClkMux
    port map (
            O => \N__73158\,
            I => \N__72833\
        );

    \I__17966\ : ClkMux
    port map (
            O => \N__73157\,
            I => \N__72833\
        );

    \I__17965\ : ClkMux
    port map (
            O => \N__73156\,
            I => \N__72833\
        );

    \I__17964\ : ClkMux
    port map (
            O => \N__73155\,
            I => \N__72833\
        );

    \I__17963\ : ClkMux
    port map (
            O => \N__73154\,
            I => \N__72833\
        );

    \I__17962\ : ClkMux
    port map (
            O => \N__73153\,
            I => \N__72833\
        );

    \I__17961\ : ClkMux
    port map (
            O => \N__73152\,
            I => \N__72833\
        );

    \I__17960\ : ClkMux
    port map (
            O => \N__73151\,
            I => \N__72833\
        );

    \I__17959\ : ClkMux
    port map (
            O => \N__73150\,
            I => \N__72833\
        );

    \I__17958\ : ClkMux
    port map (
            O => \N__73149\,
            I => \N__72833\
        );

    \I__17957\ : ClkMux
    port map (
            O => \N__73148\,
            I => \N__72833\
        );

    \I__17956\ : ClkMux
    port map (
            O => \N__73147\,
            I => \N__72833\
        );

    \I__17955\ : ClkMux
    port map (
            O => \N__73146\,
            I => \N__72833\
        );

    \I__17954\ : ClkMux
    port map (
            O => \N__73145\,
            I => \N__72833\
        );

    \I__17953\ : ClkMux
    port map (
            O => \N__73144\,
            I => \N__72833\
        );

    \I__17952\ : ClkMux
    port map (
            O => \N__73143\,
            I => \N__72833\
        );

    \I__17951\ : ClkMux
    port map (
            O => \N__73142\,
            I => \N__72833\
        );

    \I__17950\ : ClkMux
    port map (
            O => \N__73141\,
            I => \N__72833\
        );

    \I__17949\ : ClkMux
    port map (
            O => \N__73140\,
            I => \N__72833\
        );

    \I__17948\ : ClkMux
    port map (
            O => \N__73139\,
            I => \N__72833\
        );

    \I__17947\ : ClkMux
    port map (
            O => \N__73138\,
            I => \N__72833\
        );

    \I__17946\ : GlobalMux
    port map (
            O => \N__72833\,
            I => \N__72830\
        );

    \I__17945\ : gio2CtrlBuf
    port map (
            O => \N__72830\,
            I => \CLK_c_g\
        );

    \I__17944\ : InMux
    port map (
            O => \N__72827\,
            I => \N__72824\
        );

    \I__17943\ : LocalMux
    port map (
            O => \N__72824\,
            I => \N__72821\
        );

    \I__17942\ : Span4Mux_v
    port map (
            O => \N__72821\,
            I => \N__72818\
        );

    \I__17941\ : Odrv4
    port map (
            O => \N__72818\,
            I => \PROM.ROMDATA.m181\
        );

    \I__17940\ : InMux
    port map (
            O => \N__72815\,
            I => \N__72812\
        );

    \I__17939\ : LocalMux
    port map (
            O => \N__72812\,
            I => \PROM.ROMDATA.m480_bm\
        );

    \I__17938\ : CascadeMux
    port map (
            O => \N__72809\,
            I => \PROM.ROMDATA.m480_am_cascade_\
        );

    \I__17937\ : InMux
    port map (
            O => \N__72806\,
            I => \N__72803\
        );

    \I__17936\ : LocalMux
    port map (
            O => \N__72803\,
            I => \N__72800\
        );

    \I__17935\ : Span4Mux_h
    port map (
            O => \N__72800\,
            I => \N__72797\
        );

    \I__17934\ : Span4Mux_h
    port map (
            O => \N__72797\,
            I => \N__72794\
        );

    \I__17933\ : Odrv4
    port map (
            O => \N__72794\,
            I => \PROM.ROMDATA.N_551_mux\
        );

    \I__17932\ : CascadeMux
    port map (
            O => \N__72791\,
            I => \N__72786\
        );

    \I__17931\ : CascadeMux
    port map (
            O => \N__72790\,
            I => \N__72781\
        );

    \I__17930\ : CascadeMux
    port map (
            O => \N__72789\,
            I => \N__72778\
        );

    \I__17929\ : InMux
    port map (
            O => \N__72786\,
            I => \N__72761\
        );

    \I__17928\ : InMux
    port map (
            O => \N__72785\,
            I => \N__72761\
        );

    \I__17927\ : InMux
    port map (
            O => \N__72784\,
            I => \N__72761\
        );

    \I__17926\ : InMux
    port map (
            O => \N__72781\,
            I => \N__72752\
        );

    \I__17925\ : InMux
    port map (
            O => \N__72778\,
            I => \N__72752\
        );

    \I__17924\ : InMux
    port map (
            O => \N__72777\,
            I => \N__72752\
        );

    \I__17923\ : InMux
    port map (
            O => \N__72776\,
            I => \N__72752\
        );

    \I__17922\ : InMux
    port map (
            O => \N__72775\,
            I => \N__72749\
        );

    \I__17921\ : InMux
    port map (
            O => \N__72774\,
            I => \N__72746\
        );

    \I__17920\ : InMux
    port map (
            O => \N__72773\,
            I => \N__72743\
        );

    \I__17919\ : CascadeMux
    port map (
            O => \N__72772\,
            I => \N__72738\
        );

    \I__17918\ : InMux
    port map (
            O => \N__72771\,
            I => \N__72732\
        );

    \I__17917\ : InMux
    port map (
            O => \N__72770\,
            I => \N__72732\
        );

    \I__17916\ : CascadeMux
    port map (
            O => \N__72769\,
            I => \N__72717\
        );

    \I__17915\ : CascadeMux
    port map (
            O => \N__72768\,
            I => \N__72714\
        );

    \I__17914\ : LocalMux
    port map (
            O => \N__72761\,
            I => \N__72707\
        );

    \I__17913\ : LocalMux
    port map (
            O => \N__72752\,
            I => \N__72707\
        );

    \I__17912\ : LocalMux
    port map (
            O => \N__72749\,
            I => \N__72704\
        );

    \I__17911\ : LocalMux
    port map (
            O => \N__72746\,
            I => \N__72699\
        );

    \I__17910\ : LocalMux
    port map (
            O => \N__72743\,
            I => \N__72699\
        );

    \I__17909\ : CascadeMux
    port map (
            O => \N__72742\,
            I => \N__72685\
        );

    \I__17908\ : InMux
    port map (
            O => \N__72741\,
            I => \N__72676\
        );

    \I__17907\ : InMux
    port map (
            O => \N__72738\,
            I => \N__72676\
        );

    \I__17906\ : InMux
    port map (
            O => \N__72737\,
            I => \N__72673\
        );

    \I__17905\ : LocalMux
    port map (
            O => \N__72732\,
            I => \N__72669\
        );

    \I__17904\ : InMux
    port map (
            O => \N__72731\,
            I => \N__72666\
        );

    \I__17903\ : InMux
    port map (
            O => \N__72730\,
            I => \N__72657\
        );

    \I__17902\ : InMux
    port map (
            O => \N__72729\,
            I => \N__72657\
        );

    \I__17901\ : InMux
    port map (
            O => \N__72728\,
            I => \N__72657\
        );

    \I__17900\ : InMux
    port map (
            O => \N__72727\,
            I => \N__72657\
        );

    \I__17899\ : CascadeMux
    port map (
            O => \N__72726\,
            I => \N__72652\
        );

    \I__17898\ : CascadeMux
    port map (
            O => \N__72725\,
            I => \N__72649\
        );

    \I__17897\ : InMux
    port map (
            O => \N__72724\,
            I => \N__72637\
        );

    \I__17896\ : InMux
    port map (
            O => \N__72723\,
            I => \N__72637\
        );

    \I__17895\ : InMux
    port map (
            O => \N__72722\,
            I => \N__72637\
        );

    \I__17894\ : InMux
    port map (
            O => \N__72721\,
            I => \N__72637\
        );

    \I__17893\ : InMux
    port map (
            O => \N__72720\,
            I => \N__72637\
        );

    \I__17892\ : InMux
    port map (
            O => \N__72717\,
            I => \N__72630\
        );

    \I__17891\ : InMux
    port map (
            O => \N__72714\,
            I => \N__72630\
        );

    \I__17890\ : InMux
    port map (
            O => \N__72713\,
            I => \N__72630\
        );

    \I__17889\ : InMux
    port map (
            O => \N__72712\,
            I => \N__72627\
        );

    \I__17888\ : Span4Mux_v
    port map (
            O => \N__72707\,
            I => \N__72619\
        );

    \I__17887\ : Span4Mux_v
    port map (
            O => \N__72704\,
            I => \N__72619\
        );

    \I__17886\ : Span4Mux_v
    port map (
            O => \N__72699\,
            I => \N__72619\
        );

    \I__17885\ : CascadeMux
    port map (
            O => \N__72698\,
            I => \N__72615\
        );

    \I__17884\ : InMux
    port map (
            O => \N__72697\,
            I => \N__72612\
        );

    \I__17883\ : InMux
    port map (
            O => \N__72696\,
            I => \N__72609\
        );

    \I__17882\ : InMux
    port map (
            O => \N__72695\,
            I => \N__72603\
        );

    \I__17881\ : InMux
    port map (
            O => \N__72694\,
            I => \N__72600\
        );

    \I__17880\ : InMux
    port map (
            O => \N__72693\,
            I => \N__72597\
        );

    \I__17879\ : InMux
    port map (
            O => \N__72692\,
            I => \N__72588\
        );

    \I__17878\ : InMux
    port map (
            O => \N__72691\,
            I => \N__72588\
        );

    \I__17877\ : InMux
    port map (
            O => \N__72690\,
            I => \N__72588\
        );

    \I__17876\ : InMux
    port map (
            O => \N__72689\,
            I => \N__72588\
        );

    \I__17875\ : InMux
    port map (
            O => \N__72688\,
            I => \N__72583\
        );

    \I__17874\ : InMux
    port map (
            O => \N__72685\,
            I => \N__72583\
        );

    \I__17873\ : InMux
    port map (
            O => \N__72684\,
            I => \N__72580\
        );

    \I__17872\ : InMux
    port map (
            O => \N__72683\,
            I => \N__72577\
        );

    \I__17871\ : InMux
    port map (
            O => \N__72682\,
            I => \N__72572\
        );

    \I__17870\ : InMux
    port map (
            O => \N__72681\,
            I => \N__72572\
        );

    \I__17869\ : LocalMux
    port map (
            O => \N__72676\,
            I => \N__72567\
        );

    \I__17868\ : LocalMux
    port map (
            O => \N__72673\,
            I => \N__72567\
        );

    \I__17867\ : CascadeMux
    port map (
            O => \N__72672\,
            I => \N__72564\
        );

    \I__17866\ : Span4Mux_h
    port map (
            O => \N__72669\,
            I => \N__72560\
        );

    \I__17865\ : LocalMux
    port map (
            O => \N__72666\,
            I => \N__72557\
        );

    \I__17864\ : LocalMux
    port map (
            O => \N__72657\,
            I => \N__72554\
        );

    \I__17863\ : InMux
    port map (
            O => \N__72656\,
            I => \N__72549\
        );

    \I__17862\ : InMux
    port map (
            O => \N__72655\,
            I => \N__72549\
        );

    \I__17861\ : InMux
    port map (
            O => \N__72652\,
            I => \N__72546\
        );

    \I__17860\ : InMux
    port map (
            O => \N__72649\,
            I => \N__72541\
        );

    \I__17859\ : InMux
    port map (
            O => \N__72648\,
            I => \N__72541\
        );

    \I__17858\ : LocalMux
    port map (
            O => \N__72637\,
            I => \N__72538\
        );

    \I__17857\ : LocalMux
    port map (
            O => \N__72630\,
            I => \N__72535\
        );

    \I__17856\ : LocalMux
    port map (
            O => \N__72627\,
            I => \N__72532\
        );

    \I__17855\ : CascadeMux
    port map (
            O => \N__72626\,
            I => \N__72529\
        );

    \I__17854\ : Span4Mux_h
    port map (
            O => \N__72619\,
            I => \N__72526\
        );

    \I__17853\ : InMux
    port map (
            O => \N__72618\,
            I => \N__72523\
        );

    \I__17852\ : InMux
    port map (
            O => \N__72615\,
            I => \N__72520\
        );

    \I__17851\ : LocalMux
    port map (
            O => \N__72612\,
            I => \N__72515\
        );

    \I__17850\ : LocalMux
    port map (
            O => \N__72609\,
            I => \N__72515\
        );

    \I__17849\ : InMux
    port map (
            O => \N__72608\,
            I => \N__72512\
        );

    \I__17848\ : CascadeMux
    port map (
            O => \N__72607\,
            I => \N__72508\
        );

    \I__17847\ : CascadeMux
    port map (
            O => \N__72606\,
            I => \N__72505\
        );

    \I__17846\ : LocalMux
    port map (
            O => \N__72603\,
            I => \N__72500\
        );

    \I__17845\ : LocalMux
    port map (
            O => \N__72600\,
            I => \N__72495\
        );

    \I__17844\ : LocalMux
    port map (
            O => \N__72597\,
            I => \N__72495\
        );

    \I__17843\ : LocalMux
    port map (
            O => \N__72588\,
            I => \N__72490\
        );

    \I__17842\ : LocalMux
    port map (
            O => \N__72583\,
            I => \N__72490\
        );

    \I__17841\ : LocalMux
    port map (
            O => \N__72580\,
            I => \N__72485\
        );

    \I__17840\ : LocalMux
    port map (
            O => \N__72577\,
            I => \N__72485\
        );

    \I__17839\ : LocalMux
    port map (
            O => \N__72572\,
            I => \N__72480\
        );

    \I__17838\ : Span4Mux_v
    port map (
            O => \N__72567\,
            I => \N__72480\
        );

    \I__17837\ : InMux
    port map (
            O => \N__72564\,
            I => \N__72475\
        );

    \I__17836\ : InMux
    port map (
            O => \N__72563\,
            I => \N__72475\
        );

    \I__17835\ : Span4Mux_v
    port map (
            O => \N__72560\,
            I => \N__72470\
        );

    \I__17834\ : Span4Mux_v
    port map (
            O => \N__72557\,
            I => \N__72470\
        );

    \I__17833\ : Span4Mux_v
    port map (
            O => \N__72554\,
            I => \N__72461\
        );

    \I__17832\ : LocalMux
    port map (
            O => \N__72549\,
            I => \N__72461\
        );

    \I__17831\ : LocalMux
    port map (
            O => \N__72546\,
            I => \N__72461\
        );

    \I__17830\ : LocalMux
    port map (
            O => \N__72541\,
            I => \N__72461\
        );

    \I__17829\ : Span4Mux_v
    port map (
            O => \N__72538\,
            I => \N__72454\
        );

    \I__17828\ : Span4Mux_h
    port map (
            O => \N__72535\,
            I => \N__72454\
        );

    \I__17827\ : Span4Mux_h
    port map (
            O => \N__72532\,
            I => \N__72454\
        );

    \I__17826\ : InMux
    port map (
            O => \N__72529\,
            I => \N__72451\
        );

    \I__17825\ : Span4Mux_h
    port map (
            O => \N__72526\,
            I => \N__72446\
        );

    \I__17824\ : LocalMux
    port map (
            O => \N__72523\,
            I => \N__72446\
        );

    \I__17823\ : LocalMux
    port map (
            O => \N__72520\,
            I => \N__72439\
        );

    \I__17822\ : Span12Mux_h
    port map (
            O => \N__72515\,
            I => \N__72439\
        );

    \I__17821\ : LocalMux
    port map (
            O => \N__72512\,
            I => \N__72439\
        );

    \I__17820\ : InMux
    port map (
            O => \N__72511\,
            I => \N__72436\
        );

    \I__17819\ : InMux
    port map (
            O => \N__72508\,
            I => \N__72433\
        );

    \I__17818\ : InMux
    port map (
            O => \N__72505\,
            I => \N__72430\
        );

    \I__17817\ : InMux
    port map (
            O => \N__72504\,
            I => \N__72427\
        );

    \I__17816\ : InMux
    port map (
            O => \N__72503\,
            I => \N__72424\
        );

    \I__17815\ : Span4Mux_h
    port map (
            O => \N__72500\,
            I => \N__72415\
        );

    \I__17814\ : Span4Mux_v
    port map (
            O => \N__72495\,
            I => \N__72415\
        );

    \I__17813\ : Span4Mux_v
    port map (
            O => \N__72490\,
            I => \N__72415\
        );

    \I__17812\ : Span4Mux_h
    port map (
            O => \N__72485\,
            I => \N__72415\
        );

    \I__17811\ : Span4Mux_h
    port map (
            O => \N__72480\,
            I => \N__72404\
        );

    \I__17810\ : LocalMux
    port map (
            O => \N__72475\,
            I => \N__72404\
        );

    \I__17809\ : Span4Mux_h
    port map (
            O => \N__72470\,
            I => \N__72404\
        );

    \I__17808\ : Span4Mux_v
    port map (
            O => \N__72461\,
            I => \N__72404\
        );

    \I__17807\ : Span4Mux_v
    port map (
            O => \N__72454\,
            I => \N__72404\
        );

    \I__17806\ : LocalMux
    port map (
            O => \N__72451\,
            I => \progRomAddress_7\
        );

    \I__17805\ : Odrv4
    port map (
            O => \N__72446\,
            I => \progRomAddress_7\
        );

    \I__17804\ : Odrv12
    port map (
            O => \N__72439\,
            I => \progRomAddress_7\
        );

    \I__17803\ : LocalMux
    port map (
            O => \N__72436\,
            I => \progRomAddress_7\
        );

    \I__17802\ : LocalMux
    port map (
            O => \N__72433\,
            I => \progRomAddress_7\
        );

    \I__17801\ : LocalMux
    port map (
            O => \N__72430\,
            I => \progRomAddress_7\
        );

    \I__17800\ : LocalMux
    port map (
            O => \N__72427\,
            I => \progRomAddress_7\
        );

    \I__17799\ : LocalMux
    port map (
            O => \N__72424\,
            I => \progRomAddress_7\
        );

    \I__17798\ : Odrv4
    port map (
            O => \N__72415\,
            I => \progRomAddress_7\
        );

    \I__17797\ : Odrv4
    port map (
            O => \N__72404\,
            I => \progRomAddress_7\
        );

    \I__17796\ : CascadeMux
    port map (
            O => \N__72383\,
            I => \PROM.ROMDATA.m480_ns_cascade_\
        );

    \I__17795\ : InMux
    port map (
            O => \N__72380\,
            I => \N__72377\
        );

    \I__17794\ : LocalMux
    port map (
            O => \N__72377\,
            I => \N__72373\
        );

    \I__17793\ : InMux
    port map (
            O => \N__72376\,
            I => \N__72370\
        );

    \I__17792\ : Span4Mux_h
    port map (
            O => \N__72373\,
            I => \N__72367\
        );

    \I__17791\ : LocalMux
    port map (
            O => \N__72370\,
            I => \N__72364\
        );

    \I__17790\ : Span4Mux_h
    port map (
            O => \N__72367\,
            I => \N__72361\
        );

    \I__17789\ : Span12Mux_h
    port map (
            O => \N__72364\,
            I => \N__72358\
        );

    \I__17788\ : Odrv4
    port map (
            O => \N__72361\,
            I => \PROM_ROMDATA_dintern_25ro\
        );

    \I__17787\ : Odrv12
    port map (
            O => \N__72358\,
            I => \PROM_ROMDATA_dintern_25ro\
        );

    \I__17786\ : InMux
    port map (
            O => \N__72353\,
            I => \N__72349\
        );

    \I__17785\ : InMux
    port map (
            O => \N__72352\,
            I => \N__72345\
        );

    \I__17784\ : LocalMux
    port map (
            O => \N__72349\,
            I => \N__72342\
        );

    \I__17783\ : InMux
    port map (
            O => \N__72348\,
            I => \N__72339\
        );

    \I__17782\ : LocalMux
    port map (
            O => \N__72345\,
            I => \N__72336\
        );

    \I__17781\ : Span4Mux_h
    port map (
            O => \N__72342\,
            I => \N__72331\
        );

    \I__17780\ : LocalMux
    port map (
            O => \N__72339\,
            I => \N__72331\
        );

    \I__17779\ : Span4Mux_h
    port map (
            O => \N__72336\,
            I => \N__72328\
        );

    \I__17778\ : Span4Mux_h
    port map (
            O => \N__72331\,
            I => \N__72325\
        );

    \I__17777\ : Odrv4
    port map (
            O => \N__72328\,
            I => g_9
        );

    \I__17776\ : Odrv4
    port map (
            O => \N__72325\,
            I => g_9
        );

    \I__17775\ : CascadeMux
    port map (
            O => \N__72320\,
            I => \N__72312\
        );

    \I__17774\ : CascadeMux
    port map (
            O => \N__72319\,
            I => \N__72308\
        );

    \I__17773\ : InMux
    port map (
            O => \N__72318\,
            I => \N__72301\
        );

    \I__17772\ : CascadeMux
    port map (
            O => \N__72317\,
            I => \N__72294\
        );

    \I__17771\ : CascadeMux
    port map (
            O => \N__72316\,
            I => \N__72290\
        );

    \I__17770\ : CascadeMux
    port map (
            O => \N__72315\,
            I => \N__72285\
        );

    \I__17769\ : InMux
    port map (
            O => \N__72312\,
            I => \N__72281\
        );

    \I__17768\ : InMux
    port map (
            O => \N__72311\,
            I => \N__72274\
        );

    \I__17767\ : InMux
    port map (
            O => \N__72308\,
            I => \N__72274\
        );

    \I__17766\ : InMux
    port map (
            O => \N__72307\,
            I => \N__72274\
        );

    \I__17765\ : CascadeMux
    port map (
            O => \N__72306\,
            I => \N__72268\
        );

    \I__17764\ : CascadeMux
    port map (
            O => \N__72305\,
            I => \N__72265\
        );

    \I__17763\ : InMux
    port map (
            O => \N__72304\,
            I => \N__72257\
        );

    \I__17762\ : LocalMux
    port map (
            O => \N__72301\,
            I => \N__72253\
        );

    \I__17761\ : InMux
    port map (
            O => \N__72300\,
            I => \N__72244\
        );

    \I__17760\ : InMux
    port map (
            O => \N__72299\,
            I => \N__72239\
        );

    \I__17759\ : InMux
    port map (
            O => \N__72298\,
            I => \N__72239\
        );

    \I__17758\ : InMux
    port map (
            O => \N__72297\,
            I => \N__72236\
        );

    \I__17757\ : InMux
    port map (
            O => \N__72294\,
            I => \N__72231\
        );

    \I__17756\ : InMux
    port map (
            O => \N__72293\,
            I => \N__72231\
        );

    \I__17755\ : InMux
    port map (
            O => \N__72290\,
            I => \N__72228\
        );

    \I__17754\ : CascadeMux
    port map (
            O => \N__72289\,
            I => \N__72217\
        );

    \I__17753\ : CascadeMux
    port map (
            O => \N__72288\,
            I => \N__72214\
        );

    \I__17752\ : InMux
    port map (
            O => \N__72285\,
            I => \N__72209\
        );

    \I__17751\ : CascadeMux
    port map (
            O => \N__72284\,
            I => \N__72206\
        );

    \I__17750\ : LocalMux
    port map (
            O => \N__72281\,
            I => \N__72201\
        );

    \I__17749\ : LocalMux
    port map (
            O => \N__72274\,
            I => \N__72201\
        );

    \I__17748\ : InMux
    port map (
            O => \N__72273\,
            I => \N__72198\
        );

    \I__17747\ : InMux
    port map (
            O => \N__72272\,
            I => \N__72195\
        );

    \I__17746\ : InMux
    port map (
            O => \N__72271\,
            I => \N__72185\
        );

    \I__17745\ : InMux
    port map (
            O => \N__72268\,
            I => \N__72182\
        );

    \I__17744\ : InMux
    port map (
            O => \N__72265\,
            I => \N__72171\
        );

    \I__17743\ : InMux
    port map (
            O => \N__72264\,
            I => \N__72171\
        );

    \I__17742\ : InMux
    port map (
            O => \N__72263\,
            I => \N__72166\
        );

    \I__17741\ : InMux
    port map (
            O => \N__72262\,
            I => \N__72166\
        );

    \I__17740\ : InMux
    port map (
            O => \N__72261\,
            I => \N__72161\
        );

    \I__17739\ : InMux
    port map (
            O => \N__72260\,
            I => \N__72161\
        );

    \I__17738\ : LocalMux
    port map (
            O => \N__72257\,
            I => \N__72158\
        );

    \I__17737\ : InMux
    port map (
            O => \N__72256\,
            I => \N__72155\
        );

    \I__17736\ : Span4Mux_h
    port map (
            O => \N__72253\,
            I => \N__72152\
        );

    \I__17735\ : InMux
    port map (
            O => \N__72252\,
            I => \N__72149\
        );

    \I__17734\ : InMux
    port map (
            O => \N__72251\,
            I => \N__72146\
        );

    \I__17733\ : InMux
    port map (
            O => \N__72250\,
            I => \N__72141\
        );

    \I__17732\ : InMux
    port map (
            O => \N__72249\,
            I => \N__72141\
        );

    \I__17731\ : InMux
    port map (
            O => \N__72248\,
            I => \N__72137\
        );

    \I__17730\ : InMux
    port map (
            O => \N__72247\,
            I => \N__72134\
        );

    \I__17729\ : LocalMux
    port map (
            O => \N__72244\,
            I => \N__72123\
        );

    \I__17728\ : LocalMux
    port map (
            O => \N__72239\,
            I => \N__72123\
        );

    \I__17727\ : LocalMux
    port map (
            O => \N__72236\,
            I => \N__72118\
        );

    \I__17726\ : LocalMux
    port map (
            O => \N__72231\,
            I => \N__72118\
        );

    \I__17725\ : LocalMux
    port map (
            O => \N__72228\,
            I => \N__72115\
        );

    \I__17724\ : InMux
    port map (
            O => \N__72227\,
            I => \N__72110\
        );

    \I__17723\ : InMux
    port map (
            O => \N__72226\,
            I => \N__72110\
        );

    \I__17722\ : InMux
    port map (
            O => \N__72225\,
            I => \N__72105\
        );

    \I__17721\ : InMux
    port map (
            O => \N__72224\,
            I => \N__72105\
        );

    \I__17720\ : InMux
    port map (
            O => \N__72223\,
            I => \N__72097\
        );

    \I__17719\ : InMux
    port map (
            O => \N__72222\,
            I => \N__72092\
        );

    \I__17718\ : InMux
    port map (
            O => \N__72221\,
            I => \N__72092\
        );

    \I__17717\ : InMux
    port map (
            O => \N__72220\,
            I => \N__72081\
        );

    \I__17716\ : InMux
    port map (
            O => \N__72217\,
            I => \N__72081\
        );

    \I__17715\ : InMux
    port map (
            O => \N__72214\,
            I => \N__72081\
        );

    \I__17714\ : InMux
    port map (
            O => \N__72213\,
            I => \N__72081\
        );

    \I__17713\ : InMux
    port map (
            O => \N__72212\,
            I => \N__72081\
        );

    \I__17712\ : LocalMux
    port map (
            O => \N__72209\,
            I => \N__72078\
        );

    \I__17711\ : InMux
    port map (
            O => \N__72206\,
            I => \N__72075\
        );

    \I__17710\ : Span4Mux_v
    port map (
            O => \N__72201\,
            I => \N__72068\
        );

    \I__17709\ : LocalMux
    port map (
            O => \N__72198\,
            I => \N__72068\
        );

    \I__17708\ : LocalMux
    port map (
            O => \N__72195\,
            I => \N__72068\
        );

    \I__17707\ : InMux
    port map (
            O => \N__72194\,
            I => \N__72061\
        );

    \I__17706\ : InMux
    port map (
            O => \N__72193\,
            I => \N__72061\
        );

    \I__17705\ : InMux
    port map (
            O => \N__72192\,
            I => \N__72061\
        );

    \I__17704\ : InMux
    port map (
            O => \N__72191\,
            I => \N__72052\
        );

    \I__17703\ : InMux
    port map (
            O => \N__72190\,
            I => \N__72052\
        );

    \I__17702\ : InMux
    port map (
            O => \N__72189\,
            I => \N__72052\
        );

    \I__17701\ : InMux
    port map (
            O => \N__72188\,
            I => \N__72052\
        );

    \I__17700\ : LocalMux
    port map (
            O => \N__72185\,
            I => \N__72047\
        );

    \I__17699\ : LocalMux
    port map (
            O => \N__72182\,
            I => \N__72047\
        );

    \I__17698\ : InMux
    port map (
            O => \N__72181\,
            I => \N__72044\
        );

    \I__17697\ : InMux
    port map (
            O => \N__72180\,
            I => \N__72033\
        );

    \I__17696\ : InMux
    port map (
            O => \N__72179\,
            I => \N__72033\
        );

    \I__17695\ : InMux
    port map (
            O => \N__72178\,
            I => \N__72033\
        );

    \I__17694\ : InMux
    port map (
            O => \N__72177\,
            I => \N__72033\
        );

    \I__17693\ : InMux
    port map (
            O => \N__72176\,
            I => \N__72033\
        );

    \I__17692\ : LocalMux
    port map (
            O => \N__72171\,
            I => \N__72026\
        );

    \I__17691\ : LocalMux
    port map (
            O => \N__72166\,
            I => \N__72026\
        );

    \I__17690\ : LocalMux
    port map (
            O => \N__72161\,
            I => \N__72026\
        );

    \I__17689\ : Span4Mux_h
    port map (
            O => \N__72158\,
            I => \N__72013\
        );

    \I__17688\ : LocalMux
    port map (
            O => \N__72155\,
            I => \N__72013\
        );

    \I__17687\ : Span4Mux_h
    port map (
            O => \N__72152\,
            I => \N__72013\
        );

    \I__17686\ : LocalMux
    port map (
            O => \N__72149\,
            I => \N__72013\
        );

    \I__17685\ : LocalMux
    port map (
            O => \N__72146\,
            I => \N__72013\
        );

    \I__17684\ : LocalMux
    port map (
            O => \N__72141\,
            I => \N__72013\
        );

    \I__17683\ : CascadeMux
    port map (
            O => \N__72140\,
            I => \N__72010\
        );

    \I__17682\ : LocalMux
    port map (
            O => \N__72137\,
            I => \N__72005\
        );

    \I__17681\ : LocalMux
    port map (
            O => \N__72134\,
            I => \N__72002\
        );

    \I__17680\ : InMux
    port map (
            O => \N__72133\,
            I => \N__71997\
        );

    \I__17679\ : InMux
    port map (
            O => \N__72132\,
            I => \N__71997\
        );

    \I__17678\ : InMux
    port map (
            O => \N__72131\,
            I => \N__71994\
        );

    \I__17677\ : InMux
    port map (
            O => \N__72130\,
            I => \N__71987\
        );

    \I__17676\ : InMux
    port map (
            O => \N__72129\,
            I => \N__71987\
        );

    \I__17675\ : InMux
    port map (
            O => \N__72128\,
            I => \N__71987\
        );

    \I__17674\ : Span12Mux_h
    port map (
            O => \N__72123\,
            I => \N__71976\
        );

    \I__17673\ : Sp12to4
    port map (
            O => \N__72118\,
            I => \N__71976\
        );

    \I__17672\ : Sp12to4
    port map (
            O => \N__72115\,
            I => \N__71976\
        );

    \I__17671\ : LocalMux
    port map (
            O => \N__72110\,
            I => \N__71976\
        );

    \I__17670\ : LocalMux
    port map (
            O => \N__72105\,
            I => \N__71976\
        );

    \I__17669\ : InMux
    port map (
            O => \N__72104\,
            I => \N__71973\
        );

    \I__17668\ : InMux
    port map (
            O => \N__72103\,
            I => \N__71968\
        );

    \I__17667\ : InMux
    port map (
            O => \N__72102\,
            I => \N__71968\
        );

    \I__17666\ : InMux
    port map (
            O => \N__72101\,
            I => \N__71963\
        );

    \I__17665\ : InMux
    port map (
            O => \N__72100\,
            I => \N__71963\
        );

    \I__17664\ : LocalMux
    port map (
            O => \N__72097\,
            I => \N__71960\
        );

    \I__17663\ : LocalMux
    port map (
            O => \N__72092\,
            I => \N__71951\
        );

    \I__17662\ : LocalMux
    port map (
            O => \N__72081\,
            I => \N__71951\
        );

    \I__17661\ : Span4Mux_h
    port map (
            O => \N__72078\,
            I => \N__71951\
        );

    \I__17660\ : LocalMux
    port map (
            O => \N__72075\,
            I => \N__71951\
        );

    \I__17659\ : Span4Mux_v
    port map (
            O => \N__72068\,
            I => \N__71948\
        );

    \I__17658\ : LocalMux
    port map (
            O => \N__72061\,
            I => \N__71935\
        );

    \I__17657\ : LocalMux
    port map (
            O => \N__72052\,
            I => \N__71935\
        );

    \I__17656\ : Span4Mux_v
    port map (
            O => \N__72047\,
            I => \N__71935\
        );

    \I__17655\ : LocalMux
    port map (
            O => \N__72044\,
            I => \N__71935\
        );

    \I__17654\ : LocalMux
    port map (
            O => \N__72033\,
            I => \N__71935\
        );

    \I__17653\ : Span4Mux_h
    port map (
            O => \N__72026\,
            I => \N__71935\
        );

    \I__17652\ : Span4Mux_h
    port map (
            O => \N__72013\,
            I => \N__71932\
        );

    \I__17651\ : InMux
    port map (
            O => \N__72010\,
            I => \N__71925\
        );

    \I__17650\ : InMux
    port map (
            O => \N__72009\,
            I => \N__71925\
        );

    \I__17649\ : InMux
    port map (
            O => \N__72008\,
            I => \N__71925\
        );

    \I__17648\ : Span4Mux_v
    port map (
            O => \N__72005\,
            I => \N__71922\
        );

    \I__17647\ : Span4Mux_h
    port map (
            O => \N__72002\,
            I => \N__71915\
        );

    \I__17646\ : LocalMux
    port map (
            O => \N__71997\,
            I => \N__71915\
        );

    \I__17645\ : LocalMux
    port map (
            O => \N__71994\,
            I => \N__71915\
        );

    \I__17644\ : LocalMux
    port map (
            O => \N__71987\,
            I => \N__71910\
        );

    \I__17643\ : Span12Mux_v
    port map (
            O => \N__71976\,
            I => \N__71910\
        );

    \I__17642\ : LocalMux
    port map (
            O => \N__71973\,
            I => \N__71895\
        );

    \I__17641\ : LocalMux
    port map (
            O => \N__71968\,
            I => \N__71895\
        );

    \I__17640\ : LocalMux
    port map (
            O => \N__71963\,
            I => \N__71895\
        );

    \I__17639\ : Span4Mux_v
    port map (
            O => \N__71960\,
            I => \N__71895\
        );

    \I__17638\ : Span4Mux_v
    port map (
            O => \N__71951\,
            I => \N__71895\
        );

    \I__17637\ : Span4Mux_h
    port map (
            O => \N__71948\,
            I => \N__71895\
        );

    \I__17636\ : Span4Mux_v
    port map (
            O => \N__71935\,
            I => \N__71895\
        );

    \I__17635\ : Span4Mux_h
    port map (
            O => \N__71932\,
            I => \N__71892\
        );

    \I__17634\ : LocalMux
    port map (
            O => \N__71925\,
            I => \PROM_ROMDATA_dintern_adflt\
        );

    \I__17633\ : Odrv4
    port map (
            O => \N__71922\,
            I => \PROM_ROMDATA_dintern_adflt\
        );

    \I__17632\ : Odrv4
    port map (
            O => \N__71915\,
            I => \PROM_ROMDATA_dintern_adflt\
        );

    \I__17631\ : Odrv12
    port map (
            O => \N__71910\,
            I => \PROM_ROMDATA_dintern_adflt\
        );

    \I__17630\ : Odrv4
    port map (
            O => \N__71895\,
            I => \PROM_ROMDATA_dintern_adflt\
        );

    \I__17629\ : Odrv4
    port map (
            O => \N__71892\,
            I => \PROM_ROMDATA_dintern_adflt\
        );

    \I__17628\ : CascadeMux
    port map (
            O => \N__71879\,
            I => \PROM_ROMDATA_dintern_25ro_cascade_\
        );

    \I__17627\ : CascadeMux
    port map (
            O => \N__71876\,
            I => \N__71863\
        );

    \I__17626\ : InMux
    port map (
            O => \N__71875\,
            I => \N__71860\
        );

    \I__17625\ : InMux
    port map (
            O => \N__71874\,
            I => \N__71855\
        );

    \I__17624\ : InMux
    port map (
            O => \N__71873\,
            I => \N__71855\
        );

    \I__17623\ : InMux
    port map (
            O => \N__71872\,
            I => \N__71849\
        );

    \I__17622\ : InMux
    port map (
            O => \N__71871\,
            I => \N__71842\
        );

    \I__17621\ : InMux
    port map (
            O => \N__71870\,
            I => \N__71842\
        );

    \I__17620\ : InMux
    port map (
            O => \N__71869\,
            I => \N__71842\
        );

    \I__17619\ : InMux
    port map (
            O => \N__71868\,
            I => \N__71835\
        );

    \I__17618\ : InMux
    port map (
            O => \N__71867\,
            I => \N__71835\
        );

    \I__17617\ : InMux
    port map (
            O => \N__71866\,
            I => \N__71835\
        );

    \I__17616\ : InMux
    port map (
            O => \N__71863\,
            I => \N__71832\
        );

    \I__17615\ : LocalMux
    port map (
            O => \N__71860\,
            I => \N__71816\
        );

    \I__17614\ : LocalMux
    port map (
            O => \N__71855\,
            I => \N__71813\
        );

    \I__17613\ : InMux
    port map (
            O => \N__71854\,
            I => \N__71810\
        );

    \I__17612\ : CascadeMux
    port map (
            O => \N__71853\,
            I => \N__71807\
        );

    \I__17611\ : CascadeMux
    port map (
            O => \N__71852\,
            I => \N__71799\
        );

    \I__17610\ : LocalMux
    port map (
            O => \N__71849\,
            I => \N__71792\
        );

    \I__17609\ : LocalMux
    port map (
            O => \N__71842\,
            I => \N__71792\
        );

    \I__17608\ : LocalMux
    port map (
            O => \N__71835\,
            I => \N__71792\
        );

    \I__17607\ : LocalMux
    port map (
            O => \N__71832\,
            I => \N__71789\
        );

    \I__17606\ : InMux
    port map (
            O => \N__71831\,
            I => \N__71786\
        );

    \I__17605\ : InMux
    port map (
            O => \N__71830\,
            I => \N__71783\
        );

    \I__17604\ : InMux
    port map (
            O => \N__71829\,
            I => \N__71776\
        );

    \I__17603\ : InMux
    port map (
            O => \N__71828\,
            I => \N__71776\
        );

    \I__17602\ : InMux
    port map (
            O => \N__71827\,
            I => \N__71776\
        );

    \I__17601\ : InMux
    port map (
            O => \N__71826\,
            I => \N__71765\
        );

    \I__17600\ : InMux
    port map (
            O => \N__71825\,
            I => \N__71765\
        );

    \I__17599\ : InMux
    port map (
            O => \N__71824\,
            I => \N__71765\
        );

    \I__17598\ : InMux
    port map (
            O => \N__71823\,
            I => \N__71765\
        );

    \I__17597\ : InMux
    port map (
            O => \N__71822\,
            I => \N__71765\
        );

    \I__17596\ : CascadeMux
    port map (
            O => \N__71821\,
            I => \N__71762\
        );

    \I__17595\ : InMux
    port map (
            O => \N__71820\,
            I => \N__71759\
        );

    \I__17594\ : CascadeMux
    port map (
            O => \N__71819\,
            I => \N__71755\
        );

    \I__17593\ : Span4Mux_h
    port map (
            O => \N__71816\,
            I => \N__71752\
        );

    \I__17592\ : Span4Mux_v
    port map (
            O => \N__71813\,
            I => \N__71749\
        );

    \I__17591\ : LocalMux
    port map (
            O => \N__71810\,
            I => \N__71746\
        );

    \I__17590\ : InMux
    port map (
            O => \N__71807\,
            I => \N__71742\
        );

    \I__17589\ : InMux
    port map (
            O => \N__71806\,
            I => \N__71739\
        );

    \I__17588\ : InMux
    port map (
            O => \N__71805\,
            I => \N__71730\
        );

    \I__17587\ : InMux
    port map (
            O => \N__71804\,
            I => \N__71730\
        );

    \I__17586\ : InMux
    port map (
            O => \N__71803\,
            I => \N__71730\
        );

    \I__17585\ : InMux
    port map (
            O => \N__71802\,
            I => \N__71730\
        );

    \I__17584\ : InMux
    port map (
            O => \N__71799\,
            I => \N__71727\
        );

    \I__17583\ : Span4Mux_v
    port map (
            O => \N__71792\,
            I => \N__71722\
        );

    \I__17582\ : Span4Mux_v
    port map (
            O => \N__71789\,
            I => \N__71722\
        );

    \I__17581\ : LocalMux
    port map (
            O => \N__71786\,
            I => \N__71715\
        );

    \I__17580\ : LocalMux
    port map (
            O => \N__71783\,
            I => \N__71715\
        );

    \I__17579\ : LocalMux
    port map (
            O => \N__71776\,
            I => \N__71715\
        );

    \I__17578\ : LocalMux
    port map (
            O => \N__71765\,
            I => \N__71712\
        );

    \I__17577\ : InMux
    port map (
            O => \N__71762\,
            I => \N__71709\
        );

    \I__17576\ : LocalMux
    port map (
            O => \N__71759\,
            I => \N__71706\
        );

    \I__17575\ : InMux
    port map (
            O => \N__71758\,
            I => \N__71701\
        );

    \I__17574\ : InMux
    port map (
            O => \N__71755\,
            I => \N__71701\
        );

    \I__17573\ : Span4Mux_h
    port map (
            O => \N__71752\,
            I => \N__71698\
        );

    \I__17572\ : Span4Mux_h
    port map (
            O => \N__71749\,
            I => \N__71693\
        );

    \I__17571\ : Span4Mux_v
    port map (
            O => \N__71746\,
            I => \N__71693\
        );

    \I__17570\ : InMux
    port map (
            O => \N__71745\,
            I => \N__71690\
        );

    \I__17569\ : LocalMux
    port map (
            O => \N__71742\,
            I => \N__71683\
        );

    \I__17568\ : LocalMux
    port map (
            O => \N__71739\,
            I => \N__71683\
        );

    \I__17567\ : LocalMux
    port map (
            O => \N__71730\,
            I => \N__71683\
        );

    \I__17566\ : LocalMux
    port map (
            O => \N__71727\,
            I => \N__71676\
        );

    \I__17565\ : Span4Mux_h
    port map (
            O => \N__71722\,
            I => \N__71676\
        );

    \I__17564\ : Span4Mux_v
    port map (
            O => \N__71715\,
            I => \N__71676\
        );

    \I__17563\ : Odrv12
    port map (
            O => \N__71712\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17562\ : LocalMux
    port map (
            O => \N__71709\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17561\ : Odrv4
    port map (
            O => \N__71706\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17560\ : LocalMux
    port map (
            O => \N__71701\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17559\ : Odrv4
    port map (
            O => \N__71698\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17558\ : Odrv4
    port map (
            O => \N__71693\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17557\ : LocalMux
    port map (
            O => \N__71690\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17556\ : Odrv4
    port map (
            O => \N__71683\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17555\ : Odrv4
    port map (
            O => \N__71676\,
            I => \PROM_ROMDATA_dintern_3ro\
        );

    \I__17554\ : CascadeMux
    port map (
            O => \N__71657\,
            I => \N__71654\
        );

    \I__17553\ : CascadeBuf
    port map (
            O => \N__71654\,
            I => \N__71651\
        );

    \I__17552\ : CascadeMux
    port map (
            O => \N__71651\,
            I => \N__71648\
        );

    \I__17551\ : CascadeBuf
    port map (
            O => \N__71648\,
            I => \N__71645\
        );

    \I__17550\ : CascadeMux
    port map (
            O => \N__71645\,
            I => \N__71642\
        );

    \I__17549\ : CascadeBuf
    port map (
            O => \N__71642\,
            I => \N__71639\
        );

    \I__17548\ : CascadeMux
    port map (
            O => \N__71639\,
            I => \N__71636\
        );

    \I__17547\ : InMux
    port map (
            O => \N__71636\,
            I => \N__71633\
        );

    \I__17546\ : LocalMux
    port map (
            O => \N__71633\,
            I => \N__71630\
        );

    \I__17545\ : Span4Mux_v
    port map (
            O => \N__71630\,
            I => \N__71627\
        );

    \I__17544\ : Sp12to4
    port map (
            O => \N__71627\,
            I => \N__71624\
        );

    \I__17543\ : Span12Mux_v
    port map (
            O => \N__71624\,
            I => \N__71621\
        );

    \I__17542\ : Span12Mux_h
    port map (
            O => \N__71621\,
            I => \N__71618\
        );

    \I__17541\ : Odrv12
    port map (
            O => \N__71618\,
            I => \CONTROL_romAddReg_7_9\
        );

    \I__17540\ : InMux
    port map (
            O => \N__71615\,
            I => \N__71612\
        );

    \I__17539\ : LocalMux
    port map (
            O => \N__71612\,
            I => \N__71609\
        );

    \I__17538\ : Span4Mux_h
    port map (
            O => \N__71609\,
            I => \N__71606\
        );

    \I__17537\ : Odrv4
    port map (
            O => \N__71606\,
            I => \PROM.ROMDATA.m446_bm\
        );

    \I__17536\ : InMux
    port map (
            O => \N__71603\,
            I => \N__71600\
        );

    \I__17535\ : LocalMux
    port map (
            O => \N__71600\,
            I => \N__71597\
        );

    \I__17534\ : Span4Mux_h
    port map (
            O => \N__71597\,
            I => \N__71594\
        );

    \I__17533\ : Span4Mux_h
    port map (
            O => \N__71594\,
            I => \N__71591\
        );

    \I__17532\ : Odrv4
    port map (
            O => \N__71591\,
            I => \PROM.ROMDATA.m447_ns_1\
        );

    \I__17531\ : CascadeMux
    port map (
            O => \N__71588\,
            I => \N__71585\
        );

    \I__17530\ : InMux
    port map (
            O => \N__71585\,
            I => \N__71582\
        );

    \I__17529\ : LocalMux
    port map (
            O => \N__71582\,
            I => \PROM.ROMDATA.m446_am\
        );

    \I__17528\ : InMux
    port map (
            O => \N__71579\,
            I => \N__71573\
        );

    \I__17527\ : InMux
    port map (
            O => \N__71578\,
            I => \N__71573\
        );

    \I__17526\ : LocalMux
    port map (
            O => \N__71573\,
            I => \N__71570\
        );

    \I__17525\ : Span4Mux_v
    port map (
            O => \N__71570\,
            I => \N__71567\
        );

    \I__17524\ : Sp12to4
    port map (
            O => \N__71567\,
            I => \N__71564\
        );

    \I__17523\ : Span12Mux_h
    port map (
            O => \N__71564\,
            I => \N__71561\
        );

    \I__17522\ : Odrv12
    port map (
            O => \N__71561\,
            I => \PROM.ROMDATA.m447_ns\
        );

    \I__17521\ : CEMux
    port map (
            O => \N__71558\,
            I => \N__71555\
        );

    \I__17520\ : LocalMux
    port map (
            O => \N__71555\,
            I => \N__71550\
        );

    \I__17519\ : CEMux
    port map (
            O => \N__71554\,
            I => \N__71547\
        );

    \I__17518\ : CEMux
    port map (
            O => \N__71553\,
            I => \N__71544\
        );

    \I__17517\ : Span4Mux_h
    port map (
            O => \N__71550\,
            I => \N__71539\
        );

    \I__17516\ : LocalMux
    port map (
            O => \N__71547\,
            I => \N__71539\
        );

    \I__17515\ : LocalMux
    port map (
            O => \N__71544\,
            I => \N__71536\
        );

    \I__17514\ : Span4Mux_h
    port map (
            O => \N__71539\,
            I => \N__71533\
        );

    \I__17513\ : Span4Mux_v
    port map (
            O => \N__71536\,
            I => \N__71530\
        );

    \I__17512\ : Span4Mux_h
    port map (
            O => \N__71533\,
            I => \N__71527\
        );

    \I__17511\ : Span4Mux_h
    port map (
            O => \N__71530\,
            I => \N__71522\
        );

    \I__17510\ : Span4Mux_h
    port map (
            O => \N__71527\,
            I => \N__71522\
        );

    \I__17509\ : Odrv4
    port map (
            O => \N__71522\,
            I => \ALU.un1_a41_7_0\
        );

    \I__17508\ : InMux
    port map (
            O => \N__71519\,
            I => \N__71516\
        );

    \I__17507\ : LocalMux
    port map (
            O => \N__71516\,
            I => \N__71512\
        );

    \I__17506\ : InMux
    port map (
            O => \N__71515\,
            I => \N__71509\
        );

    \I__17505\ : Odrv4
    port map (
            O => \N__71512\,
            I => \ALU.un1_operation_13Z0Z_2\
        );

    \I__17504\ : LocalMux
    port map (
            O => \N__71509\,
            I => \ALU.un1_operation_13Z0Z_2\
        );

    \I__17503\ : CascadeMux
    port map (
            O => \N__71504\,
            I => \N__71501\
        );

    \I__17502\ : InMux
    port map (
            O => \N__71501\,
            I => \N__71495\
        );

    \I__17501\ : InMux
    port map (
            O => \N__71500\,
            I => \N__71495\
        );

    \I__17500\ : LocalMux
    port map (
            O => \N__71495\,
            I => \N__71492\
        );

    \I__17499\ : Sp12to4
    port map (
            O => \N__71492\,
            I => \N__71487\
        );

    \I__17498\ : InMux
    port map (
            O => \N__71491\,
            I => \N__71484\
        );

    \I__17497\ : InMux
    port map (
            O => \N__71490\,
            I => \N__71481\
        );

    \I__17496\ : Span12Mux_v
    port map (
            O => \N__71487\,
            I => \N__71478\
        );

    \I__17495\ : LocalMux
    port map (
            O => \N__71484\,
            I => \ALU.un1_operation_10_0\
        );

    \I__17494\ : LocalMux
    port map (
            O => \N__71481\,
            I => \ALU.un1_operation_10_0\
        );

    \I__17493\ : Odrv12
    port map (
            O => \N__71478\,
            I => \ALU.un1_operation_10_0\
        );

    \I__17492\ : InMux
    port map (
            O => \N__71471\,
            I => \N__71464\
        );

    \I__17491\ : InMux
    port map (
            O => \N__71470\,
            I => \N__71460\
        );

    \I__17490\ : InMux
    port map (
            O => \N__71469\,
            I => \N__71455\
        );

    \I__17489\ : InMux
    port map (
            O => \N__71468\,
            I => \N__71455\
        );

    \I__17488\ : InMux
    port map (
            O => \N__71467\,
            I => \N__71445\
        );

    \I__17487\ : LocalMux
    port map (
            O => \N__71464\,
            I => \N__71442\
        );

    \I__17486\ : InMux
    port map (
            O => \N__71463\,
            I => \N__71437\
        );

    \I__17485\ : LocalMux
    port map (
            O => \N__71460\,
            I => \N__71432\
        );

    \I__17484\ : LocalMux
    port map (
            O => \N__71455\,
            I => \N__71429\
        );

    \I__17483\ : InMux
    port map (
            O => \N__71454\,
            I => \N__71426\
        );

    \I__17482\ : InMux
    port map (
            O => \N__71453\,
            I => \N__71418\
        );

    \I__17481\ : InMux
    port map (
            O => \N__71452\,
            I => \N__71418\
        );

    \I__17480\ : InMux
    port map (
            O => \N__71451\,
            I => \N__71411\
        );

    \I__17479\ : InMux
    port map (
            O => \N__71450\,
            I => \N__71411\
        );

    \I__17478\ : InMux
    port map (
            O => \N__71449\,
            I => \N__71411\
        );

    \I__17477\ : CascadeMux
    port map (
            O => \N__71448\,
            I => \N__71407\
        );

    \I__17476\ : LocalMux
    port map (
            O => \N__71445\,
            I => \N__71402\
        );

    \I__17475\ : Span4Mux_v
    port map (
            O => \N__71442\,
            I => \N__71402\
        );

    \I__17474\ : InMux
    port map (
            O => \N__71441\,
            I => \N__71396\
        );

    \I__17473\ : InMux
    port map (
            O => \N__71440\,
            I => \N__71391\
        );

    \I__17472\ : LocalMux
    port map (
            O => \N__71437\,
            I => \N__71388\
        );

    \I__17471\ : InMux
    port map (
            O => \N__71436\,
            I => \N__71385\
        );

    \I__17470\ : CascadeMux
    port map (
            O => \N__71435\,
            I => \N__71381\
        );

    \I__17469\ : Span4Mux_v
    port map (
            O => \N__71432\,
            I => \N__71377\
        );

    \I__17468\ : Span4Mux_h
    port map (
            O => \N__71429\,
            I => \N__71372\
        );

    \I__17467\ : LocalMux
    port map (
            O => \N__71426\,
            I => \N__71372\
        );

    \I__17466\ : InMux
    port map (
            O => \N__71425\,
            I => \N__71367\
        );

    \I__17465\ : InMux
    port map (
            O => \N__71424\,
            I => \N__71367\
        );

    \I__17464\ : InMux
    port map (
            O => \N__71423\,
            I => \N__71364\
        );

    \I__17463\ : LocalMux
    port map (
            O => \N__71418\,
            I => \N__71361\
        );

    \I__17462\ : LocalMux
    port map (
            O => \N__71411\,
            I => \N__71358\
        );

    \I__17461\ : InMux
    port map (
            O => \N__71410\,
            I => \N__71353\
        );

    \I__17460\ : InMux
    port map (
            O => \N__71407\,
            I => \N__71353\
        );

    \I__17459\ : Span4Mux_v
    port map (
            O => \N__71402\,
            I => \N__71350\
        );

    \I__17458\ : InMux
    port map (
            O => \N__71401\,
            I => \N__71347\
        );

    \I__17457\ : InMux
    port map (
            O => \N__71400\,
            I => \N__71344\
        );

    \I__17456\ : InMux
    port map (
            O => \N__71399\,
            I => \N__71341\
        );

    \I__17455\ : LocalMux
    port map (
            O => \N__71396\,
            I => \N__71338\
        );

    \I__17454\ : InMux
    port map (
            O => \N__71395\,
            I => \N__71333\
        );

    \I__17453\ : InMux
    port map (
            O => \N__71394\,
            I => \N__71333\
        );

    \I__17452\ : LocalMux
    port map (
            O => \N__71391\,
            I => \N__71330\
        );

    \I__17451\ : Span4Mux_v
    port map (
            O => \N__71388\,
            I => \N__71327\
        );

    \I__17450\ : LocalMux
    port map (
            O => \N__71385\,
            I => \N__71324\
        );

    \I__17449\ : CascadeMux
    port map (
            O => \N__71384\,
            I => \N__71321\
        );

    \I__17448\ : InMux
    port map (
            O => \N__71381\,
            I => \N__71315\
        );

    \I__17447\ : InMux
    port map (
            O => \N__71380\,
            I => \N__71315\
        );

    \I__17446\ : Span4Mux_h
    port map (
            O => \N__71377\,
            I => \N__71309\
        );

    \I__17445\ : Span4Mux_v
    port map (
            O => \N__71372\,
            I => \N__71309\
        );

    \I__17444\ : LocalMux
    port map (
            O => \N__71367\,
            I => \N__71304\
        );

    \I__17443\ : LocalMux
    port map (
            O => \N__71364\,
            I => \N__71304\
        );

    \I__17442\ : Span4Mux_v
    port map (
            O => \N__71361\,
            I => \N__71297\
        );

    \I__17441\ : Span4Mux_h
    port map (
            O => \N__71358\,
            I => \N__71297\
        );

    \I__17440\ : LocalMux
    port map (
            O => \N__71353\,
            I => \N__71297\
        );

    \I__17439\ : Span4Mux_v
    port map (
            O => \N__71350\,
            I => \N__71292\
        );

    \I__17438\ : LocalMux
    port map (
            O => \N__71347\,
            I => \N__71292\
        );

    \I__17437\ : LocalMux
    port map (
            O => \N__71344\,
            I => \N__71289\
        );

    \I__17436\ : LocalMux
    port map (
            O => \N__71341\,
            I => \N__71282\
        );

    \I__17435\ : Span4Mux_h
    port map (
            O => \N__71338\,
            I => \N__71282\
        );

    \I__17434\ : LocalMux
    port map (
            O => \N__71333\,
            I => \N__71282\
        );

    \I__17433\ : Span4Mux_v
    port map (
            O => \N__71330\,
            I => \N__71279\
        );

    \I__17432\ : Span4Mux_h
    port map (
            O => \N__71327\,
            I => \N__71274\
        );

    \I__17431\ : Span4Mux_v
    port map (
            O => \N__71324\,
            I => \N__71274\
        );

    \I__17430\ : InMux
    port map (
            O => \N__71321\,
            I => \N__71269\
        );

    \I__17429\ : InMux
    port map (
            O => \N__71320\,
            I => \N__71269\
        );

    \I__17428\ : LocalMux
    port map (
            O => \N__71315\,
            I => \N__71266\
        );

    \I__17427\ : InMux
    port map (
            O => \N__71314\,
            I => \N__71263\
        );

    \I__17426\ : Span4Mux_h
    port map (
            O => \N__71309\,
            I => \N__71260\
        );

    \I__17425\ : Span4Mux_v
    port map (
            O => \N__71304\,
            I => \N__71257\
        );

    \I__17424\ : Span4Mux_h
    port map (
            O => \N__71297\,
            I => \N__71254\
        );

    \I__17423\ : Span4Mux_h
    port map (
            O => \N__71292\,
            I => \N__71251\
        );

    \I__17422\ : Span4Mux_h
    port map (
            O => \N__71289\,
            I => \N__71248\
        );

    \I__17421\ : Span4Mux_v
    port map (
            O => \N__71282\,
            I => \N__71245\
        );

    \I__17420\ : Span4Mux_v
    port map (
            O => \N__71279\,
            I => \N__71236\
        );

    \I__17419\ : Span4Mux_h
    port map (
            O => \N__71274\,
            I => \N__71236\
        );

    \I__17418\ : LocalMux
    port map (
            O => \N__71269\,
            I => \N__71236\
        );

    \I__17417\ : Span4Mux_v
    port map (
            O => \N__71266\,
            I => \N__71236\
        );

    \I__17416\ : LocalMux
    port map (
            O => \N__71263\,
            I => \aluReadBus\
        );

    \I__17415\ : Odrv4
    port map (
            O => \N__71260\,
            I => \aluReadBus\
        );

    \I__17414\ : Odrv4
    port map (
            O => \N__71257\,
            I => \aluReadBus\
        );

    \I__17413\ : Odrv4
    port map (
            O => \N__71254\,
            I => \aluReadBus\
        );

    \I__17412\ : Odrv4
    port map (
            O => \N__71251\,
            I => \aluReadBus\
        );

    \I__17411\ : Odrv4
    port map (
            O => \N__71248\,
            I => \aluReadBus\
        );

    \I__17410\ : Odrv4
    port map (
            O => \N__71245\,
            I => \aluReadBus\
        );

    \I__17409\ : Odrv4
    port map (
            O => \N__71236\,
            I => \aluReadBus\
        );

    \I__17408\ : CascadeMux
    port map (
            O => \N__71219\,
            I => \ALU.un1_operation_13_0_cascade_\
        );

    \I__17407\ : CEMux
    port map (
            O => \N__71216\,
            I => \N__71208\
        );

    \I__17406\ : CEMux
    port map (
            O => \N__71215\,
            I => \N__71204\
        );

    \I__17405\ : CEMux
    port map (
            O => \N__71214\,
            I => \N__71201\
        );

    \I__17404\ : CEMux
    port map (
            O => \N__71213\,
            I => \N__71194\
        );

    \I__17403\ : CEMux
    port map (
            O => \N__71212\,
            I => \N__71190\
        );

    \I__17402\ : CEMux
    port map (
            O => \N__71211\,
            I => \N__71186\
        );

    \I__17401\ : LocalMux
    port map (
            O => \N__71208\,
            I => \N__71183\
        );

    \I__17400\ : CEMux
    port map (
            O => \N__71207\,
            I => \N__71180\
        );

    \I__17399\ : LocalMux
    port map (
            O => \N__71204\,
            I => \N__71177\
        );

    \I__17398\ : LocalMux
    port map (
            O => \N__71201\,
            I => \N__71173\
        );

    \I__17397\ : CEMux
    port map (
            O => \N__71200\,
            I => \N__71170\
        );

    \I__17396\ : CEMux
    port map (
            O => \N__71199\,
            I => \N__71167\
        );

    \I__17395\ : CEMux
    port map (
            O => \N__71198\,
            I => \N__71164\
        );

    \I__17394\ : CEMux
    port map (
            O => \N__71197\,
            I => \N__71160\
        );

    \I__17393\ : LocalMux
    port map (
            O => \N__71194\,
            I => \N__71157\
        );

    \I__17392\ : CEMux
    port map (
            O => \N__71193\,
            I => \N__71154\
        );

    \I__17391\ : LocalMux
    port map (
            O => \N__71190\,
            I => \N__71151\
        );

    \I__17390\ : CEMux
    port map (
            O => \N__71189\,
            I => \N__71148\
        );

    \I__17389\ : LocalMux
    port map (
            O => \N__71186\,
            I => \N__71145\
        );

    \I__17388\ : Span4Mux_h
    port map (
            O => \N__71183\,
            I => \N__71140\
        );

    \I__17387\ : LocalMux
    port map (
            O => \N__71180\,
            I => \N__71140\
        );

    \I__17386\ : Span4Mux_v
    port map (
            O => \N__71177\,
            I => \N__71137\
        );

    \I__17385\ : CEMux
    port map (
            O => \N__71176\,
            I => \N__71134\
        );

    \I__17384\ : Span4Mux_v
    port map (
            O => \N__71173\,
            I => \N__71131\
        );

    \I__17383\ : LocalMux
    port map (
            O => \N__71170\,
            I => \N__71128\
        );

    \I__17382\ : LocalMux
    port map (
            O => \N__71167\,
            I => \N__71125\
        );

    \I__17381\ : LocalMux
    port map (
            O => \N__71164\,
            I => \N__71122\
        );

    \I__17380\ : CEMux
    port map (
            O => \N__71163\,
            I => \N__71119\
        );

    \I__17379\ : LocalMux
    port map (
            O => \N__71160\,
            I => \N__71116\
        );

    \I__17378\ : Span4Mux_h
    port map (
            O => \N__71157\,
            I => \N__71113\
        );

    \I__17377\ : LocalMux
    port map (
            O => \N__71154\,
            I => \N__71110\
        );

    \I__17376\ : Span4Mux_h
    port map (
            O => \N__71151\,
            I => \N__71105\
        );

    \I__17375\ : LocalMux
    port map (
            O => \N__71148\,
            I => \N__71105\
        );

    \I__17374\ : Span4Mux_v
    port map (
            O => \N__71145\,
            I => \N__71102\
        );

    \I__17373\ : Span4Mux_v
    port map (
            O => \N__71140\,
            I => \N__71097\
        );

    \I__17372\ : Span4Mux_h
    port map (
            O => \N__71137\,
            I => \N__71097\
        );

    \I__17371\ : LocalMux
    port map (
            O => \N__71134\,
            I => \N__71094\
        );

    \I__17370\ : Span4Mux_h
    port map (
            O => \N__71131\,
            I => \N__71089\
        );

    \I__17369\ : Span4Mux_h
    port map (
            O => \N__71128\,
            I => \N__71089\
        );

    \I__17368\ : Span4Mux_v
    port map (
            O => \N__71125\,
            I => \N__71084\
        );

    \I__17367\ : Span4Mux_v
    port map (
            O => \N__71122\,
            I => \N__71084\
        );

    \I__17366\ : LocalMux
    port map (
            O => \N__71119\,
            I => \N__71081\
        );

    \I__17365\ : Span4Mux_v
    port map (
            O => \N__71116\,
            I => \N__71076\
        );

    \I__17364\ : Span4Mux_h
    port map (
            O => \N__71113\,
            I => \N__71076\
        );

    \I__17363\ : Span4Mux_v
    port map (
            O => \N__71110\,
            I => \N__71071\
        );

    \I__17362\ : Span4Mux_h
    port map (
            O => \N__71105\,
            I => \N__71071\
        );

    \I__17361\ : Span4Mux_h
    port map (
            O => \N__71102\,
            I => \N__71066\
        );

    \I__17360\ : Span4Mux_h
    port map (
            O => \N__71097\,
            I => \N__71066\
        );

    \I__17359\ : Span4Mux_h
    port map (
            O => \N__71094\,
            I => \N__71063\
        );

    \I__17358\ : Span4Mux_v
    port map (
            O => \N__71089\,
            I => \N__71060\
        );

    \I__17357\ : Span4Mux_v
    port map (
            O => \N__71084\,
            I => \N__71057\
        );

    \I__17356\ : Span4Mux_h
    port map (
            O => \N__71081\,
            I => \N__71052\
        );

    \I__17355\ : Span4Mux_h
    port map (
            O => \N__71076\,
            I => \N__71052\
        );

    \I__17354\ : Span4Mux_h
    port map (
            O => \N__71071\,
            I => \N__71049\
        );

    \I__17353\ : Span4Mux_h
    port map (
            O => \N__71066\,
            I => \N__71046\
        );

    \I__17352\ : Span4Mux_h
    port map (
            O => \N__71063\,
            I => \N__71043\
        );

    \I__17351\ : Span4Mux_h
    port map (
            O => \N__71060\,
            I => \N__71038\
        );

    \I__17350\ : Span4Mux_h
    port map (
            O => \N__71057\,
            I => \N__71038\
        );

    \I__17349\ : Span4Mux_h
    port map (
            O => \N__71052\,
            I => \N__71035\
        );

    \I__17348\ : Span4Mux_h
    port map (
            O => \N__71049\,
            I => \N__71030\
        );

    \I__17347\ : Span4Mux_v
    port map (
            O => \N__71046\,
            I => \N__71030\
        );

    \I__17346\ : Odrv4
    port map (
            O => \N__71043\,
            I => \ALU.un1_a41_9_0\
        );

    \I__17345\ : Odrv4
    port map (
            O => \N__71038\,
            I => \ALU.un1_a41_9_0\
        );

    \I__17344\ : Odrv4
    port map (
            O => \N__71035\,
            I => \ALU.un1_a41_9_0\
        );

    \I__17343\ : Odrv4
    port map (
            O => \N__71030\,
            I => \ALU.un1_a41_9_0\
        );

    \I__17342\ : InMux
    port map (
            O => \N__71021\,
            I => \N__71012\
        );

    \I__17341\ : InMux
    port map (
            O => \N__71020\,
            I => \N__71012\
        );

    \I__17340\ : InMux
    port map (
            O => \N__71019\,
            I => \N__71012\
        );

    \I__17339\ : LocalMux
    port map (
            O => \N__71012\,
            I => \ALU.un1_a41_3_0_1\
        );

    \I__17338\ : InMux
    port map (
            O => \N__71009\,
            I => \N__70997\
        );

    \I__17337\ : InMux
    port map (
            O => \N__71008\,
            I => \N__70997\
        );

    \I__17336\ : InMux
    port map (
            O => \N__71007\,
            I => \N__70997\
        );

    \I__17335\ : InMux
    port map (
            O => \N__71006\,
            I => \N__70997\
        );

    \I__17334\ : LocalMux
    port map (
            O => \N__70997\,
            I => \ALU.un1_operation_13_0\
        );

    \I__17333\ : CEMux
    port map (
            O => \N__70994\,
            I => \N__70990\
        );

    \I__17332\ : CEMux
    port map (
            O => \N__70993\,
            I => \N__70987\
        );

    \I__17331\ : LocalMux
    port map (
            O => \N__70990\,
            I => \N__70983\
        );

    \I__17330\ : LocalMux
    port map (
            O => \N__70987\,
            I => \N__70980\
        );

    \I__17329\ : CEMux
    port map (
            O => \N__70986\,
            I => \N__70977\
        );

    \I__17328\ : Span4Mux_h
    port map (
            O => \N__70983\,
            I => \N__70974\
        );

    \I__17327\ : Span4Mux_v
    port map (
            O => \N__70980\,
            I => \N__70971\
        );

    \I__17326\ : LocalMux
    port map (
            O => \N__70977\,
            I => \N__70968\
        );

    \I__17325\ : Span4Mux_h
    port map (
            O => \N__70974\,
            I => \N__70965\
        );

    \I__17324\ : Span4Mux_v
    port map (
            O => \N__70971\,
            I => \N__70962\
        );

    \I__17323\ : Span4Mux_h
    port map (
            O => \N__70968\,
            I => \N__70959\
        );

    \I__17322\ : Span4Mux_h
    port map (
            O => \N__70965\,
            I => \N__70956\
        );

    \I__17321\ : Sp12to4
    port map (
            O => \N__70962\,
            I => \N__70953\
        );

    \I__17320\ : Span4Mux_h
    port map (
            O => \N__70959\,
            I => \N__70948\
        );

    \I__17319\ : Span4Mux_v
    port map (
            O => \N__70956\,
            I => \N__70948\
        );

    \I__17318\ : Odrv12
    port map (
            O => \N__70953\,
            I => \ALU.un1_a41_3_0\
        );

    \I__17317\ : Odrv4
    port map (
            O => \N__70948\,
            I => \ALU.un1_a41_3_0\
        );

    \I__17316\ : CascadeMux
    port map (
            O => \N__70943\,
            I => \N__70937\
        );

    \I__17315\ : CascadeMux
    port map (
            O => \N__70942\,
            I => \N__70932\
        );

    \I__17314\ : InMux
    port map (
            O => \N__70941\,
            I => \N__70922\
        );

    \I__17313\ : InMux
    port map (
            O => \N__70940\,
            I => \N__70922\
        );

    \I__17312\ : InMux
    port map (
            O => \N__70937\,
            I => \N__70922\
        );

    \I__17311\ : InMux
    port map (
            O => \N__70936\,
            I => \N__70922\
        );

    \I__17310\ : InMux
    port map (
            O => \N__70935\,
            I => \N__70915\
        );

    \I__17309\ : InMux
    port map (
            O => \N__70932\,
            I => \N__70915\
        );

    \I__17308\ : InMux
    port map (
            O => \N__70931\,
            I => \N__70915\
        );

    \I__17307\ : LocalMux
    port map (
            O => \N__70922\,
            I => \N__70908\
        );

    \I__17306\ : LocalMux
    port map (
            O => \N__70915\,
            I => \N__70908\
        );

    \I__17305\ : InMux
    port map (
            O => \N__70914\,
            I => \N__70905\
        );

    \I__17304\ : InMux
    port map (
            O => \N__70913\,
            I => \N__70902\
        );

    \I__17303\ : Span4Mux_v
    port map (
            O => \N__70908\,
            I => \N__70897\
        );

    \I__17302\ : LocalMux
    port map (
            O => \N__70905\,
            I => \N__70897\
        );

    \I__17301\ : LocalMux
    port map (
            O => \N__70902\,
            I => \aluResults_2\
        );

    \I__17300\ : Odrv4
    port map (
            O => \N__70897\,
            I => \aluResults_2\
        );

    \I__17299\ : CascadeMux
    port map (
            O => \N__70892\,
            I => \N__70884\
        );

    \I__17298\ : InMux
    port map (
            O => \N__70891\,
            I => \N__70875\
        );

    \I__17297\ : InMux
    port map (
            O => \N__70890\,
            I => \N__70875\
        );

    \I__17296\ : InMux
    port map (
            O => \N__70889\,
            I => \N__70875\
        );

    \I__17295\ : InMux
    port map (
            O => \N__70888\,
            I => \N__70866\
        );

    \I__17294\ : InMux
    port map (
            O => \N__70887\,
            I => \N__70866\
        );

    \I__17293\ : InMux
    port map (
            O => \N__70884\,
            I => \N__70866\
        );

    \I__17292\ : InMux
    port map (
            O => \N__70883\,
            I => \N__70866\
        );

    \I__17291\ : InMux
    port map (
            O => \N__70882\,
            I => \N__70862\
        );

    \I__17290\ : LocalMux
    port map (
            O => \N__70875\,
            I => \N__70859\
        );

    \I__17289\ : LocalMux
    port map (
            O => \N__70866\,
            I => \N__70856\
        );

    \I__17288\ : InMux
    port map (
            O => \N__70865\,
            I => \N__70853\
        );

    \I__17287\ : LocalMux
    port map (
            O => \N__70862\,
            I => \aluResults_1\
        );

    \I__17286\ : Odrv4
    port map (
            O => \N__70859\,
            I => \aluResults_1\
        );

    \I__17285\ : Odrv4
    port map (
            O => \N__70856\,
            I => \aluResults_1\
        );

    \I__17284\ : LocalMux
    port map (
            O => \N__70853\,
            I => \aluResults_1\
        );

    \I__17283\ : CascadeMux
    port map (
            O => \N__70844\,
            I => \N__70841\
        );

    \I__17282\ : InMux
    port map (
            O => \N__70841\,
            I => \N__70838\
        );

    \I__17281\ : LocalMux
    port map (
            O => \N__70838\,
            I => \ALU.un1_a41_2Z0Z_1\
        );

    \I__17280\ : InMux
    port map (
            O => \N__70835\,
            I => \N__70832\
        );

    \I__17279\ : LocalMux
    port map (
            O => \N__70832\,
            I => \N__70829\
        );

    \I__17278\ : Span4Mux_v
    port map (
            O => \N__70829\,
            I => \N__70825\
        );

    \I__17277\ : InMux
    port map (
            O => \N__70828\,
            I => \N__70822\
        );

    \I__17276\ : Sp12to4
    port map (
            O => \N__70825\,
            I => \N__70819\
        );

    \I__17275\ : LocalMux
    port map (
            O => \N__70822\,
            I => \N__70816\
        );

    \I__17274\ : Span12Mux_h
    port map (
            O => \N__70819\,
            I => \N__70812\
        );

    \I__17273\ : Span4Mux_h
    port map (
            O => \N__70816\,
            I => \N__70809\
        );

    \I__17272\ : InMux
    port map (
            O => \N__70815\,
            I => \N__70806\
        );

    \I__17271\ : Odrv12
    port map (
            O => \N__70812\,
            I => \controlWord_22\
        );

    \I__17270\ : Odrv4
    port map (
            O => \N__70809\,
            I => \controlWord_22\
        );

    \I__17269\ : LocalMux
    port map (
            O => \N__70806\,
            I => \controlWord_22\
        );

    \I__17268\ : InMux
    port map (
            O => \N__70799\,
            I => \N__70791\
        );

    \I__17267\ : CascadeMux
    port map (
            O => \N__70798\,
            I => \N__70782\
        );

    \I__17266\ : CascadeMux
    port map (
            O => \N__70797\,
            I => \N__70779\
        );

    \I__17265\ : CascadeMux
    port map (
            O => \N__70796\,
            I => \N__70776\
        );

    \I__17264\ : InMux
    port map (
            O => \N__70795\,
            I => \N__70773\
        );

    \I__17263\ : InMux
    port map (
            O => \N__70794\,
            I => \N__70770\
        );

    \I__17262\ : LocalMux
    port map (
            O => \N__70791\,
            I => \N__70767\
        );

    \I__17261\ : InMux
    port map (
            O => \N__70790\,
            I => \N__70751\
        );

    \I__17260\ : InMux
    port map (
            O => \N__70789\,
            I => \N__70746\
        );

    \I__17259\ : InMux
    port map (
            O => \N__70788\,
            I => \N__70746\
        );

    \I__17258\ : InMux
    port map (
            O => \N__70787\,
            I => \N__70733\
        );

    \I__17257\ : InMux
    port map (
            O => \N__70786\,
            I => \N__70733\
        );

    \I__17256\ : InMux
    port map (
            O => \N__70785\,
            I => \N__70733\
        );

    \I__17255\ : InMux
    port map (
            O => \N__70782\,
            I => \N__70733\
        );

    \I__17254\ : InMux
    port map (
            O => \N__70779\,
            I => \N__70733\
        );

    \I__17253\ : InMux
    port map (
            O => \N__70776\,
            I => \N__70733\
        );

    \I__17252\ : LocalMux
    port map (
            O => \N__70773\,
            I => \N__70730\
        );

    \I__17251\ : LocalMux
    port map (
            O => \N__70770\,
            I => \N__70727\
        );

    \I__17250\ : Span4Mux_v
    port map (
            O => \N__70767\,
            I => \N__70724\
        );

    \I__17249\ : CascadeMux
    port map (
            O => \N__70766\,
            I => \N__70718\
        );

    \I__17248\ : CascadeMux
    port map (
            O => \N__70765\,
            I => \N__70715\
        );

    \I__17247\ : CascadeMux
    port map (
            O => \N__70764\,
            I => \N__70712\
        );

    \I__17246\ : InMux
    port map (
            O => \N__70763\,
            I => \N__70703\
        );

    \I__17245\ : InMux
    port map (
            O => \N__70762\,
            I => \N__70703\
        );

    \I__17244\ : InMux
    port map (
            O => \N__70761\,
            I => \N__70700\
        );

    \I__17243\ : InMux
    port map (
            O => \N__70760\,
            I => \N__70693\
        );

    \I__17242\ : InMux
    port map (
            O => \N__70759\,
            I => \N__70693\
        );

    \I__17241\ : InMux
    port map (
            O => \N__70758\,
            I => \N__70693\
        );

    \I__17240\ : InMux
    port map (
            O => \N__70757\,
            I => \N__70690\
        );

    \I__17239\ : InMux
    port map (
            O => \N__70756\,
            I => \N__70683\
        );

    \I__17238\ : InMux
    port map (
            O => \N__70755\,
            I => \N__70683\
        );

    \I__17237\ : InMux
    port map (
            O => \N__70754\,
            I => \N__70683\
        );

    \I__17236\ : LocalMux
    port map (
            O => \N__70751\,
            I => \N__70678\
        );

    \I__17235\ : LocalMux
    port map (
            O => \N__70746\,
            I => \N__70678\
        );

    \I__17234\ : LocalMux
    port map (
            O => \N__70733\,
            I => \N__70671\
        );

    \I__17233\ : Span4Mux_h
    port map (
            O => \N__70730\,
            I => \N__70671\
        );

    \I__17232\ : Span4Mux_v
    port map (
            O => \N__70727\,
            I => \N__70671\
        );

    \I__17231\ : Span4Mux_h
    port map (
            O => \N__70724\,
            I => \N__70668\
        );

    \I__17230\ : InMux
    port map (
            O => \N__70723\,
            I => \N__70661\
        );

    \I__17229\ : InMux
    port map (
            O => \N__70722\,
            I => \N__70661\
        );

    \I__17228\ : InMux
    port map (
            O => \N__70721\,
            I => \N__70661\
        );

    \I__17227\ : InMux
    port map (
            O => \N__70718\,
            I => \N__70646\
        );

    \I__17226\ : InMux
    port map (
            O => \N__70715\,
            I => \N__70646\
        );

    \I__17225\ : InMux
    port map (
            O => \N__70712\,
            I => \N__70646\
        );

    \I__17224\ : InMux
    port map (
            O => \N__70711\,
            I => \N__70646\
        );

    \I__17223\ : InMux
    port map (
            O => \N__70710\,
            I => \N__70646\
        );

    \I__17222\ : InMux
    port map (
            O => \N__70709\,
            I => \N__70646\
        );

    \I__17221\ : InMux
    port map (
            O => \N__70708\,
            I => \N__70646\
        );

    \I__17220\ : LocalMux
    port map (
            O => \N__70703\,
            I => \N__70643\
        );

    \I__17219\ : LocalMux
    port map (
            O => \N__70700\,
            I => \N__70640\
        );

    \I__17218\ : LocalMux
    port map (
            O => \N__70693\,
            I => \N__70631\
        );

    \I__17217\ : LocalMux
    port map (
            O => \N__70690\,
            I => \N__70631\
        );

    \I__17216\ : LocalMux
    port map (
            O => \N__70683\,
            I => \N__70631\
        );

    \I__17215\ : Span12Mux_h
    port map (
            O => \N__70678\,
            I => \N__70631\
        );

    \I__17214\ : Span4Mux_h
    port map (
            O => \N__70671\,
            I => \N__70626\
        );

    \I__17213\ : Span4Mux_h
    port map (
            O => \N__70668\,
            I => \N__70626\
        );

    \I__17212\ : LocalMux
    port map (
            O => \N__70661\,
            I => \CONTROL.un1_busState101_3_0_0_0\
        );

    \I__17211\ : LocalMux
    port map (
            O => \N__70646\,
            I => \CONTROL.un1_busState101_3_0_0_0\
        );

    \I__17210\ : Odrv4
    port map (
            O => \N__70643\,
            I => \CONTROL.un1_busState101_3_0_0_0\
        );

    \I__17209\ : Odrv12
    port map (
            O => \N__70640\,
            I => \CONTROL.un1_busState101_3_0_0_0\
        );

    \I__17208\ : Odrv12
    port map (
            O => \N__70631\,
            I => \CONTROL.un1_busState101_3_0_0_0\
        );

    \I__17207\ : Odrv4
    port map (
            O => \N__70626\,
            I => \CONTROL.un1_busState101_3_0_0_0\
        );

    \I__17206\ : CascadeMux
    port map (
            O => \N__70613\,
            I => \N__70610\
        );

    \I__17205\ : InMux
    port map (
            O => \N__70610\,
            I => \N__70607\
        );

    \I__17204\ : LocalMux
    port map (
            O => \N__70607\,
            I => \N__70604\
        );

    \I__17203\ : Span4Mux_v
    port map (
            O => \N__70604\,
            I => \N__70600\
        );

    \I__17202\ : InMux
    port map (
            O => \N__70603\,
            I => \N__70597\
        );

    \I__17201\ : Span4Mux_h
    port map (
            O => \N__70600\,
            I => \N__70594\
        );

    \I__17200\ : LocalMux
    port map (
            O => \N__70597\,
            I => \N__70591\
        );

    \I__17199\ : Span4Mux_h
    port map (
            O => \N__70594\,
            I => \N__70586\
        );

    \I__17198\ : Span4Mux_h
    port map (
            O => \N__70591\,
            I => \N__70586\
        );

    \I__17197\ : Span4Mux_v
    port map (
            O => \N__70586\,
            I => \N__70582\
        );

    \I__17196\ : InMux
    port map (
            O => \N__70585\,
            I => \N__70579\
        );

    \I__17195\ : Span4Mux_v
    port map (
            O => \N__70582\,
            I => \N__70576\
        );

    \I__17194\ : LocalMux
    port map (
            O => \N__70579\,
            I => \N__70573\
        );

    \I__17193\ : Sp12to4
    port map (
            O => \N__70576\,
            I => \N__70570\
        );

    \I__17192\ : Span4Mux_h
    port map (
            O => \N__70573\,
            I => \N__70567\
        );

    \I__17191\ : Span12Mux_s8_v
    port map (
            O => \N__70570\,
            I => \N__70564\
        );

    \I__17190\ : Span4Mux_h
    port map (
            O => \N__70567\,
            I => \N__70561\
        );

    \I__17189\ : Odrv12
    port map (
            O => \N__70564\,
            I => f_6
        );

    \I__17188\ : Odrv4
    port map (
            O => \N__70561\,
            I => f_6
        );

    \I__17187\ : InMux
    port map (
            O => \N__70556\,
            I => \N__70553\
        );

    \I__17186\ : LocalMux
    port map (
            O => \N__70553\,
            I => \N__70545\
        );

    \I__17185\ : InMux
    port map (
            O => \N__70552\,
            I => \N__70536\
        );

    \I__17184\ : InMux
    port map (
            O => \N__70551\,
            I => \N__70528\
        );

    \I__17183\ : InMux
    port map (
            O => \N__70550\,
            I => \N__70528\
        );

    \I__17182\ : InMux
    port map (
            O => \N__70549\,
            I => \N__70528\
        );

    \I__17181\ : InMux
    port map (
            O => \N__70548\,
            I => \N__70518\
        );

    \I__17180\ : Span4Mux_h
    port map (
            O => \N__70545\,
            I => \N__70515\
        );

    \I__17179\ : CascadeMux
    port map (
            O => \N__70544\,
            I => \N__70511\
        );

    \I__17178\ : InMux
    port map (
            O => \N__70543\,
            I => \N__70500\
        );

    \I__17177\ : InMux
    port map (
            O => \N__70542\,
            I => \N__70500\
        );

    \I__17176\ : InMux
    port map (
            O => \N__70541\,
            I => \N__70500\
        );

    \I__17175\ : InMux
    port map (
            O => \N__70540\,
            I => \N__70500\
        );

    \I__17174\ : InMux
    port map (
            O => \N__70539\,
            I => \N__70500\
        );

    \I__17173\ : LocalMux
    port map (
            O => \N__70536\,
            I => \N__70497\
        );

    \I__17172\ : InMux
    port map (
            O => \N__70535\,
            I => \N__70494\
        );

    \I__17171\ : LocalMux
    port map (
            O => \N__70528\,
            I => \N__70491\
        );

    \I__17170\ : InMux
    port map (
            O => \N__70527\,
            I => \N__70478\
        );

    \I__17169\ : InMux
    port map (
            O => \N__70526\,
            I => \N__70478\
        );

    \I__17168\ : InMux
    port map (
            O => \N__70525\,
            I => \N__70478\
        );

    \I__17167\ : InMux
    port map (
            O => \N__70524\,
            I => \N__70478\
        );

    \I__17166\ : InMux
    port map (
            O => \N__70523\,
            I => \N__70478\
        );

    \I__17165\ : InMux
    port map (
            O => \N__70522\,
            I => \N__70478\
        );

    \I__17164\ : InMux
    port map (
            O => \N__70521\,
            I => \N__70475\
        );

    \I__17163\ : LocalMux
    port map (
            O => \N__70518\,
            I => \N__70472\
        );

    \I__17162\ : Span4Mux_h
    port map (
            O => \N__70515\,
            I => \N__70469\
        );

    \I__17161\ : InMux
    port map (
            O => \N__70514\,
            I => \N__70463\
        );

    \I__17160\ : InMux
    port map (
            O => \N__70511\,
            I => \N__70452\
        );

    \I__17159\ : LocalMux
    port map (
            O => \N__70500\,
            I => \N__70445\
        );

    \I__17158\ : Span4Mux_h
    port map (
            O => \N__70497\,
            I => \N__70445\
        );

    \I__17157\ : LocalMux
    port map (
            O => \N__70494\,
            I => \N__70445\
        );

    \I__17156\ : Span4Mux_h
    port map (
            O => \N__70491\,
            I => \N__70442\
        );

    \I__17155\ : LocalMux
    port map (
            O => \N__70478\,
            I => \N__70437\
        );

    \I__17154\ : LocalMux
    port map (
            O => \N__70475\,
            I => \N__70437\
        );

    \I__17153\ : Span4Mux_h
    port map (
            O => \N__70472\,
            I => \N__70432\
        );

    \I__17152\ : Span4Mux_h
    port map (
            O => \N__70469\,
            I => \N__70432\
        );

    \I__17151\ : InMux
    port map (
            O => \N__70468\,
            I => \N__70425\
        );

    \I__17150\ : InMux
    port map (
            O => \N__70467\,
            I => \N__70425\
        );

    \I__17149\ : InMux
    port map (
            O => \N__70466\,
            I => \N__70425\
        );

    \I__17148\ : LocalMux
    port map (
            O => \N__70463\,
            I => \N__70422\
        );

    \I__17147\ : InMux
    port map (
            O => \N__70462\,
            I => \N__70417\
        );

    \I__17146\ : InMux
    port map (
            O => \N__70461\,
            I => \N__70417\
        );

    \I__17145\ : InMux
    port map (
            O => \N__70460\,
            I => \N__70404\
        );

    \I__17144\ : InMux
    port map (
            O => \N__70459\,
            I => \N__70404\
        );

    \I__17143\ : InMux
    port map (
            O => \N__70458\,
            I => \N__70404\
        );

    \I__17142\ : InMux
    port map (
            O => \N__70457\,
            I => \N__70404\
        );

    \I__17141\ : InMux
    port map (
            O => \N__70456\,
            I => \N__70404\
        );

    \I__17140\ : InMux
    port map (
            O => \N__70455\,
            I => \N__70404\
        );

    \I__17139\ : LocalMux
    port map (
            O => \N__70452\,
            I => \N__70401\
        );

    \I__17138\ : Span4Mux_h
    port map (
            O => \N__70445\,
            I => \N__70398\
        );

    \I__17137\ : Span4Mux_h
    port map (
            O => \N__70442\,
            I => \N__70395\
        );

    \I__17136\ : Span4Mux_v
    port map (
            O => \N__70437\,
            I => \N__70390\
        );

    \I__17135\ : Span4Mux_h
    port map (
            O => \N__70432\,
            I => \N__70390\
        );

    \I__17134\ : LocalMux
    port map (
            O => \N__70425\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17133\ : Odrv4
    port map (
            O => \N__70422\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17132\ : LocalMux
    port map (
            O => \N__70417\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17131\ : LocalMux
    port map (
            O => \N__70404\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17130\ : Odrv4
    port map (
            O => \N__70401\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17129\ : Odrv4
    port map (
            O => \N__70398\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17128\ : Odrv4
    port map (
            O => \N__70395\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17127\ : Odrv4
    port map (
            O => \N__70390\,
            I => \CONTROL.un1_busState101_3_0Z0Z_1\
        );

    \I__17126\ : IoInMux
    port map (
            O => \N__70373\,
            I => \N__70370\
        );

    \I__17125\ : LocalMux
    port map (
            O => \N__70370\,
            I => \N__70366\
        );

    \I__17124\ : InMux
    port map (
            O => \N__70369\,
            I => \N__70363\
        );

    \I__17123\ : Span4Mux_s3_h
    port map (
            O => \N__70366\,
            I => \N__70360\
        );

    \I__17122\ : LocalMux
    port map (
            O => \N__70363\,
            I => \N__70357\
        );

    \I__17121\ : Sp12to4
    port map (
            O => \N__70360\,
            I => \N__70354\
        );

    \I__17120\ : Span12Mux_v
    port map (
            O => \N__70357\,
            I => \N__70351\
        );

    \I__17119\ : Span12Mux_v
    port map (
            O => \N__70354\,
            I => \N__70348\
        );

    \I__17118\ : Span12Mux_h
    port map (
            O => \N__70351\,
            I => \N__70345\
        );

    \I__17117\ : Odrv12
    port map (
            O => \N__70348\,
            I => \A6_c\
        );

    \I__17116\ : Odrv12
    port map (
            O => \N__70345\,
            I => \A6_c\
        );

    \I__17115\ : CEMux
    port map (
            O => \N__70340\,
            I => \N__70337\
        );

    \I__17114\ : LocalMux
    port map (
            O => \N__70337\,
            I => \N__70334\
        );

    \I__17113\ : Span4Mux_v
    port map (
            O => \N__70334\,
            I => \N__70331\
        );

    \I__17112\ : Span4Mux_h
    port map (
            O => \N__70331\,
            I => \N__70325\
        );

    \I__17111\ : CEMux
    port map (
            O => \N__70330\,
            I => \N__70322\
        );

    \I__17110\ : CEMux
    port map (
            O => \N__70329\,
            I => \N__70319\
        );

    \I__17109\ : CEMux
    port map (
            O => \N__70328\,
            I => \N__70314\
        );

    \I__17108\ : Span4Mux_v
    port map (
            O => \N__70325\,
            I => \N__70309\
        );

    \I__17107\ : LocalMux
    port map (
            O => \N__70322\,
            I => \N__70309\
        );

    \I__17106\ : LocalMux
    port map (
            O => \N__70319\,
            I => \N__70306\
        );

    \I__17105\ : CEMux
    port map (
            O => \N__70318\,
            I => \N__70303\
        );

    \I__17104\ : CEMux
    port map (
            O => \N__70317\,
            I => \N__70300\
        );

    \I__17103\ : LocalMux
    port map (
            O => \N__70314\,
            I => \N__70297\
        );

    \I__17102\ : Span4Mux_h
    port map (
            O => \N__70309\,
            I => \N__70292\
        );

    \I__17101\ : Span4Mux_v
    port map (
            O => \N__70306\,
            I => \N__70292\
        );

    \I__17100\ : LocalMux
    port map (
            O => \N__70303\,
            I => \N__70285\
        );

    \I__17099\ : LocalMux
    port map (
            O => \N__70300\,
            I => \N__70285\
        );

    \I__17098\ : Span4Mux_v
    port map (
            O => \N__70297\,
            I => \N__70285\
        );

    \I__17097\ : Span4Mux_h
    port map (
            O => \N__70292\,
            I => \N__70282\
        );

    \I__17096\ : Span4Mux_v
    port map (
            O => \N__70285\,
            I => \N__70279\
        );

    \I__17095\ : Sp12to4
    port map (
            O => \N__70282\,
            I => \N__70276\
        );

    \I__17094\ : Odrv4
    port map (
            O => \N__70279\,
            I => \CONTROL.N_60\
        );

    \I__17093\ : Odrv12
    port map (
            O => \N__70276\,
            I => \CONTROL.N_60\
        );

    \I__17092\ : CascadeMux
    port map (
            O => \N__70271\,
            I => \PROM.ROMDATA.m281_cascade_\
        );

    \I__17091\ : InMux
    port map (
            O => \N__70268\,
            I => \N__70265\
        );

    \I__17090\ : LocalMux
    port map (
            O => \N__70265\,
            I => \ALU.un1_a41_7_0_2\
        );

    \I__17089\ : CascadeMux
    port map (
            O => \N__70262\,
            I => \ALU.un1_operation_13Z0Z_2_cascade_\
        );

    \I__17088\ : InMux
    port map (
            O => \N__70259\,
            I => \N__70256\
        );

    \I__17087\ : LocalMux
    port map (
            O => \N__70256\,
            I => \ALU.un1_a41_4_0_2\
        );

    \I__17086\ : CascadeMux
    port map (
            O => \N__70253\,
            I => \ALU.un1_a41_4_0_2_cascade_\
        );

    \I__17085\ : CEMux
    port map (
            O => \N__70250\,
            I => \N__70246\
        );

    \I__17084\ : CEMux
    port map (
            O => \N__70249\,
            I => \N__70243\
        );

    \I__17083\ : LocalMux
    port map (
            O => \N__70246\,
            I => \N__70240\
        );

    \I__17082\ : LocalMux
    port map (
            O => \N__70243\,
            I => \N__70236\
        );

    \I__17081\ : Span4Mux_h
    port map (
            O => \N__70240\,
            I => \N__70233\
        );

    \I__17080\ : CEMux
    port map (
            O => \N__70239\,
            I => \N__70230\
        );

    \I__17079\ : Span4Mux_h
    port map (
            O => \N__70236\,
            I => \N__70227\
        );

    \I__17078\ : Span4Mux_h
    port map (
            O => \N__70233\,
            I => \N__70224\
        );

    \I__17077\ : LocalMux
    port map (
            O => \N__70230\,
            I => \N__70221\
        );

    \I__17076\ : Span4Mux_h
    port map (
            O => \N__70227\,
            I => \N__70218\
        );

    \I__17075\ : Span4Mux_v
    port map (
            O => \N__70224\,
            I => \N__70215\
        );

    \I__17074\ : Span4Mux_v
    port map (
            O => \N__70221\,
            I => \N__70212\
        );

    \I__17073\ : Span4Mux_v
    port map (
            O => \N__70218\,
            I => \N__70209\
        );

    \I__17072\ : Sp12to4
    port map (
            O => \N__70215\,
            I => \N__70206\
        );

    \I__17071\ : Odrv4
    port map (
            O => \N__70212\,
            I => \ALU.un1_a41_6_0\
        );

    \I__17070\ : Odrv4
    port map (
            O => \N__70209\,
            I => \ALU.un1_a41_6_0\
        );

    \I__17069\ : Odrv12
    port map (
            O => \N__70206\,
            I => \ALU.un1_a41_6_0\
        );

    \I__17068\ : InMux
    port map (
            O => \N__70199\,
            I => \N__70192\
        );

    \I__17067\ : InMux
    port map (
            O => \N__70198\,
            I => \N__70192\
        );

    \I__17066\ : InMux
    port map (
            O => \N__70197\,
            I => \N__70188\
        );

    \I__17065\ : LocalMux
    port map (
            O => \N__70192\,
            I => \N__70181\
        );

    \I__17064\ : InMux
    port map (
            O => \N__70191\,
            I => \N__70178\
        );

    \I__17063\ : LocalMux
    port map (
            O => \N__70188\,
            I => \N__70175\
        );

    \I__17062\ : InMux
    port map (
            O => \N__70187\,
            I => \N__70172\
        );

    \I__17061\ : InMux
    port map (
            O => \N__70186\,
            I => \N__70160\
        );

    \I__17060\ : InMux
    port map (
            O => \N__70185\,
            I => \N__70160\
        );

    \I__17059\ : InMux
    port map (
            O => \N__70184\,
            I => \N__70160\
        );

    \I__17058\ : Span4Mux_v
    port map (
            O => \N__70181\,
            I => \N__70154\
        );

    \I__17057\ : LocalMux
    port map (
            O => \N__70178\,
            I => \N__70147\
        );

    \I__17056\ : Span4Mux_v
    port map (
            O => \N__70175\,
            I => \N__70147\
        );

    \I__17055\ : LocalMux
    port map (
            O => \N__70172\,
            I => \N__70147\
        );

    \I__17054\ : InMux
    port map (
            O => \N__70171\,
            I => \N__70140\
        );

    \I__17053\ : InMux
    port map (
            O => \N__70170\,
            I => \N__70140\
        );

    \I__17052\ : InMux
    port map (
            O => \N__70169\,
            I => \N__70140\
        );

    \I__17051\ : InMux
    port map (
            O => \N__70168\,
            I => \N__70134\
        );

    \I__17050\ : InMux
    port map (
            O => \N__70167\,
            I => \N__70134\
        );

    \I__17049\ : LocalMux
    port map (
            O => \N__70160\,
            I => \N__70131\
        );

    \I__17048\ : InMux
    port map (
            O => \N__70159\,
            I => \N__70128\
        );

    \I__17047\ : InMux
    port map (
            O => \N__70158\,
            I => \N__70123\
        );

    \I__17046\ : InMux
    port map (
            O => \N__70157\,
            I => \N__70123\
        );

    \I__17045\ : Span4Mux_h
    port map (
            O => \N__70154\,
            I => \N__70118\
        );

    \I__17044\ : Span4Mux_v
    port map (
            O => \N__70147\,
            I => \N__70118\
        );

    \I__17043\ : LocalMux
    port map (
            O => \N__70140\,
            I => \N__70114\
        );

    \I__17042\ : InMux
    port map (
            O => \N__70139\,
            I => \N__70111\
        );

    \I__17041\ : LocalMux
    port map (
            O => \N__70134\,
            I => \N__70106\
        );

    \I__17040\ : Span4Mux_h
    port map (
            O => \N__70131\,
            I => \N__70106\
        );

    \I__17039\ : LocalMux
    port map (
            O => \N__70128\,
            I => \N__70103\
        );

    \I__17038\ : LocalMux
    port map (
            O => \N__70123\,
            I => \N__70100\
        );

    \I__17037\ : Span4Mux_h
    port map (
            O => \N__70118\,
            I => \N__70097\
        );

    \I__17036\ : InMux
    port map (
            O => \N__70117\,
            I => \N__70091\
        );

    \I__17035\ : Span4Mux_v
    port map (
            O => \N__70114\,
            I => \N__70085\
        );

    \I__17034\ : LocalMux
    port map (
            O => \N__70111\,
            I => \N__70080\
        );

    \I__17033\ : Span4Mux_v
    port map (
            O => \N__70106\,
            I => \N__70080\
        );

    \I__17032\ : Span4Mux_v
    port map (
            O => \N__70103\,
            I => \N__70075\
        );

    \I__17031\ : Span4Mux_v
    port map (
            O => \N__70100\,
            I => \N__70075\
        );

    \I__17030\ : Sp12to4
    port map (
            O => \N__70097\,
            I => \N__70072\
        );

    \I__17029\ : InMux
    port map (
            O => \N__70096\,
            I => \N__70065\
        );

    \I__17028\ : InMux
    port map (
            O => \N__70095\,
            I => \N__70065\
        );

    \I__17027\ : InMux
    port map (
            O => \N__70094\,
            I => \N__70065\
        );

    \I__17026\ : LocalMux
    port map (
            O => \N__70091\,
            I => \N__70062\
        );

    \I__17025\ : InMux
    port map (
            O => \N__70090\,
            I => \N__70055\
        );

    \I__17024\ : InMux
    port map (
            O => \N__70089\,
            I => \N__70055\
        );

    \I__17023\ : InMux
    port map (
            O => \N__70088\,
            I => \N__70055\
        );

    \I__17022\ : Span4Mux_v
    port map (
            O => \N__70085\,
            I => \N__70047\
        );

    \I__17021\ : Span4Mux_v
    port map (
            O => \N__70080\,
            I => \N__70047\
        );

    \I__17020\ : Span4Mux_h
    port map (
            O => \N__70075\,
            I => \N__70047\
        );

    \I__17019\ : Span12Mux_h
    port map (
            O => \N__70072\,
            I => \N__70042\
        );

    \I__17018\ : LocalMux
    port map (
            O => \N__70065\,
            I => \N__70042\
        );

    \I__17017\ : Span4Mux_h
    port map (
            O => \N__70062\,
            I => \N__70037\
        );

    \I__17016\ : LocalMux
    port map (
            O => \N__70055\,
            I => \N__70037\
        );

    \I__17015\ : InMux
    port map (
            O => \N__70054\,
            I => \N__70034\
        );

    \I__17014\ : Span4Mux_h
    port map (
            O => \N__70047\,
            I => \N__70031\
        );

    \I__17013\ : Span12Mux_v
    port map (
            O => \N__70042\,
            I => \N__70028\
        );

    \I__17012\ : Sp12to4
    port map (
            O => \N__70037\,
            I => \N__70025\
        );

    \I__17011\ : LocalMux
    port map (
            O => \N__70034\,
            I => \aluOperation_2\
        );

    \I__17010\ : Odrv4
    port map (
            O => \N__70031\,
            I => \aluOperation_2\
        );

    \I__17009\ : Odrv12
    port map (
            O => \N__70028\,
            I => \aluOperation_2\
        );

    \I__17008\ : Odrv12
    port map (
            O => \N__70025\,
            I => \aluOperation_2\
        );

    \I__17007\ : CascadeMux
    port map (
            O => \N__70016\,
            I => \N__70013\
        );

    \I__17006\ : InMux
    port map (
            O => \N__70013\,
            I => \N__70008\
        );

    \I__17005\ : CascadeMux
    port map (
            O => \N__70012\,
            I => \N__70004\
        );

    \I__17004\ : CascadeMux
    port map (
            O => \N__70011\,
            I => \N__70001\
        );

    \I__17003\ : LocalMux
    port map (
            O => \N__70008\,
            I => \N__69995\
        );

    \I__17002\ : InMux
    port map (
            O => \N__70007\,
            I => \N__69992\
        );

    \I__17001\ : InMux
    port map (
            O => \N__70004\,
            I => \N__69989\
        );

    \I__17000\ : InMux
    port map (
            O => \N__70001\,
            I => \N__69983\
        );

    \I__16999\ : InMux
    port map (
            O => \N__70000\,
            I => \N__69983\
        );

    \I__16998\ : InMux
    port map (
            O => \N__69999\,
            I => \N__69978\
        );

    \I__16997\ : InMux
    port map (
            O => \N__69998\,
            I => \N__69978\
        );

    \I__16996\ : Span4Mux_v
    port map (
            O => \N__69995\,
            I => \N__69974\
        );

    \I__16995\ : LocalMux
    port map (
            O => \N__69992\,
            I => \N__69969\
        );

    \I__16994\ : LocalMux
    port map (
            O => \N__69989\,
            I => \N__69962\
        );

    \I__16993\ : InMux
    port map (
            O => \N__69988\,
            I => \N__69959\
        );

    \I__16992\ : LocalMux
    port map (
            O => \N__69983\,
            I => \N__69954\
        );

    \I__16991\ : LocalMux
    port map (
            O => \N__69978\,
            I => \N__69954\
        );

    \I__16990\ : InMux
    port map (
            O => \N__69977\,
            I => \N__69951\
        );

    \I__16989\ : Span4Mux_h
    port map (
            O => \N__69974\,
            I => \N__69948\
        );

    \I__16988\ : InMux
    port map (
            O => \N__69973\,
            I => \N__69945\
        );

    \I__16987\ : InMux
    port map (
            O => \N__69972\,
            I => \N__69940\
        );

    \I__16986\ : Span4Mux_v
    port map (
            O => \N__69969\,
            I => \N__69937\
        );

    \I__16985\ : InMux
    port map (
            O => \N__69968\,
            I => \N__69932\
        );

    \I__16984\ : InMux
    port map (
            O => \N__69967\,
            I => \N__69932\
        );

    \I__16983\ : InMux
    port map (
            O => \N__69966\,
            I => \N__69929\
        );

    \I__16982\ : CascadeMux
    port map (
            O => \N__69965\,
            I => \N__69925\
        );

    \I__16981\ : Span4Mux_v
    port map (
            O => \N__69962\,
            I => \N__69922\
        );

    \I__16980\ : LocalMux
    port map (
            O => \N__69959\,
            I => \N__69919\
        );

    \I__16979\ : Span4Mux_v
    port map (
            O => \N__69954\,
            I => \N__69914\
        );

    \I__16978\ : LocalMux
    port map (
            O => \N__69951\,
            I => \N__69914\
        );

    \I__16977\ : Span4Mux_h
    port map (
            O => \N__69948\,
            I => \N__69909\
        );

    \I__16976\ : LocalMux
    port map (
            O => \N__69945\,
            I => \N__69909\
        );

    \I__16975\ : InMux
    port map (
            O => \N__69944\,
            I => \N__69904\
        );

    \I__16974\ : InMux
    port map (
            O => \N__69943\,
            I => \N__69901\
        );

    \I__16973\ : LocalMux
    port map (
            O => \N__69940\,
            I => \N__69898\
        );

    \I__16972\ : Span4Mux_v
    port map (
            O => \N__69937\,
            I => \N__69891\
        );

    \I__16971\ : LocalMux
    port map (
            O => \N__69932\,
            I => \N__69891\
        );

    \I__16970\ : LocalMux
    port map (
            O => \N__69929\,
            I => \N__69891\
        );

    \I__16969\ : InMux
    port map (
            O => \N__69928\,
            I => \N__69886\
        );

    \I__16968\ : InMux
    port map (
            O => \N__69925\,
            I => \N__69886\
        );

    \I__16967\ : Span4Mux_v
    port map (
            O => \N__69922\,
            I => \N__69882\
        );

    \I__16966\ : Span4Mux_v
    port map (
            O => \N__69919\,
            I => \N__69879\
        );

    \I__16965\ : Sp12to4
    port map (
            O => \N__69914\,
            I => \N__69876\
        );

    \I__16964\ : Span4Mux_v
    port map (
            O => \N__69909\,
            I => \N__69873\
        );

    \I__16963\ : InMux
    port map (
            O => \N__69908\,
            I => \N__69868\
        );

    \I__16962\ : InMux
    port map (
            O => \N__69907\,
            I => \N__69868\
        );

    \I__16961\ : LocalMux
    port map (
            O => \N__69904\,
            I => \N__69863\
        );

    \I__16960\ : LocalMux
    port map (
            O => \N__69901\,
            I => \N__69863\
        );

    \I__16959\ : Span4Mux_v
    port map (
            O => \N__69898\,
            I => \N__69860\
        );

    \I__16958\ : Span4Mux_h
    port map (
            O => \N__69891\,
            I => \N__69855\
        );

    \I__16957\ : LocalMux
    port map (
            O => \N__69886\,
            I => \N__69855\
        );

    \I__16956\ : CascadeMux
    port map (
            O => \N__69885\,
            I => \N__69852\
        );

    \I__16955\ : Span4Mux_v
    port map (
            O => \N__69882\,
            I => \N__69849\
        );

    \I__16954\ : Span4Mux_h
    port map (
            O => \N__69879\,
            I => \N__69846\
        );

    \I__16953\ : Span12Mux_s9_v
    port map (
            O => \N__69876\,
            I => \N__69839\
        );

    \I__16952\ : Sp12to4
    port map (
            O => \N__69873\,
            I => \N__69839\
        );

    \I__16951\ : LocalMux
    port map (
            O => \N__69868\,
            I => \N__69839\
        );

    \I__16950\ : Span4Mux_v
    port map (
            O => \N__69863\,
            I => \N__69836\
        );

    \I__16949\ : Span4Mux_h
    port map (
            O => \N__69860\,
            I => \N__69833\
        );

    \I__16948\ : Span4Mux_h
    port map (
            O => \N__69855\,
            I => \N__69830\
        );

    \I__16947\ : InMux
    port map (
            O => \N__69852\,
            I => \N__69827\
        );

    \I__16946\ : Span4Mux_h
    port map (
            O => \N__69849\,
            I => \N__69822\
        );

    \I__16945\ : Span4Mux_h
    port map (
            O => \N__69846\,
            I => \N__69822\
        );

    \I__16944\ : Span12Mux_h
    port map (
            O => \N__69839\,
            I => \N__69819\
        );

    \I__16943\ : Span4Mux_v
    port map (
            O => \N__69836\,
            I => \N__69812\
        );

    \I__16942\ : Span4Mux_h
    port map (
            O => \N__69833\,
            I => \N__69812\
        );

    \I__16941\ : Span4Mux_v
    port map (
            O => \N__69830\,
            I => \N__69812\
        );

    \I__16940\ : LocalMux
    port map (
            O => \N__69827\,
            I => \aluOperation_4\
        );

    \I__16939\ : Odrv4
    port map (
            O => \N__69822\,
            I => \aluOperation_4\
        );

    \I__16938\ : Odrv12
    port map (
            O => \N__69819\,
            I => \aluOperation_4\
        );

    \I__16937\ : Odrv4
    port map (
            O => \N__69812\,
            I => \aluOperation_4\
        );

    \I__16936\ : CascadeMux
    port map (
            O => \N__69803\,
            I => \N__69800\
        );

    \I__16935\ : InMux
    port map (
            O => \N__69800\,
            I => \N__69791\
        );

    \I__16934\ : InMux
    port map (
            O => \N__69799\,
            I => \N__69791\
        );

    \I__16933\ : InMux
    port map (
            O => \N__69798\,
            I => \N__69791\
        );

    \I__16932\ : LocalMux
    port map (
            O => \N__69791\,
            I => \N__69786\
        );

    \I__16931\ : InMux
    port map (
            O => \N__69790\,
            I => \N__69783\
        );

    \I__16930\ : InMux
    port map (
            O => \N__69789\,
            I => \N__69780\
        );

    \I__16929\ : Span4Mux_h
    port map (
            O => \N__69786\,
            I => \N__69773\
        );

    \I__16928\ : LocalMux
    port map (
            O => \N__69783\,
            I => \N__69773\
        );

    \I__16927\ : LocalMux
    port map (
            O => \N__69780\,
            I => \N__69773\
        );

    \I__16926\ : Span4Mux_h
    port map (
            O => \N__69773\,
            I => \N__69770\
        );

    \I__16925\ : Span4Mux_h
    port map (
            O => \N__69770\,
            I => \N__69767\
        );

    \I__16924\ : Span4Mux_h
    port map (
            O => \N__69767\,
            I => \N__69763\
        );

    \I__16923\ : InMux
    port map (
            O => \N__69766\,
            I => \N__69760\
        );

    \I__16922\ : Span4Mux_h
    port map (
            O => \N__69763\,
            I => \N__69757\
        );

    \I__16921\ : LocalMux
    port map (
            O => \N__69760\,
            I => \aluOperation_3\
        );

    \I__16920\ : Odrv4
    port map (
            O => \N__69757\,
            I => \aluOperation_3\
        );

    \I__16919\ : CascadeMux
    port map (
            O => \N__69752\,
            I => \N__69749\
        );

    \I__16918\ : InMux
    port map (
            O => \N__69749\,
            I => \N__69739\
        );

    \I__16917\ : InMux
    port map (
            O => \N__69748\,
            I => \N__69739\
        );

    \I__16916\ : CascadeMux
    port map (
            O => \N__69747\,
            I => \N__69736\
        );

    \I__16915\ : CascadeMux
    port map (
            O => \N__69746\,
            I => \N__69733\
        );

    \I__16914\ : CascadeMux
    port map (
            O => \N__69745\,
            I => \N__69730\
        );

    \I__16913\ : CascadeMux
    port map (
            O => \N__69744\,
            I => \N__69726\
        );

    \I__16912\ : LocalMux
    port map (
            O => \N__69739\,
            I => \N__69723\
        );

    \I__16911\ : InMux
    port map (
            O => \N__69736\,
            I => \N__69720\
        );

    \I__16910\ : InMux
    port map (
            O => \N__69733\,
            I => \N__69717\
        );

    \I__16909\ : InMux
    port map (
            O => \N__69730\,
            I => \N__69712\
        );

    \I__16908\ : InMux
    port map (
            O => \N__69729\,
            I => \N__69707\
        );

    \I__16907\ : InMux
    port map (
            O => \N__69726\,
            I => \N__69707\
        );

    \I__16906\ : Span4Mux_v
    port map (
            O => \N__69723\,
            I => \N__69700\
        );

    \I__16905\ : LocalMux
    port map (
            O => \N__69720\,
            I => \N__69700\
        );

    \I__16904\ : LocalMux
    port map (
            O => \N__69717\,
            I => \N__69700\
        );

    \I__16903\ : CascadeMux
    port map (
            O => \N__69716\,
            I => \N__69694\
        );

    \I__16902\ : CascadeMux
    port map (
            O => \N__69715\,
            I => \N__69691\
        );

    \I__16901\ : LocalMux
    port map (
            O => \N__69712\,
            I => \N__69684\
        );

    \I__16900\ : LocalMux
    port map (
            O => \N__69707\,
            I => \N__69684\
        );

    \I__16899\ : Span4Mux_v
    port map (
            O => \N__69700\,
            I => \N__69681\
        );

    \I__16898\ : CascadeMux
    port map (
            O => \N__69699\,
            I => \N__69675\
        );

    \I__16897\ : CascadeMux
    port map (
            O => \N__69698\,
            I => \N__69672\
        );

    \I__16896\ : InMux
    port map (
            O => \N__69697\,
            I => \N__69667\
        );

    \I__16895\ : InMux
    port map (
            O => \N__69694\,
            I => \N__69667\
        );

    \I__16894\ : InMux
    port map (
            O => \N__69691\,
            I => \N__69661\
        );

    \I__16893\ : InMux
    port map (
            O => \N__69690\,
            I => \N__69661\
        );

    \I__16892\ : CascadeMux
    port map (
            O => \N__69689\,
            I => \N__69658\
        );

    \I__16891\ : Span4Mux_v
    port map (
            O => \N__69684\,
            I => \N__69655\
        );

    \I__16890\ : Span4Mux_v
    port map (
            O => \N__69681\,
            I => \N__69652\
        );

    \I__16889\ : CascadeMux
    port map (
            O => \N__69680\,
            I => \N__69648\
        );

    \I__16888\ : CascadeMux
    port map (
            O => \N__69679\,
            I => \N__69642\
        );

    \I__16887\ : CascadeMux
    port map (
            O => \N__69678\,
            I => \N__69637\
        );

    \I__16886\ : InMux
    port map (
            O => \N__69675\,
            I => \N__69634\
        );

    \I__16885\ : InMux
    port map (
            O => \N__69672\,
            I => \N__69631\
        );

    \I__16884\ : LocalMux
    port map (
            O => \N__69667\,
            I => \N__69628\
        );

    \I__16883\ : CascadeMux
    port map (
            O => \N__69666\,
            I => \N__69624\
        );

    \I__16882\ : LocalMux
    port map (
            O => \N__69661\,
            I => \N__69621\
        );

    \I__16881\ : InMux
    port map (
            O => \N__69658\,
            I => \N__69618\
        );

    \I__16880\ : Span4Mux_h
    port map (
            O => \N__69655\,
            I => \N__69613\
        );

    \I__16879\ : Span4Mux_h
    port map (
            O => \N__69652\,
            I => \N__69613\
        );

    \I__16878\ : InMux
    port map (
            O => \N__69651\,
            I => \N__69610\
        );

    \I__16877\ : InMux
    port map (
            O => \N__69648\,
            I => \N__69603\
        );

    \I__16876\ : InMux
    port map (
            O => \N__69647\,
            I => \N__69603\
        );

    \I__16875\ : InMux
    port map (
            O => \N__69646\,
            I => \N__69603\
        );

    \I__16874\ : InMux
    port map (
            O => \N__69645\,
            I => \N__69596\
        );

    \I__16873\ : InMux
    port map (
            O => \N__69642\,
            I => \N__69596\
        );

    \I__16872\ : InMux
    port map (
            O => \N__69641\,
            I => \N__69596\
        );

    \I__16871\ : InMux
    port map (
            O => \N__69640\,
            I => \N__69593\
        );

    \I__16870\ : InMux
    port map (
            O => \N__69637\,
            I => \N__69590\
        );

    \I__16869\ : LocalMux
    port map (
            O => \N__69634\,
            I => \N__69583\
        );

    \I__16868\ : LocalMux
    port map (
            O => \N__69631\,
            I => \N__69583\
        );

    \I__16867\ : Span4Mux_h
    port map (
            O => \N__69628\,
            I => \N__69583\
        );

    \I__16866\ : InMux
    port map (
            O => \N__69627\,
            I => \N__69580\
        );

    \I__16865\ : InMux
    port map (
            O => \N__69624\,
            I => \N__69577\
        );

    \I__16864\ : Span4Mux_v
    port map (
            O => \N__69621\,
            I => \N__69574\
        );

    \I__16863\ : LocalMux
    port map (
            O => \N__69618\,
            I => \N__69563\
        );

    \I__16862\ : Span4Mux_v
    port map (
            O => \N__69613\,
            I => \N__69563\
        );

    \I__16861\ : LocalMux
    port map (
            O => \N__69610\,
            I => \N__69563\
        );

    \I__16860\ : LocalMux
    port map (
            O => \N__69603\,
            I => \N__69563\
        );

    \I__16859\ : LocalMux
    port map (
            O => \N__69596\,
            I => \N__69563\
        );

    \I__16858\ : LocalMux
    port map (
            O => \N__69593\,
            I => \N__69560\
        );

    \I__16857\ : LocalMux
    port map (
            O => \N__69590\,
            I => \N__69555\
        );

    \I__16856\ : Span4Mux_h
    port map (
            O => \N__69583\,
            I => \N__69555\
        );

    \I__16855\ : LocalMux
    port map (
            O => \N__69580\,
            I => \N__69552\
        );

    \I__16854\ : LocalMux
    port map (
            O => \N__69577\,
            I => \N__69547\
        );

    \I__16853\ : Span4Mux_h
    port map (
            O => \N__69574\,
            I => \N__69547\
        );

    \I__16852\ : Span4Mux_v
    port map (
            O => \N__69563\,
            I => \N__69544\
        );

    \I__16851\ : Span4Mux_h
    port map (
            O => \N__69560\,
            I => \N__69539\
        );

    \I__16850\ : Span4Mux_v
    port map (
            O => \N__69555\,
            I => \N__69539\
        );

    \I__16849\ : Odrv12
    port map (
            O => \N__69552\,
            I => \ALU.a32Z0Z_0\
        );

    \I__16848\ : Odrv4
    port map (
            O => \N__69547\,
            I => \ALU.a32Z0Z_0\
        );

    \I__16847\ : Odrv4
    port map (
            O => \N__69544\,
            I => \ALU.a32Z0Z_0\
        );

    \I__16846\ : Odrv4
    port map (
            O => \N__69539\,
            I => \ALU.a32Z0Z_0\
        );

    \I__16845\ : InMux
    port map (
            O => \N__69530\,
            I => \N__69526\
        );

    \I__16844\ : InMux
    port map (
            O => \N__69529\,
            I => \N__69523\
        );

    \I__16843\ : LocalMux
    port map (
            O => \N__69526\,
            I => \N__69520\
        );

    \I__16842\ : LocalMux
    port map (
            O => \N__69523\,
            I => \N__69514\
        );

    \I__16841\ : Sp12to4
    port map (
            O => \N__69520\,
            I => \N__69514\
        );

    \I__16840\ : InMux
    port map (
            O => \N__69519\,
            I => \N__69509\
        );

    \I__16839\ : Span12Mux_v
    port map (
            O => \N__69514\,
            I => \N__69506\
        );

    \I__16838\ : InMux
    port map (
            O => \N__69513\,
            I => \N__69503\
        );

    \I__16837\ : InMux
    port map (
            O => \N__69512\,
            I => \N__69500\
        );

    \I__16836\ : LocalMux
    port map (
            O => \N__69509\,
            I => \N__69497\
        );

    \I__16835\ : Span12Mux_h
    port map (
            O => \N__69506\,
            I => \N__69493\
        );

    \I__16834\ : LocalMux
    port map (
            O => \N__69503\,
            I => \N__69490\
        );

    \I__16833\ : LocalMux
    port map (
            O => \N__69500\,
            I => \N__69487\
        );

    \I__16832\ : Span4Mux_h
    port map (
            O => \N__69497\,
            I => \N__69484\
        );

    \I__16831\ : CascadeMux
    port map (
            O => \N__69496\,
            I => \N__69481\
        );

    \I__16830\ : Span12Mux_v
    port map (
            O => \N__69493\,
            I => \N__69478\
        );

    \I__16829\ : Span4Mux_v
    port map (
            O => \N__69490\,
            I => \N__69473\
        );

    \I__16828\ : Span4Mux_h
    port map (
            O => \N__69487\,
            I => \N__69473\
        );

    \I__16827\ : Span4Mux_h
    port map (
            O => \N__69484\,
            I => \N__69470\
        );

    \I__16826\ : InMux
    port map (
            O => \N__69481\,
            I => \N__69467\
        );

    \I__16825\ : Odrv12
    port map (
            O => \N__69478\,
            I => \ALU.un1_operationZ0Z_7\
        );

    \I__16824\ : Odrv4
    port map (
            O => \N__69473\,
            I => \ALU.un1_operationZ0Z_7\
        );

    \I__16823\ : Odrv4
    port map (
            O => \N__69470\,
            I => \ALU.un1_operationZ0Z_7\
        );

    \I__16822\ : LocalMux
    port map (
            O => \N__69467\,
            I => \ALU.un1_operationZ0Z_7\
        );

    \I__16821\ : CEMux
    port map (
            O => \N__69458\,
            I => \N__69455\
        );

    \I__16820\ : LocalMux
    port map (
            O => \N__69455\,
            I => \N__69446\
        );

    \I__16819\ : CEMux
    port map (
            O => \N__69454\,
            I => \N__69443\
        );

    \I__16818\ : CEMux
    port map (
            O => \N__69453\,
            I => \N__69440\
        );

    \I__16817\ : CEMux
    port map (
            O => \N__69452\,
            I => \N__69437\
        );

    \I__16816\ : CEMux
    port map (
            O => \N__69451\,
            I => \N__69434\
        );

    \I__16815\ : CEMux
    port map (
            O => \N__69450\,
            I => \N__69431\
        );

    \I__16814\ : CEMux
    port map (
            O => \N__69449\,
            I => \N__69428\
        );

    \I__16813\ : Span4Mux_v
    port map (
            O => \N__69446\,
            I => \N__69425\
        );

    \I__16812\ : LocalMux
    port map (
            O => \N__69443\,
            I => \N__69422\
        );

    \I__16811\ : LocalMux
    port map (
            O => \N__69440\,
            I => \N__69419\
        );

    \I__16810\ : LocalMux
    port map (
            O => \N__69437\,
            I => \N__69416\
        );

    \I__16809\ : LocalMux
    port map (
            O => \N__69434\,
            I => \N__69413\
        );

    \I__16808\ : LocalMux
    port map (
            O => \N__69431\,
            I => \N__69408\
        );

    \I__16807\ : LocalMux
    port map (
            O => \N__69428\,
            I => \N__69408\
        );

    \I__16806\ : Span4Mux_v
    port map (
            O => \N__69425\,
            I => \N__69405\
        );

    \I__16805\ : Span4Mux_h
    port map (
            O => \N__69422\,
            I => \N__69402\
        );

    \I__16804\ : Span4Mux_h
    port map (
            O => \N__69419\,
            I => \N__69399\
        );

    \I__16803\ : Span4Mux_h
    port map (
            O => \N__69416\,
            I => \N__69396\
        );

    \I__16802\ : Span4Mux_h
    port map (
            O => \N__69413\,
            I => \N__69393\
        );

    \I__16801\ : Span4Mux_h
    port map (
            O => \N__69408\,
            I => \N__69390\
        );

    \I__16800\ : Sp12to4
    port map (
            O => \N__69405\,
            I => \N__69387\
        );

    \I__16799\ : Span4Mux_h
    port map (
            O => \N__69402\,
            I => \N__69382\
        );

    \I__16798\ : Span4Mux_h
    port map (
            O => \N__69399\,
            I => \N__69382\
        );

    \I__16797\ : Span4Mux_h
    port map (
            O => \N__69396\,
            I => \N__69379\
        );

    \I__16796\ : Span4Mux_h
    port map (
            O => \N__69393\,
            I => \N__69376\
        );

    \I__16795\ : Sp12to4
    port map (
            O => \N__69390\,
            I => \N__69373\
        );

    \I__16794\ : Span12Mux_h
    port map (
            O => \N__69387\,
            I => \N__69370\
        );

    \I__16793\ : Odrv4
    port map (
            O => \N__69382\,
            I => \ALU.un1_a41_2_0\
        );

    \I__16792\ : Odrv4
    port map (
            O => \N__69379\,
            I => \ALU.un1_a41_2_0\
        );

    \I__16791\ : Odrv4
    port map (
            O => \N__69376\,
            I => \ALU.un1_a41_2_0\
        );

    \I__16790\ : Odrv12
    port map (
            O => \N__69373\,
            I => \ALU.un1_a41_2_0\
        );

    \I__16789\ : Odrv12
    port map (
            O => \N__69370\,
            I => \ALU.un1_a41_2_0\
        );

    \I__16788\ : CascadeMux
    port map (
            O => \N__69359\,
            I => \N__69356\
        );

    \I__16787\ : InMux
    port map (
            O => \N__69356\,
            I => \N__69353\
        );

    \I__16786\ : LocalMux
    port map (
            O => \N__69353\,
            I => \N__69350\
        );

    \I__16785\ : Span4Mux_h
    port map (
            O => \N__69350\,
            I => \N__69347\
        );

    \I__16784\ : Span4Mux_h
    port map (
            O => \N__69347\,
            I => \N__69344\
        );

    \I__16783\ : Span4Mux_v
    port map (
            O => \N__69344\,
            I => \N__69341\
        );

    \I__16782\ : Odrv4
    port map (
            O => \N__69341\,
            I => \PROM.ROMDATA.m160\
        );

    \I__16781\ : CascadeMux
    port map (
            O => \N__69338\,
            I => \N__69334\
        );

    \I__16780\ : InMux
    port map (
            O => \N__69337\,
            I => \N__69324\
        );

    \I__16779\ : InMux
    port map (
            O => \N__69334\,
            I => \N__69324\
        );

    \I__16778\ : InMux
    port map (
            O => \N__69333\,
            I => \N__69324\
        );

    \I__16777\ : InMux
    port map (
            O => \N__69332\,
            I => \N__69319\
        );

    \I__16776\ : InMux
    port map (
            O => \N__69331\,
            I => \N__69319\
        );

    \I__16775\ : LocalMux
    port map (
            O => \N__69324\,
            I => \N__69312\
        );

    \I__16774\ : LocalMux
    port map (
            O => \N__69319\,
            I => \N__69312\
        );

    \I__16773\ : InMux
    port map (
            O => \N__69318\,
            I => \N__69309\
        );

    \I__16772\ : InMux
    port map (
            O => \N__69317\,
            I => \N__69306\
        );

    \I__16771\ : Span4Mux_v
    port map (
            O => \N__69312\,
            I => \N__69303\
        );

    \I__16770\ : LocalMux
    port map (
            O => \N__69309\,
            I => \N__69298\
        );

    \I__16769\ : LocalMux
    port map (
            O => \N__69306\,
            I => \N__69298\
        );

    \I__16768\ : Span4Mux_h
    port map (
            O => \N__69303\,
            I => \N__69295\
        );

    \I__16767\ : Span12Mux_v
    port map (
            O => \N__69298\,
            I => \N__69292\
        );

    \I__16766\ : Span4Mux_h
    port map (
            O => \N__69295\,
            I => \N__69289\
        );

    \I__16765\ : Odrv12
    port map (
            O => \N__69292\,
            I => \aluOperation_6\
        );

    \I__16764\ : Odrv4
    port map (
            O => \N__69289\,
            I => \aluOperation_6\
        );

    \I__16763\ : InMux
    port map (
            O => \N__69284\,
            I => \N__69276\
        );

    \I__16762\ : InMux
    port map (
            O => \N__69283\,
            I => \N__69276\
        );

    \I__16761\ : InMux
    port map (
            O => \N__69282\,
            I => \N__69271\
        );

    \I__16760\ : InMux
    port map (
            O => \N__69281\,
            I => \N__69271\
        );

    \I__16759\ : LocalMux
    port map (
            O => \N__69276\,
            I => \N__69267\
        );

    \I__16758\ : LocalMux
    port map (
            O => \N__69271\,
            I => \N__69264\
        );

    \I__16757\ : InMux
    port map (
            O => \N__69270\,
            I => \N__69261\
        );

    \I__16756\ : Span4Mux_v
    port map (
            O => \N__69267\,
            I => \N__69258\
        );

    \I__16755\ : Span4Mux_h
    port map (
            O => \N__69264\,
            I => \N__69255\
        );

    \I__16754\ : LocalMux
    port map (
            O => \N__69261\,
            I => \aluResults_0\
        );

    \I__16753\ : Odrv4
    port map (
            O => \N__69258\,
            I => \aluResults_0\
        );

    \I__16752\ : Odrv4
    port map (
            O => \N__69255\,
            I => \aluResults_0\
        );

    \I__16751\ : CascadeMux
    port map (
            O => \N__69248\,
            I => \ALU.un1_a41_3_0_1_cascade_\
        );

    \I__16750\ : CEMux
    port map (
            O => \N__69245\,
            I => \N__69240\
        );

    \I__16749\ : CEMux
    port map (
            O => \N__69244\,
            I => \N__69237\
        );

    \I__16748\ : CEMux
    port map (
            O => \N__69243\,
            I => \N__69234\
        );

    \I__16747\ : LocalMux
    port map (
            O => \N__69240\,
            I => \N__69231\
        );

    \I__16746\ : LocalMux
    port map (
            O => \N__69237\,
            I => \N__69228\
        );

    \I__16745\ : LocalMux
    port map (
            O => \N__69234\,
            I => \N__69225\
        );

    \I__16744\ : Span4Mux_h
    port map (
            O => \N__69231\,
            I => \N__69222\
        );

    \I__16743\ : Span4Mux_v
    port map (
            O => \N__69228\,
            I => \N__69219\
        );

    \I__16742\ : Span4Mux_v
    port map (
            O => \N__69225\,
            I => \N__69216\
        );

    \I__16741\ : Span4Mux_v
    port map (
            O => \N__69222\,
            I => \N__69213\
        );

    \I__16740\ : Span4Mux_h
    port map (
            O => \N__69219\,
            I => \N__69210\
        );

    \I__16739\ : Span4Mux_h
    port map (
            O => \N__69216\,
            I => \N__69207\
        );

    \I__16738\ : Span4Mux_h
    port map (
            O => \N__69213\,
            I => \N__69204\
        );

    \I__16737\ : Span4Mux_h
    port map (
            O => \N__69210\,
            I => \N__69201\
        );

    \I__16736\ : Span4Mux_h
    port map (
            O => \N__69207\,
            I => \N__69198\
        );

    \I__16735\ : Span4Mux_h
    port map (
            O => \N__69204\,
            I => \N__69195\
        );

    \I__16734\ : Odrv4
    port map (
            O => \N__69201\,
            I => \ALU.un1_a41_5_0\
        );

    \I__16733\ : Odrv4
    port map (
            O => \N__69198\,
            I => \ALU.un1_a41_5_0\
        );

    \I__16732\ : Odrv4
    port map (
            O => \N__69195\,
            I => \ALU.un1_a41_5_0\
        );

    \I__16731\ : InMux
    port map (
            O => \N__69188\,
            I => \N__69185\
        );

    \I__16730\ : LocalMux
    port map (
            O => \N__69185\,
            I => \N__69182\
        );

    \I__16729\ : Span4Mux_v
    port map (
            O => \N__69182\,
            I => \N__69179\
        );

    \I__16728\ : Odrv4
    port map (
            O => \N__69179\,
            I => \ALU.N_863\
        );

    \I__16727\ : CascadeMux
    port map (
            O => \N__69176\,
            I => \ALU.N_859_cascade_\
        );

    \I__16726\ : CascadeMux
    port map (
            O => \N__69173\,
            I => \ALU.rshift_15_ns_1_1_cascade_\
        );

    \I__16725\ : InMux
    port map (
            O => \N__69170\,
            I => \N__69165\
        );

    \I__16724\ : InMux
    port map (
            O => \N__69169\,
            I => \N__69162\
        );

    \I__16723\ : CascadeMux
    port map (
            O => \N__69168\,
            I => \N__69157\
        );

    \I__16722\ : LocalMux
    port map (
            O => \N__69165\,
            I => \N__69151\
        );

    \I__16721\ : LocalMux
    port map (
            O => \N__69162\,
            I => \N__69151\
        );

    \I__16720\ : InMux
    port map (
            O => \N__69161\,
            I => \N__69146\
        );

    \I__16719\ : InMux
    port map (
            O => \N__69160\,
            I => \N__69143\
        );

    \I__16718\ : InMux
    port map (
            O => \N__69157\,
            I => \N__69140\
        );

    \I__16717\ : InMux
    port map (
            O => \N__69156\,
            I => \N__69137\
        );

    \I__16716\ : Span4Mux_v
    port map (
            O => \N__69151\,
            I => \N__69134\
        );

    \I__16715\ : InMux
    port map (
            O => \N__69150\,
            I => \N__69131\
        );

    \I__16714\ : InMux
    port map (
            O => \N__69149\,
            I => \N__69128\
        );

    \I__16713\ : LocalMux
    port map (
            O => \N__69146\,
            I => \N__69121\
        );

    \I__16712\ : LocalMux
    port map (
            O => \N__69143\,
            I => \N__69121\
        );

    \I__16711\ : LocalMux
    port map (
            O => \N__69140\,
            I => \N__69121\
        );

    \I__16710\ : LocalMux
    port map (
            O => \N__69137\,
            I => \N__69118\
        );

    \I__16709\ : Span4Mux_h
    port map (
            O => \N__69134\,
            I => \N__69112\
        );

    \I__16708\ : LocalMux
    port map (
            O => \N__69131\,
            I => \N__69112\
        );

    \I__16707\ : LocalMux
    port map (
            O => \N__69128\,
            I => \N__69107\
        );

    \I__16706\ : Span4Mux_v
    port map (
            O => \N__69121\,
            I => \N__69107\
        );

    \I__16705\ : Span4Mux_v
    port map (
            O => \N__69118\,
            I => \N__69103\
        );

    \I__16704\ : InMux
    port map (
            O => \N__69117\,
            I => \N__69100\
        );

    \I__16703\ : Span4Mux_v
    port map (
            O => \N__69112\,
            I => \N__69095\
        );

    \I__16702\ : Span4Mux_h
    port map (
            O => \N__69107\,
            I => \N__69095\
        );

    \I__16701\ : InMux
    port map (
            O => \N__69106\,
            I => \N__69092\
        );

    \I__16700\ : Span4Mux_h
    port map (
            O => \N__69103\,
            I => \N__69089\
        );

    \I__16699\ : LocalMux
    port map (
            O => \N__69100\,
            I => \N__69084\
        );

    \I__16698\ : Span4Mux_h
    port map (
            O => \N__69095\,
            I => \N__69084\
        );

    \I__16697\ : LocalMux
    port map (
            O => \N__69092\,
            I => \ALU.a_15_m2_sZ0Z_1\
        );

    \I__16696\ : Odrv4
    port map (
            O => \N__69089\,
            I => \ALU.a_15_m2_sZ0Z_1\
        );

    \I__16695\ : Odrv4
    port map (
            O => \N__69084\,
            I => \ALU.a_15_m2_sZ0Z_1\
        );

    \I__16694\ : CascadeMux
    port map (
            O => \N__69077\,
            I => \ALU.rshift_1_cascade_\
        );

    \I__16693\ : IoInMux
    port map (
            O => \N__69074\,
            I => \N__69071\
        );

    \I__16692\ : LocalMux
    port map (
            O => \N__69071\,
            I => \N__69067\
        );

    \I__16691\ : IoInMux
    port map (
            O => \N__69070\,
            I => \N__69064\
        );

    \I__16690\ : IoSpan4Mux
    port map (
            O => \N__69067\,
            I => \N__69061\
        );

    \I__16689\ : LocalMux
    port map (
            O => \N__69064\,
            I => \N__69058\
        );

    \I__16688\ : IoSpan4Mux
    port map (
            O => \N__69061\,
            I => \N__69054\
        );

    \I__16687\ : IoSpan4Mux
    port map (
            O => \N__69058\,
            I => \N__69051\
        );

    \I__16686\ : InMux
    port map (
            O => \N__69057\,
            I => \N__69048\
        );

    \I__16685\ : Sp12to4
    port map (
            O => \N__69054\,
            I => \N__69045\
        );

    \I__16684\ : Span4Mux_s2_h
    port map (
            O => \N__69051\,
            I => \N__69042\
        );

    \I__16683\ : LocalMux
    port map (
            O => \N__69048\,
            I => \N__69039\
        );

    \I__16682\ : Span12Mux_s7_h
    port map (
            O => \N__69045\,
            I => \N__69036\
        );

    \I__16681\ : Sp12to4
    port map (
            O => \N__69042\,
            I => \N__69033\
        );

    \I__16680\ : Span4Mux_v
    port map (
            O => \N__69039\,
            I => \N__69030\
        );

    \I__16679\ : Span12Mux_h
    port map (
            O => \N__69036\,
            I => \N__69027\
        );

    \I__16678\ : Span12Mux_v
    port map (
            O => \N__69033\,
            I => \N__69024\
        );

    \I__16677\ : Sp12to4
    port map (
            O => \N__69030\,
            I => \N__69021\
        );

    \I__16676\ : Odrv12
    port map (
            O => \N__69027\,
            I => bus_1
        );

    \I__16675\ : Odrv12
    port map (
            O => \N__69024\,
            I => bus_1
        );

    \I__16674\ : Odrv12
    port map (
            O => \N__69021\,
            I => bus_1
        );

    \I__16673\ : InMux
    port map (
            O => \N__69014\,
            I => \N__69006\
        );

    \I__16672\ : InMux
    port map (
            O => \N__69013\,
            I => \N__69003\
        );

    \I__16671\ : InMux
    port map (
            O => \N__69012\,
            I => \N__68999\
        );

    \I__16670\ : InMux
    port map (
            O => \N__69011\,
            I => \N__68996\
        );

    \I__16669\ : InMux
    port map (
            O => \N__69010\,
            I => \N__68993\
        );

    \I__16668\ : InMux
    port map (
            O => \N__69009\,
            I => \N__68990\
        );

    \I__16667\ : LocalMux
    port map (
            O => \N__69006\,
            I => \N__68986\
        );

    \I__16666\ : LocalMux
    port map (
            O => \N__69003\,
            I => \N__68983\
        );

    \I__16665\ : InMux
    port map (
            O => \N__69002\,
            I => \N__68980\
        );

    \I__16664\ : LocalMux
    port map (
            O => \N__68999\,
            I => \N__68977\
        );

    \I__16663\ : LocalMux
    port map (
            O => \N__68996\,
            I => \N__68970\
        );

    \I__16662\ : LocalMux
    port map (
            O => \N__68993\,
            I => \N__68970\
        );

    \I__16661\ : LocalMux
    port map (
            O => \N__68990\,
            I => \N__68970\
        );

    \I__16660\ : InMux
    port map (
            O => \N__68989\,
            I => \N__68967\
        );

    \I__16659\ : Span4Mux_v
    port map (
            O => \N__68986\,
            I => \N__68962\
        );

    \I__16658\ : Span4Mux_v
    port map (
            O => \N__68983\,
            I => \N__68962\
        );

    \I__16657\ : LocalMux
    port map (
            O => \N__68980\,
            I => \N__68955\
        );

    \I__16656\ : Span4Mux_v
    port map (
            O => \N__68977\,
            I => \N__68955\
        );

    \I__16655\ : Span4Mux_v
    port map (
            O => \N__68970\,
            I => \N__68955\
        );

    \I__16654\ : LocalMux
    port map (
            O => \N__68967\,
            I => \N__68950\
        );

    \I__16653\ : Span4Mux_h
    port map (
            O => \N__68962\,
            I => \N__68950\
        );

    \I__16652\ : Odrv4
    port map (
            O => \N__68955\,
            I => \ALU.c_RNI98D92DZ0Z_15\
        );

    \I__16651\ : Odrv4
    port map (
            O => \N__68950\,
            I => \ALU.c_RNI98D92DZ0Z_15\
        );

    \I__16650\ : InMux
    port map (
            O => \N__68945\,
            I => \N__68936\
        );

    \I__16649\ : InMux
    port map (
            O => \N__68944\,
            I => \N__68914\
        );

    \I__16648\ : InMux
    port map (
            O => \N__68943\,
            I => \N__68911\
        );

    \I__16647\ : InMux
    port map (
            O => \N__68942\,
            I => \N__68901\
        );

    \I__16646\ : InMux
    port map (
            O => \N__68941\,
            I => \N__68901\
        );

    \I__16645\ : InMux
    port map (
            O => \N__68940\,
            I => \N__68901\
        );

    \I__16644\ : InMux
    port map (
            O => \N__68939\,
            I => \N__68898\
        );

    \I__16643\ : LocalMux
    port map (
            O => \N__68936\,
            I => \N__68891\
        );

    \I__16642\ : InMux
    port map (
            O => \N__68935\,
            I => \N__68886\
        );

    \I__16641\ : InMux
    port map (
            O => \N__68934\,
            I => \N__68886\
        );

    \I__16640\ : InMux
    port map (
            O => \N__68933\,
            I => \N__68883\
        );

    \I__16639\ : CascadeMux
    port map (
            O => \N__68932\,
            I => \N__68880\
        );

    \I__16638\ : InMux
    port map (
            O => \N__68931\,
            I => \N__68875\
        );

    \I__16637\ : InMux
    port map (
            O => \N__68930\,
            I => \N__68875\
        );

    \I__16636\ : InMux
    port map (
            O => \N__68929\,
            I => \N__68872\
        );

    \I__16635\ : InMux
    port map (
            O => \N__68928\,
            I => \N__68867\
        );

    \I__16634\ : InMux
    port map (
            O => \N__68927\,
            I => \N__68867\
        );

    \I__16633\ : InMux
    port map (
            O => \N__68926\,
            I => \N__68860\
        );

    \I__16632\ : InMux
    port map (
            O => \N__68925\,
            I => \N__68860\
        );

    \I__16631\ : InMux
    port map (
            O => \N__68924\,
            I => \N__68860\
        );

    \I__16630\ : InMux
    port map (
            O => \N__68923\,
            I => \N__68855\
        );

    \I__16629\ : InMux
    port map (
            O => \N__68922\,
            I => \N__68855\
        );

    \I__16628\ : InMux
    port map (
            O => \N__68921\,
            I => \N__68852\
        );

    \I__16627\ : InMux
    port map (
            O => \N__68920\,
            I => \N__68847\
        );

    \I__16626\ : InMux
    port map (
            O => \N__68919\,
            I => \N__68847\
        );

    \I__16625\ : InMux
    port map (
            O => \N__68918\,
            I => \N__68836\
        );

    \I__16624\ : InMux
    port map (
            O => \N__68917\,
            I => \N__68836\
        );

    \I__16623\ : LocalMux
    port map (
            O => \N__68914\,
            I => \N__68831\
        );

    \I__16622\ : LocalMux
    port map (
            O => \N__68911\,
            I => \N__68831\
        );

    \I__16621\ : InMux
    port map (
            O => \N__68910\,
            I => \N__68826\
        );

    \I__16620\ : InMux
    port map (
            O => \N__68909\,
            I => \N__68826\
        );

    \I__16619\ : CascadeMux
    port map (
            O => \N__68908\,
            I => \N__68819\
        );

    \I__16618\ : LocalMux
    port map (
            O => \N__68901\,
            I => \N__68816\
        );

    \I__16617\ : LocalMux
    port map (
            O => \N__68898\,
            I => \N__68813\
        );

    \I__16616\ : InMux
    port map (
            O => \N__68897\,
            I => \N__68804\
        );

    \I__16615\ : InMux
    port map (
            O => \N__68896\,
            I => \N__68804\
        );

    \I__16614\ : InMux
    port map (
            O => \N__68895\,
            I => \N__68799\
        );

    \I__16613\ : InMux
    port map (
            O => \N__68894\,
            I => \N__68799\
        );

    \I__16612\ : Span4Mux_v
    port map (
            O => \N__68891\,
            I => \N__68796\
        );

    \I__16611\ : LocalMux
    port map (
            O => \N__68886\,
            I => \N__68791\
        );

    \I__16610\ : LocalMux
    port map (
            O => \N__68883\,
            I => \N__68791\
        );

    \I__16609\ : InMux
    port map (
            O => \N__68880\,
            I => \N__68786\
        );

    \I__16608\ : LocalMux
    port map (
            O => \N__68875\,
            I => \N__68783\
        );

    \I__16607\ : LocalMux
    port map (
            O => \N__68872\,
            I => \N__68774\
        );

    \I__16606\ : LocalMux
    port map (
            O => \N__68867\,
            I => \N__68774\
        );

    \I__16605\ : LocalMux
    port map (
            O => \N__68860\,
            I => \N__68774\
        );

    \I__16604\ : LocalMux
    port map (
            O => \N__68855\,
            I => \N__68774\
        );

    \I__16603\ : LocalMux
    port map (
            O => \N__68852\,
            I => \N__68769\
        );

    \I__16602\ : LocalMux
    port map (
            O => \N__68847\,
            I => \N__68769\
        );

    \I__16601\ : InMux
    port map (
            O => \N__68846\,
            I => \N__68762\
        );

    \I__16600\ : InMux
    port map (
            O => \N__68845\,
            I => \N__68762\
        );

    \I__16599\ : InMux
    port map (
            O => \N__68844\,
            I => \N__68762\
        );

    \I__16598\ : InMux
    port map (
            O => \N__68843\,
            I => \N__68755\
        );

    \I__16597\ : InMux
    port map (
            O => \N__68842\,
            I => \N__68755\
        );

    \I__16596\ : InMux
    port map (
            O => \N__68841\,
            I => \N__68755\
        );

    \I__16595\ : LocalMux
    port map (
            O => \N__68836\,
            I => \N__68752\
        );

    \I__16594\ : Span4Mux_h
    port map (
            O => \N__68831\,
            I => \N__68747\
        );

    \I__16593\ : LocalMux
    port map (
            O => \N__68826\,
            I => \N__68747\
        );

    \I__16592\ : InMux
    port map (
            O => \N__68825\,
            I => \N__68741\
        );

    \I__16591\ : InMux
    port map (
            O => \N__68824\,
            I => \N__68734\
        );

    \I__16590\ : InMux
    port map (
            O => \N__68823\,
            I => \N__68734\
        );

    \I__16589\ : InMux
    port map (
            O => \N__68822\,
            I => \N__68734\
        );

    \I__16588\ : InMux
    port map (
            O => \N__68819\,
            I => \N__68730\
        );

    \I__16587\ : Span4Mux_v
    port map (
            O => \N__68816\,
            I => \N__68722\
        );

    \I__16586\ : Span4Mux_h
    port map (
            O => \N__68813\,
            I => \N__68722\
        );

    \I__16585\ : InMux
    port map (
            O => \N__68812\,
            I => \N__68712\
        );

    \I__16584\ : InMux
    port map (
            O => \N__68811\,
            I => \N__68712\
        );

    \I__16583\ : InMux
    port map (
            O => \N__68810\,
            I => \N__68712\
        );

    \I__16582\ : InMux
    port map (
            O => \N__68809\,
            I => \N__68709\
        );

    \I__16581\ : LocalMux
    port map (
            O => \N__68804\,
            I => \N__68706\
        );

    \I__16580\ : LocalMux
    port map (
            O => \N__68799\,
            I => \N__68703\
        );

    \I__16579\ : Span4Mux_v
    port map (
            O => \N__68796\,
            I => \N__68698\
        );

    \I__16578\ : Span4Mux_v
    port map (
            O => \N__68791\,
            I => \N__68698\
        );

    \I__16577\ : InMux
    port map (
            O => \N__68790\,
            I => \N__68693\
        );

    \I__16576\ : InMux
    port map (
            O => \N__68789\,
            I => \N__68693\
        );

    \I__16575\ : LocalMux
    port map (
            O => \N__68786\,
            I => \N__68690\
        );

    \I__16574\ : Span4Mux_v
    port map (
            O => \N__68783\,
            I => \N__68679\
        );

    \I__16573\ : Span4Mux_h
    port map (
            O => \N__68774\,
            I => \N__68679\
        );

    \I__16572\ : Span4Mux_v
    port map (
            O => \N__68769\,
            I => \N__68679\
        );

    \I__16571\ : LocalMux
    port map (
            O => \N__68762\,
            I => \N__68679\
        );

    \I__16570\ : LocalMux
    port map (
            O => \N__68755\,
            I => \N__68679\
        );

    \I__16569\ : Span4Mux_h
    port map (
            O => \N__68752\,
            I => \N__68674\
        );

    \I__16568\ : Span4Mux_h
    port map (
            O => \N__68747\,
            I => \N__68674\
        );

    \I__16567\ : InMux
    port map (
            O => \N__68746\,
            I => \N__68667\
        );

    \I__16566\ : InMux
    port map (
            O => \N__68745\,
            I => \N__68667\
        );

    \I__16565\ : InMux
    port map (
            O => \N__68744\,
            I => \N__68667\
        );

    \I__16564\ : LocalMux
    port map (
            O => \N__68741\,
            I => \N__68662\
        );

    \I__16563\ : LocalMux
    port map (
            O => \N__68734\,
            I => \N__68662\
        );

    \I__16562\ : CascadeMux
    port map (
            O => \N__68733\,
            I => \N__68655\
        );

    \I__16561\ : LocalMux
    port map (
            O => \N__68730\,
            I => \N__68652\
        );

    \I__16560\ : InMux
    port map (
            O => \N__68729\,
            I => \N__68649\
        );

    \I__16559\ : InMux
    port map (
            O => \N__68728\,
            I => \N__68646\
        );

    \I__16558\ : InMux
    port map (
            O => \N__68727\,
            I => \N__68643\
        );

    \I__16557\ : Span4Mux_v
    port map (
            O => \N__68722\,
            I => \N__68640\
        );

    \I__16556\ : InMux
    port map (
            O => \N__68721\,
            I => \N__68637\
        );

    \I__16555\ : InMux
    port map (
            O => \N__68720\,
            I => \N__68632\
        );

    \I__16554\ : InMux
    port map (
            O => \N__68719\,
            I => \N__68632\
        );

    \I__16553\ : LocalMux
    port map (
            O => \N__68712\,
            I => \N__68619\
        );

    \I__16552\ : LocalMux
    port map (
            O => \N__68709\,
            I => \N__68619\
        );

    \I__16551\ : Span12Mux_s11_h
    port map (
            O => \N__68706\,
            I => \N__68619\
        );

    \I__16550\ : Span12Mux_v
    port map (
            O => \N__68703\,
            I => \N__68619\
        );

    \I__16549\ : Sp12to4
    port map (
            O => \N__68698\,
            I => \N__68619\
        );

    \I__16548\ : LocalMux
    port map (
            O => \N__68693\,
            I => \N__68619\
        );

    \I__16547\ : Span4Mux_v
    port map (
            O => \N__68690\,
            I => \N__68614\
        );

    \I__16546\ : Span4Mux_h
    port map (
            O => \N__68679\,
            I => \N__68614\
        );

    \I__16545\ : Span4Mux_h
    port map (
            O => \N__68674\,
            I => \N__68607\
        );

    \I__16544\ : LocalMux
    port map (
            O => \N__68667\,
            I => \N__68607\
        );

    \I__16543\ : Span4Mux_h
    port map (
            O => \N__68662\,
            I => \N__68607\
        );

    \I__16542\ : InMux
    port map (
            O => \N__68661\,
            I => \N__68600\
        );

    \I__16541\ : InMux
    port map (
            O => \N__68660\,
            I => \N__68600\
        );

    \I__16540\ : InMux
    port map (
            O => \N__68659\,
            I => \N__68600\
        );

    \I__16539\ : InMux
    port map (
            O => \N__68658\,
            I => \N__68595\
        );

    \I__16538\ : InMux
    port map (
            O => \N__68655\,
            I => \N__68595\
        );

    \I__16537\ : Span4Mux_h
    port map (
            O => \N__68652\,
            I => \N__68588\
        );

    \I__16536\ : LocalMux
    port map (
            O => \N__68649\,
            I => \N__68588\
        );

    \I__16535\ : LocalMux
    port map (
            O => \N__68646\,
            I => \N__68588\
        );

    \I__16534\ : LocalMux
    port map (
            O => \N__68643\,
            I => \ALU.status_19_1\
        );

    \I__16533\ : Odrv4
    port map (
            O => \N__68640\,
            I => \ALU.status_19_1\
        );

    \I__16532\ : LocalMux
    port map (
            O => \N__68637\,
            I => \ALU.status_19_1\
        );

    \I__16531\ : LocalMux
    port map (
            O => \N__68632\,
            I => \ALU.status_19_1\
        );

    \I__16530\ : Odrv12
    port map (
            O => \N__68619\,
            I => \ALU.status_19_1\
        );

    \I__16529\ : Odrv4
    port map (
            O => \N__68614\,
            I => \ALU.status_19_1\
        );

    \I__16528\ : Odrv4
    port map (
            O => \N__68607\,
            I => \ALU.status_19_1\
        );

    \I__16527\ : LocalMux
    port map (
            O => \N__68600\,
            I => \ALU.status_19_1\
        );

    \I__16526\ : LocalMux
    port map (
            O => \N__68595\,
            I => \ALU.status_19_1\
        );

    \I__16525\ : Odrv4
    port map (
            O => \N__68588\,
            I => \ALU.status_19_1\
        );

    \I__16524\ : InMux
    port map (
            O => \N__68567\,
            I => \N__68560\
        );

    \I__16523\ : InMux
    port map (
            O => \N__68566\,
            I => \N__68560\
        );

    \I__16522\ : InMux
    port map (
            O => \N__68565\,
            I => \N__68557\
        );

    \I__16521\ : LocalMux
    port map (
            O => \N__68560\,
            I => \N__68553\
        );

    \I__16520\ : LocalMux
    port map (
            O => \N__68557\,
            I => \N__68550\
        );

    \I__16519\ : CascadeMux
    port map (
            O => \N__68556\,
            I => \N__68547\
        );

    \I__16518\ : Span4Mux_v
    port map (
            O => \N__68553\,
            I => \N__68544\
        );

    \I__16517\ : Span4Mux_v
    port map (
            O => \N__68550\,
            I => \N__68541\
        );

    \I__16516\ : InMux
    port map (
            O => \N__68547\,
            I => \N__68538\
        );

    \I__16515\ : Odrv4
    port map (
            O => \N__68544\,
            I => \ALU.N_968\
        );

    \I__16514\ : Odrv4
    port map (
            O => \N__68541\,
            I => \ALU.N_968\
        );

    \I__16513\ : LocalMux
    port map (
            O => \N__68538\,
            I => \ALU.N_968\
        );

    \I__16512\ : CascadeMux
    port map (
            O => \N__68531\,
            I => \N__68518\
        );

    \I__16511\ : CascadeMux
    port map (
            O => \N__68530\,
            I => \N__68512\
        );

    \I__16510\ : InMux
    port map (
            O => \N__68529\,
            I => \N__68502\
        );

    \I__16509\ : InMux
    port map (
            O => \N__68528\,
            I => \N__68499\
        );

    \I__16508\ : InMux
    port map (
            O => \N__68527\,
            I => \N__68494\
        );

    \I__16507\ : InMux
    port map (
            O => \N__68526\,
            I => \N__68494\
        );

    \I__16506\ : InMux
    port map (
            O => \N__68525\,
            I => \N__68491\
        );

    \I__16505\ : InMux
    port map (
            O => \N__68524\,
            I => \N__68485\
        );

    \I__16504\ : InMux
    port map (
            O => \N__68523\,
            I => \N__68485\
        );

    \I__16503\ : InMux
    port map (
            O => \N__68522\,
            I => \N__68472\
        );

    \I__16502\ : InMux
    port map (
            O => \N__68521\,
            I => \N__68472\
        );

    \I__16501\ : InMux
    port map (
            O => \N__68518\,
            I => \N__68472\
        );

    \I__16500\ : CascadeMux
    port map (
            O => \N__68517\,
            I => \N__68469\
        );

    \I__16499\ : InMux
    port map (
            O => \N__68516\,
            I => \N__68465\
        );

    \I__16498\ : InMux
    port map (
            O => \N__68515\,
            I => \N__68461\
        );

    \I__16497\ : InMux
    port map (
            O => \N__68512\,
            I => \N__68455\
        );

    \I__16496\ : InMux
    port map (
            O => \N__68511\,
            I => \N__68452\
        );

    \I__16495\ : InMux
    port map (
            O => \N__68510\,
            I => \N__68445\
        );

    \I__16494\ : InMux
    port map (
            O => \N__68509\,
            I => \N__68445\
        );

    \I__16493\ : InMux
    port map (
            O => \N__68508\,
            I => \N__68445\
        );

    \I__16492\ : InMux
    port map (
            O => \N__68507\,
            I => \N__68442\
        );

    \I__16491\ : CascadeMux
    port map (
            O => \N__68506\,
            I => \N__68435\
        );

    \I__16490\ : CascadeMux
    port map (
            O => \N__68505\,
            I => \N__68432\
        );

    \I__16489\ : LocalMux
    port map (
            O => \N__68502\,
            I => \N__68426\
        );

    \I__16488\ : LocalMux
    port map (
            O => \N__68499\,
            I => \N__68426\
        );

    \I__16487\ : LocalMux
    port map (
            O => \N__68494\,
            I => \N__68423\
        );

    \I__16486\ : LocalMux
    port map (
            O => \N__68491\,
            I => \N__68420\
        );

    \I__16485\ : InMux
    port map (
            O => \N__68490\,
            I => \N__68417\
        );

    \I__16484\ : LocalMux
    port map (
            O => \N__68485\,
            I => \N__68414\
        );

    \I__16483\ : InMux
    port map (
            O => \N__68484\,
            I => \N__68411\
        );

    \I__16482\ : InMux
    port map (
            O => \N__68483\,
            I => \N__68404\
        );

    \I__16481\ : InMux
    port map (
            O => \N__68482\,
            I => \N__68404\
        );

    \I__16480\ : InMux
    port map (
            O => \N__68481\,
            I => \N__68404\
        );

    \I__16479\ : InMux
    port map (
            O => \N__68480\,
            I => \N__68399\
        );

    \I__16478\ : InMux
    port map (
            O => \N__68479\,
            I => \N__68399\
        );

    \I__16477\ : LocalMux
    port map (
            O => \N__68472\,
            I => \N__68396\
        );

    \I__16476\ : InMux
    port map (
            O => \N__68469\,
            I => \N__68391\
        );

    \I__16475\ : InMux
    port map (
            O => \N__68468\,
            I => \N__68388\
        );

    \I__16474\ : LocalMux
    port map (
            O => \N__68465\,
            I => \N__68385\
        );

    \I__16473\ : InMux
    port map (
            O => \N__68464\,
            I => \N__68382\
        );

    \I__16472\ : LocalMux
    port map (
            O => \N__68461\,
            I => \N__68379\
        );

    \I__16471\ : CascadeMux
    port map (
            O => \N__68460\,
            I => \N__68375\
        );

    \I__16470\ : InMux
    port map (
            O => \N__68459\,
            I => \N__68371\
        );

    \I__16469\ : InMux
    port map (
            O => \N__68458\,
            I => \N__68368\
        );

    \I__16468\ : LocalMux
    port map (
            O => \N__68455\,
            I => \N__68359\
        );

    \I__16467\ : LocalMux
    port map (
            O => \N__68452\,
            I => \N__68359\
        );

    \I__16466\ : LocalMux
    port map (
            O => \N__68445\,
            I => \N__68359\
        );

    \I__16465\ : LocalMux
    port map (
            O => \N__68442\,
            I => \N__68359\
        );

    \I__16464\ : InMux
    port map (
            O => \N__68441\,
            I => \N__68352\
        );

    \I__16463\ : InMux
    port map (
            O => \N__68440\,
            I => \N__68352\
        );

    \I__16462\ : InMux
    port map (
            O => \N__68439\,
            I => \N__68352\
        );

    \I__16461\ : InMux
    port map (
            O => \N__68438\,
            I => \N__68349\
        );

    \I__16460\ : InMux
    port map (
            O => \N__68435\,
            I => \N__68346\
        );

    \I__16459\ : InMux
    port map (
            O => \N__68432\,
            I => \N__68343\
        );

    \I__16458\ : InMux
    port map (
            O => \N__68431\,
            I => \N__68340\
        );

    \I__16457\ : Span4Mux_v
    port map (
            O => \N__68426\,
            I => \N__68329\
        );

    \I__16456\ : Span4Mux_v
    port map (
            O => \N__68423\,
            I => \N__68329\
        );

    \I__16455\ : Span4Mux_v
    port map (
            O => \N__68420\,
            I => \N__68329\
        );

    \I__16454\ : LocalMux
    port map (
            O => \N__68417\,
            I => \N__68329\
        );

    \I__16453\ : Span4Mux_v
    port map (
            O => \N__68414\,
            I => \N__68329\
        );

    \I__16452\ : LocalMux
    port map (
            O => \N__68411\,
            I => \N__68322\
        );

    \I__16451\ : LocalMux
    port map (
            O => \N__68404\,
            I => \N__68322\
        );

    \I__16450\ : LocalMux
    port map (
            O => \N__68399\,
            I => \N__68322\
        );

    \I__16449\ : Span4Mux_v
    port map (
            O => \N__68396\,
            I => \N__68319\
        );

    \I__16448\ : InMux
    port map (
            O => \N__68395\,
            I => \N__68316\
        );

    \I__16447\ : CascadeMux
    port map (
            O => \N__68394\,
            I => \N__68312\
        );

    \I__16446\ : LocalMux
    port map (
            O => \N__68391\,
            I => \N__68309\
        );

    \I__16445\ : LocalMux
    port map (
            O => \N__68388\,
            I => \N__68306\
        );

    \I__16444\ : Span4Mux_v
    port map (
            O => \N__68385\,
            I => \N__68299\
        );

    \I__16443\ : LocalMux
    port map (
            O => \N__68382\,
            I => \N__68299\
        );

    \I__16442\ : Span4Mux_h
    port map (
            O => \N__68379\,
            I => \N__68299\
        );

    \I__16441\ : InMux
    port map (
            O => \N__68378\,
            I => \N__68292\
        );

    \I__16440\ : InMux
    port map (
            O => \N__68375\,
            I => \N__68292\
        );

    \I__16439\ : InMux
    port map (
            O => \N__68374\,
            I => \N__68292\
        );

    \I__16438\ : LocalMux
    port map (
            O => \N__68371\,
            I => \N__68285\
        );

    \I__16437\ : LocalMux
    port map (
            O => \N__68368\,
            I => \N__68285\
        );

    \I__16436\ : Span4Mux_v
    port map (
            O => \N__68359\,
            I => \N__68285\
        );

    \I__16435\ : LocalMux
    port map (
            O => \N__68352\,
            I => \N__68282\
        );

    \I__16434\ : LocalMux
    port map (
            O => \N__68349\,
            I => \N__68271\
        );

    \I__16433\ : LocalMux
    port map (
            O => \N__68346\,
            I => \N__68271\
        );

    \I__16432\ : LocalMux
    port map (
            O => \N__68343\,
            I => \N__68271\
        );

    \I__16431\ : LocalMux
    port map (
            O => \N__68340\,
            I => \N__68271\
        );

    \I__16430\ : Sp12to4
    port map (
            O => \N__68329\,
            I => \N__68267\
        );

    \I__16429\ : Span4Mux_v
    port map (
            O => \N__68322\,
            I => \N__68260\
        );

    \I__16428\ : Span4Mux_h
    port map (
            O => \N__68319\,
            I => \N__68260\
        );

    \I__16427\ : LocalMux
    port map (
            O => \N__68316\,
            I => \N__68260\
        );

    \I__16426\ : InMux
    port map (
            O => \N__68315\,
            I => \N__68257\
        );

    \I__16425\ : InMux
    port map (
            O => \N__68312\,
            I => \N__68253\
        );

    \I__16424\ : Span4Mux_h
    port map (
            O => \N__68309\,
            I => \N__68240\
        );

    \I__16423\ : Span4Mux_v
    port map (
            O => \N__68306\,
            I => \N__68240\
        );

    \I__16422\ : Span4Mux_v
    port map (
            O => \N__68299\,
            I => \N__68240\
        );

    \I__16421\ : LocalMux
    port map (
            O => \N__68292\,
            I => \N__68240\
        );

    \I__16420\ : Span4Mux_h
    port map (
            O => \N__68285\,
            I => \N__68240\
        );

    \I__16419\ : Span4Mux_h
    port map (
            O => \N__68282\,
            I => \N__68240\
        );

    \I__16418\ : InMux
    port map (
            O => \N__68281\,
            I => \N__68237\
        );

    \I__16417\ : CascadeMux
    port map (
            O => \N__68280\,
            I => \N__68234\
        );

    \I__16416\ : Span4Mux_v
    port map (
            O => \N__68271\,
            I => \N__68225\
        );

    \I__16415\ : InMux
    port map (
            O => \N__68270\,
            I => \N__68222\
        );

    \I__16414\ : Span12Mux_h
    port map (
            O => \N__68267\,
            I => \N__68215\
        );

    \I__16413\ : Sp12to4
    port map (
            O => \N__68260\,
            I => \N__68215\
        );

    \I__16412\ : LocalMux
    port map (
            O => \N__68257\,
            I => \N__68215\
        );

    \I__16411\ : InMux
    port map (
            O => \N__68256\,
            I => \N__68212\
        );

    \I__16410\ : LocalMux
    port map (
            O => \N__68253\,
            I => \N__68205\
        );

    \I__16409\ : Span4Mux_h
    port map (
            O => \N__68240\,
            I => \N__68205\
        );

    \I__16408\ : LocalMux
    port map (
            O => \N__68237\,
            I => \N__68205\
        );

    \I__16407\ : InMux
    port map (
            O => \N__68234\,
            I => \N__68196\
        );

    \I__16406\ : InMux
    port map (
            O => \N__68233\,
            I => \N__68196\
        );

    \I__16405\ : InMux
    port map (
            O => \N__68232\,
            I => \N__68196\
        );

    \I__16404\ : InMux
    port map (
            O => \N__68231\,
            I => \N__68196\
        );

    \I__16403\ : InMux
    port map (
            O => \N__68230\,
            I => \N__68189\
        );

    \I__16402\ : InMux
    port map (
            O => \N__68229\,
            I => \N__68189\
        );

    \I__16401\ : InMux
    port map (
            O => \N__68228\,
            I => \N__68189\
        );

    \I__16400\ : Odrv4
    port map (
            O => \N__68225\,
            I => \ALU.status_19_2\
        );

    \I__16399\ : LocalMux
    port map (
            O => \N__68222\,
            I => \ALU.status_19_2\
        );

    \I__16398\ : Odrv12
    port map (
            O => \N__68215\,
            I => \ALU.status_19_2\
        );

    \I__16397\ : LocalMux
    port map (
            O => \N__68212\,
            I => \ALU.status_19_2\
        );

    \I__16396\ : Odrv4
    port map (
            O => \N__68205\,
            I => \ALU.status_19_2\
        );

    \I__16395\ : LocalMux
    port map (
            O => \N__68196\,
            I => \ALU.status_19_2\
        );

    \I__16394\ : LocalMux
    port map (
            O => \N__68189\,
            I => \ALU.status_19_2\
        );

    \I__16393\ : InMux
    port map (
            O => \N__68174\,
            I => \N__68171\
        );

    \I__16392\ : LocalMux
    port map (
            O => \N__68171\,
            I => \N__68168\
        );

    \I__16391\ : Span4Mux_v
    port map (
            O => \N__68168\,
            I => \N__68163\
        );

    \I__16390\ : InMux
    port map (
            O => \N__68167\,
            I => \N__68158\
        );

    \I__16389\ : InMux
    port map (
            O => \N__68166\,
            I => \N__68158\
        );

    \I__16388\ : Sp12to4
    port map (
            O => \N__68163\,
            I => \N__68153\
        );

    \I__16387\ : LocalMux
    port map (
            O => \N__68158\,
            I => \N__68153\
        );

    \I__16386\ : Odrv12
    port map (
            O => \N__68153\,
            I => \ALU.N_867\
        );

    \I__16385\ : InMux
    port map (
            O => \N__68150\,
            I => \N__68147\
        );

    \I__16384\ : LocalMux
    port map (
            O => \N__68147\,
            I => \ALU.c_RNICBIG85Z0Z_15\
        );

    \I__16383\ : InMux
    port map (
            O => \N__68144\,
            I => \N__68141\
        );

    \I__16382\ : LocalMux
    port map (
            O => \N__68141\,
            I => \N__68133\
        );

    \I__16381\ : InMux
    port map (
            O => \N__68140\,
            I => \N__68130\
        );

    \I__16380\ : InMux
    port map (
            O => \N__68139\,
            I => \N__68127\
        );

    \I__16379\ : InMux
    port map (
            O => \N__68138\,
            I => \N__68124\
        );

    \I__16378\ : InMux
    port map (
            O => \N__68137\,
            I => \N__68119\
        );

    \I__16377\ : InMux
    port map (
            O => \N__68136\,
            I => \N__68116\
        );

    \I__16376\ : Span4Mux_v
    port map (
            O => \N__68133\,
            I => \N__68109\
        );

    \I__16375\ : LocalMux
    port map (
            O => \N__68130\,
            I => \N__68109\
        );

    \I__16374\ : LocalMux
    port map (
            O => \N__68127\,
            I => \N__68109\
        );

    \I__16373\ : LocalMux
    port map (
            O => \N__68124\,
            I => \N__68106\
        );

    \I__16372\ : InMux
    port map (
            O => \N__68123\,
            I => \N__68103\
        );

    \I__16371\ : InMux
    port map (
            O => \N__68122\,
            I => \N__68100\
        );

    \I__16370\ : LocalMux
    port map (
            O => \N__68119\,
            I => \ALU.a_15_ns_snZ0Z_14\
        );

    \I__16369\ : LocalMux
    port map (
            O => \N__68116\,
            I => \ALU.a_15_ns_snZ0Z_14\
        );

    \I__16368\ : Odrv4
    port map (
            O => \N__68109\,
            I => \ALU.a_15_ns_snZ0Z_14\
        );

    \I__16367\ : Odrv4
    port map (
            O => \N__68106\,
            I => \ALU.a_15_ns_snZ0Z_14\
        );

    \I__16366\ : LocalMux
    port map (
            O => \N__68103\,
            I => \ALU.a_15_ns_snZ0Z_14\
        );

    \I__16365\ : LocalMux
    port map (
            O => \N__68100\,
            I => \ALU.a_15_ns_snZ0Z_14\
        );

    \I__16364\ : InMux
    port map (
            O => \N__68087\,
            I => \N__68083\
        );

    \I__16363\ : InMux
    port map (
            O => \N__68086\,
            I => \N__68080\
        );

    \I__16362\ : LocalMux
    port map (
            O => \N__68083\,
            I => \N__68071\
        );

    \I__16361\ : LocalMux
    port map (
            O => \N__68080\,
            I => \N__68071\
        );

    \I__16360\ : InMux
    port map (
            O => \N__68079\,
            I => \N__68068\
        );

    \I__16359\ : InMux
    port map (
            O => \N__68078\,
            I => \N__68065\
        );

    \I__16358\ : InMux
    port map (
            O => \N__68077\,
            I => \N__68062\
        );

    \I__16357\ : InMux
    port map (
            O => \N__68076\,
            I => \N__68059\
        );

    \I__16356\ : Span4Mux_h
    port map (
            O => \N__68071\,
            I => \N__68054\
        );

    \I__16355\ : LocalMux
    port map (
            O => \N__68068\,
            I => \N__68049\
        );

    \I__16354\ : LocalMux
    port map (
            O => \N__68065\,
            I => \N__68049\
        );

    \I__16353\ : LocalMux
    port map (
            O => \N__68062\,
            I => \N__68046\
        );

    \I__16352\ : LocalMux
    port map (
            O => \N__68059\,
            I => \N__68043\
        );

    \I__16351\ : InMux
    port map (
            O => \N__68058\,
            I => \N__68040\
        );

    \I__16350\ : InMux
    port map (
            O => \N__68057\,
            I => \N__68037\
        );

    \I__16349\ : Span4Mux_h
    port map (
            O => \N__68054\,
            I => \N__68034\
        );

    \I__16348\ : Span4Mux_v
    port map (
            O => \N__68049\,
            I => \N__68023\
        );

    \I__16347\ : Span4Mux_v
    port map (
            O => \N__68046\,
            I => \N__68023\
        );

    \I__16346\ : Span4Mux_h
    port map (
            O => \N__68043\,
            I => \N__68023\
        );

    \I__16345\ : LocalMux
    port map (
            O => \N__68040\,
            I => \N__68023\
        );

    \I__16344\ : LocalMux
    port map (
            O => \N__68037\,
            I => \N__68023\
        );

    \I__16343\ : Span4Mux_h
    port map (
            O => \N__68034\,
            I => \N__68020\
        );

    \I__16342\ : Span4Mux_h
    port map (
            O => \N__68023\,
            I => \N__68017\
        );

    \I__16341\ : Odrv4
    port map (
            O => \N__68020\,
            I => \ALU.lshift_14\
        );

    \I__16340\ : Odrv4
    port map (
            O => \N__68017\,
            I => \ALU.lshift_14\
        );

    \I__16339\ : InMux
    port map (
            O => \N__68012\,
            I => \N__68008\
        );

    \I__16338\ : InMux
    port map (
            O => \N__68011\,
            I => \N__68005\
        );

    \I__16337\ : LocalMux
    port map (
            O => \N__68008\,
            I => \N__67997\
        );

    \I__16336\ : LocalMux
    port map (
            O => \N__68005\,
            I => \N__67994\
        );

    \I__16335\ : InMux
    port map (
            O => \N__68004\,
            I => \N__67991\
        );

    \I__16334\ : InMux
    port map (
            O => \N__68003\,
            I => \N__67988\
        );

    \I__16333\ : InMux
    port map (
            O => \N__68002\,
            I => \N__67985\
        );

    \I__16332\ : InMux
    port map (
            O => \N__68001\,
            I => \N__67982\
        );

    \I__16331\ : InMux
    port map (
            O => \N__68000\,
            I => \N__67979\
        );

    \I__16330\ : Odrv4
    port map (
            O => \N__67997\,
            I => \ALU.a_15_ns_rn_0_14\
        );

    \I__16329\ : Odrv4
    port map (
            O => \N__67994\,
            I => \ALU.a_15_ns_rn_0_14\
        );

    \I__16328\ : LocalMux
    port map (
            O => \N__67991\,
            I => \ALU.a_15_ns_rn_0_14\
        );

    \I__16327\ : LocalMux
    port map (
            O => \N__67988\,
            I => \ALU.a_15_ns_rn_0_14\
        );

    \I__16326\ : LocalMux
    port map (
            O => \N__67985\,
            I => \ALU.a_15_ns_rn_0_14\
        );

    \I__16325\ : LocalMux
    port map (
            O => \N__67982\,
            I => \ALU.a_15_ns_rn_0_14\
        );

    \I__16324\ : LocalMux
    port map (
            O => \N__67979\,
            I => \ALU.a_15_ns_rn_0_14\
        );

    \I__16323\ : InMux
    port map (
            O => \N__67964\,
            I => \N__67960\
        );

    \I__16322\ : InMux
    port map (
            O => \N__67963\,
            I => \N__67957\
        );

    \I__16321\ : LocalMux
    port map (
            O => \N__67960\,
            I => \N__67952\
        );

    \I__16320\ : LocalMux
    port map (
            O => \N__67957\,
            I => \N__67952\
        );

    \I__16319\ : Span4Mux_v
    port map (
            O => \N__67952\,
            I => \N__67949\
        );

    \I__16318\ : Span4Mux_h
    port map (
            O => \N__67949\,
            I => \N__67946\
        );

    \I__16317\ : Odrv4
    port map (
            O => \N__67946\,
            I => \ALU.bZ0Z_14\
        );

    \I__16316\ : CEMux
    port map (
            O => \N__67943\,
            I => \N__67939\
        );

    \I__16315\ : CEMux
    port map (
            O => \N__67942\,
            I => \N__67935\
        );

    \I__16314\ : LocalMux
    port map (
            O => \N__67939\,
            I => \N__67932\
        );

    \I__16313\ : CEMux
    port map (
            O => \N__67938\,
            I => \N__67928\
        );

    \I__16312\ : LocalMux
    port map (
            O => \N__67935\,
            I => \N__67925\
        );

    \I__16311\ : Span4Mux_v
    port map (
            O => \N__67932\,
            I => \N__67922\
        );

    \I__16310\ : CEMux
    port map (
            O => \N__67931\,
            I => \N__67918\
        );

    \I__16309\ : LocalMux
    port map (
            O => \N__67928\,
            I => \N__67915\
        );

    \I__16308\ : Span4Mux_v
    port map (
            O => \N__67925\,
            I => \N__67912\
        );

    \I__16307\ : Span4Mux_h
    port map (
            O => \N__67922\,
            I => \N__67909\
        );

    \I__16306\ : CEMux
    port map (
            O => \N__67921\,
            I => \N__67906\
        );

    \I__16305\ : LocalMux
    port map (
            O => \N__67918\,
            I => \N__67903\
        );

    \I__16304\ : Span4Mux_h
    port map (
            O => \N__67915\,
            I => \N__67900\
        );

    \I__16303\ : Span4Mux_h
    port map (
            O => \N__67912\,
            I => \N__67897\
        );

    \I__16302\ : Span4Mux_v
    port map (
            O => \N__67909\,
            I => \N__67894\
        );

    \I__16301\ : LocalMux
    port map (
            O => \N__67906\,
            I => \N__67891\
        );

    \I__16300\ : Span4Mux_h
    port map (
            O => \N__67903\,
            I => \N__67888\
        );

    \I__16299\ : Span4Mux_h
    port map (
            O => \N__67900\,
            I => \N__67885\
        );

    \I__16298\ : Span4Mux_v
    port map (
            O => \N__67897\,
            I => \N__67880\
        );

    \I__16297\ : Span4Mux_h
    port map (
            O => \N__67894\,
            I => \N__67880\
        );

    \I__16296\ : Odrv12
    port map (
            O => \N__67891\,
            I => \ALU.un1_a41_8_0\
        );

    \I__16295\ : Odrv4
    port map (
            O => \N__67888\,
            I => \ALU.un1_a41_8_0\
        );

    \I__16294\ : Odrv4
    port map (
            O => \N__67885\,
            I => \ALU.un1_a41_8_0\
        );

    \I__16293\ : Odrv4
    port map (
            O => \N__67880\,
            I => \ALU.un1_a41_8_0\
        );

    \I__16292\ : CEMux
    port map (
            O => \N__67871\,
            I => \N__67868\
        );

    \I__16291\ : LocalMux
    port map (
            O => \N__67868\,
            I => \N__67865\
        );

    \I__16290\ : Span4Mux_v
    port map (
            O => \N__67865\,
            I => \N__67861\
        );

    \I__16289\ : CEMux
    port map (
            O => \N__67864\,
            I => \N__67857\
        );

    \I__16288\ : Span4Mux_h
    port map (
            O => \N__67861\,
            I => \N__67854\
        );

    \I__16287\ : CEMux
    port map (
            O => \N__67860\,
            I => \N__67851\
        );

    \I__16286\ : LocalMux
    port map (
            O => \N__67857\,
            I => \N__67848\
        );

    \I__16285\ : Span4Mux_h
    port map (
            O => \N__67854\,
            I => \N__67845\
        );

    \I__16284\ : LocalMux
    port map (
            O => \N__67851\,
            I => \N__67842\
        );

    \I__16283\ : Sp12to4
    port map (
            O => \N__67848\,
            I => \N__67839\
        );

    \I__16282\ : Span4Mux_h
    port map (
            O => \N__67845\,
            I => \N__67836\
        );

    \I__16281\ : Span4Mux_v
    port map (
            O => \N__67842\,
            I => \N__67833\
        );

    \I__16280\ : Span12Mux_s11_v
    port map (
            O => \N__67839\,
            I => \N__67830\
        );

    \I__16279\ : Sp12to4
    port map (
            O => \N__67836\,
            I => \N__67827\
        );

    \I__16278\ : Odrv4
    port map (
            O => \N__67833\,
            I => \ALU.un1_a41_4_0\
        );

    \I__16277\ : Odrv12
    port map (
            O => \N__67830\,
            I => \ALU.un1_a41_4_0\
        );

    \I__16276\ : Odrv12
    port map (
            O => \N__67827\,
            I => \ALU.un1_a41_4_0\
        );

    \I__16275\ : InMux
    port map (
            O => \N__67820\,
            I => \N__67817\
        );

    \I__16274\ : LocalMux
    port map (
            O => \N__67817\,
            I => \N__67814\
        );

    \I__16273\ : Span12Mux_v
    port map (
            O => \N__67814\,
            I => \N__67811\
        );

    \I__16272\ : Odrv12
    port map (
            O => \N__67811\,
            I => \ALU.un1_operation_5_0\
        );

    \I__16271\ : CascadeMux
    port map (
            O => \N__67808\,
            I => \N__67805\
        );

    \I__16270\ : InMux
    port map (
            O => \N__67805\,
            I => \N__67802\
        );

    \I__16269\ : LocalMux
    port map (
            O => \N__67802\,
            I => \N__67799\
        );

    \I__16268\ : Span4Mux_v
    port map (
            O => \N__67799\,
            I => \N__67796\
        );

    \I__16267\ : Sp12to4
    port map (
            O => \N__67796\,
            I => \N__67793\
        );

    \I__16266\ : Span12Mux_h
    port map (
            O => \N__67793\,
            I => \N__67790\
        );

    \I__16265\ : Odrv12
    port map (
            O => \N__67790\,
            I => \aluOperation_5\
        );

    \I__16264\ : CascadeMux
    port map (
            O => \N__67787\,
            I => \ALU.un1_operation_10_0_cascade_\
        );

    \I__16263\ : InMux
    port map (
            O => \N__67784\,
            I => \N__67780\
        );

    \I__16262\ : InMux
    port map (
            O => \N__67783\,
            I => \N__67777\
        );

    \I__16261\ : LocalMux
    port map (
            O => \N__67780\,
            I => \N__67774\
        );

    \I__16260\ : LocalMux
    port map (
            O => \N__67777\,
            I => \N__67771\
        );

    \I__16259\ : Span4Mux_v
    port map (
            O => \N__67774\,
            I => \N__67766\
        );

    \I__16258\ : Span4Mux_h
    port map (
            O => \N__67771\,
            I => \N__67766\
        );

    \I__16257\ : Span4Mux_h
    port map (
            O => \N__67766\,
            I => \N__67763\
        );

    \I__16256\ : Sp12to4
    port map (
            O => \N__67763\,
            I => \N__67760\
        );

    \I__16255\ : Odrv12
    port map (
            O => \N__67760\,
            I => \ALU.dZ0Z_14\
        );

    \I__16254\ : InMux
    port map (
            O => \N__67757\,
            I => \N__67750\
        );

    \I__16253\ : InMux
    port map (
            O => \N__67756\,
            I => \N__67747\
        );

    \I__16252\ : InMux
    port map (
            O => \N__67755\,
            I => \N__67744\
        );

    \I__16251\ : InMux
    port map (
            O => \N__67754\,
            I => \N__67738\
        );

    \I__16250\ : InMux
    port map (
            O => \N__67753\,
            I => \N__67735\
        );

    \I__16249\ : LocalMux
    port map (
            O => \N__67750\,
            I => \N__67732\
        );

    \I__16248\ : LocalMux
    port map (
            O => \N__67747\,
            I => \N__67729\
        );

    \I__16247\ : LocalMux
    port map (
            O => \N__67744\,
            I => \N__67726\
        );

    \I__16246\ : InMux
    port map (
            O => \N__67743\,
            I => \N__67723\
        );

    \I__16245\ : InMux
    port map (
            O => \N__67742\,
            I => \N__67720\
        );

    \I__16244\ : InMux
    port map (
            O => \N__67741\,
            I => \N__67717\
        );

    \I__16243\ : LocalMux
    port map (
            O => \N__67738\,
            I => \N__67712\
        );

    \I__16242\ : LocalMux
    port map (
            O => \N__67735\,
            I => \N__67712\
        );

    \I__16241\ : Span4Mux_h
    port map (
            O => \N__67732\,
            I => \N__67707\
        );

    \I__16240\ : Span4Mux_h
    port map (
            O => \N__67729\,
            I => \N__67707\
        );

    \I__16239\ : Span12Mux_v
    port map (
            O => \N__67726\,
            I => \N__67704\
        );

    \I__16238\ : LocalMux
    port map (
            O => \N__67723\,
            I => \ALU.c_RNIBRG4Q9Z0Z_12\
        );

    \I__16237\ : LocalMux
    port map (
            O => \N__67720\,
            I => \ALU.c_RNIBRG4Q9Z0Z_12\
        );

    \I__16236\ : LocalMux
    port map (
            O => \N__67717\,
            I => \ALU.c_RNIBRG4Q9Z0Z_12\
        );

    \I__16235\ : Odrv12
    port map (
            O => \N__67712\,
            I => \ALU.c_RNIBRG4Q9Z0Z_12\
        );

    \I__16234\ : Odrv4
    port map (
            O => \N__67707\,
            I => \ALU.c_RNIBRG4Q9Z0Z_12\
        );

    \I__16233\ : Odrv12
    port map (
            O => \N__67704\,
            I => \ALU.c_RNIBRG4Q9Z0Z_12\
        );

    \I__16232\ : InMux
    port map (
            O => \N__67691\,
            I => \N__67688\
        );

    \I__16231\ : LocalMux
    port map (
            O => \N__67688\,
            I => \N__67682\
        );

    \I__16230\ : InMux
    port map (
            O => \N__67687\,
            I => \N__67679\
        );

    \I__16229\ : InMux
    port map (
            O => \N__67686\,
            I => \N__67676\
        );

    \I__16228\ : InMux
    port map (
            O => \N__67685\,
            I => \N__67673\
        );

    \I__16227\ : Span4Mux_v
    port map (
            O => \N__67682\,
            I => \N__67669\
        );

    \I__16226\ : LocalMux
    port map (
            O => \N__67679\,
            I => \N__67665\
        );

    \I__16225\ : LocalMux
    port map (
            O => \N__67676\,
            I => \N__67662\
        );

    \I__16224\ : LocalMux
    port map (
            O => \N__67673\,
            I => \N__67659\
        );

    \I__16223\ : InMux
    port map (
            O => \N__67672\,
            I => \N__67656\
        );

    \I__16222\ : Span4Mux_h
    port map (
            O => \N__67669\,
            I => \N__67651\
        );

    \I__16221\ : InMux
    port map (
            O => \N__67668\,
            I => \N__67648\
        );

    \I__16220\ : Span4Mux_v
    port map (
            O => \N__67665\,
            I => \N__67639\
        );

    \I__16219\ : Span4Mux_v
    port map (
            O => \N__67662\,
            I => \N__67639\
        );

    \I__16218\ : Span4Mux_h
    port map (
            O => \N__67659\,
            I => \N__67639\
        );

    \I__16217\ : LocalMux
    port map (
            O => \N__67656\,
            I => \N__67639\
        );

    \I__16216\ : InMux
    port map (
            O => \N__67655\,
            I => \N__67636\
        );

    \I__16215\ : InMux
    port map (
            O => \N__67654\,
            I => \N__67633\
        );

    \I__16214\ : Odrv4
    port map (
            O => \N__67651\,
            I => \ALU.c_RNIBRG4Q9_0Z0Z_12\
        );

    \I__16213\ : LocalMux
    port map (
            O => \N__67648\,
            I => \ALU.c_RNIBRG4Q9_0Z0Z_12\
        );

    \I__16212\ : Odrv4
    port map (
            O => \N__67639\,
            I => \ALU.c_RNIBRG4Q9_0Z0Z_12\
        );

    \I__16211\ : LocalMux
    port map (
            O => \N__67636\,
            I => \ALU.c_RNIBRG4Q9_0Z0Z_12\
        );

    \I__16210\ : LocalMux
    port map (
            O => \N__67633\,
            I => \ALU.c_RNIBRG4Q9_0Z0Z_12\
        );

    \I__16209\ : CascadeMux
    port map (
            O => \N__67622\,
            I => \N__67618\
        );

    \I__16208\ : InMux
    port map (
            O => \N__67621\,
            I => \N__67614\
        );

    \I__16207\ : InMux
    port map (
            O => \N__67618\,
            I => \N__67611\
        );

    \I__16206\ : InMux
    port map (
            O => \N__67617\,
            I => \N__67607\
        );

    \I__16205\ : LocalMux
    port map (
            O => \N__67614\,
            I => \N__67604\
        );

    \I__16204\ : LocalMux
    port map (
            O => \N__67611\,
            I => \N__67599\
        );

    \I__16203\ : InMux
    port map (
            O => \N__67610\,
            I => \N__67596\
        );

    \I__16202\ : LocalMux
    port map (
            O => \N__67607\,
            I => \N__67590\
        );

    \I__16201\ : Span4Mux_v
    port map (
            O => \N__67604\,
            I => \N__67590\
        );

    \I__16200\ : InMux
    port map (
            O => \N__67603\,
            I => \N__67587\
        );

    \I__16199\ : CascadeMux
    port map (
            O => \N__67602\,
            I => \N__67584\
        );

    \I__16198\ : Span4Mux_v
    port map (
            O => \N__67599\,
            I => \N__67581\
        );

    \I__16197\ : LocalMux
    port map (
            O => \N__67596\,
            I => \N__67578\
        );

    \I__16196\ : InMux
    port map (
            O => \N__67595\,
            I => \N__67575\
        );

    \I__16195\ : Span4Mux_v
    port map (
            O => \N__67590\,
            I => \N__67570\
        );

    \I__16194\ : LocalMux
    port map (
            O => \N__67587\,
            I => \N__67570\
        );

    \I__16193\ : InMux
    port map (
            O => \N__67584\,
            I => \N__67567\
        );

    \I__16192\ : Odrv4
    port map (
            O => \N__67581\,
            I => \ALU.mult_555_c_RNIJF56AMZ0\
        );

    \I__16191\ : Odrv4
    port map (
            O => \N__67578\,
            I => \ALU.mult_555_c_RNIJF56AMZ0\
        );

    \I__16190\ : LocalMux
    port map (
            O => \N__67575\,
            I => \ALU.mult_555_c_RNIJF56AMZ0\
        );

    \I__16189\ : Odrv4
    port map (
            O => \N__67570\,
            I => \ALU.mult_555_c_RNIJF56AMZ0\
        );

    \I__16188\ : LocalMux
    port map (
            O => \N__67567\,
            I => \ALU.mult_555_c_RNIJF56AMZ0\
        );

    \I__16187\ : InMux
    port map (
            O => \N__67556\,
            I => \N__67553\
        );

    \I__16186\ : LocalMux
    port map (
            O => \N__67553\,
            I => \N__67550\
        );

    \I__16185\ : Span4Mux_v
    port map (
            O => \N__67550\,
            I => \N__67546\
        );

    \I__16184\ : InMux
    port map (
            O => \N__67549\,
            I => \N__67543\
        );

    \I__16183\ : Span4Mux_h
    port map (
            O => \N__67546\,
            I => \N__67538\
        );

    \I__16182\ : LocalMux
    port map (
            O => \N__67543\,
            I => \N__67538\
        );

    \I__16181\ : Span4Mux_h
    port map (
            O => \N__67538\,
            I => \N__67535\
        );

    \I__16180\ : Span4Mux_h
    port map (
            O => \N__67535\,
            I => \N__67532\
        );

    \I__16179\ : Span4Mux_h
    port map (
            O => \N__67532\,
            I => \N__67529\
        );

    \I__16178\ : Span4Mux_h
    port map (
            O => \N__67529\,
            I => \N__67526\
        );

    \I__16177\ : Span4Mux_v
    port map (
            O => \N__67526\,
            I => \N__67523\
        );

    \I__16176\ : Span4Mux_h
    port map (
            O => \N__67523\,
            I => \N__67520\
        );

    \I__16175\ : Odrv4
    port map (
            O => \N__67520\,
            I => \ALU.cZ0Z_12\
        );

    \I__16174\ : InMux
    port map (
            O => \N__67517\,
            I => \N__67513\
        );

    \I__16173\ : InMux
    port map (
            O => \N__67516\,
            I => \N__67509\
        );

    \I__16172\ : LocalMux
    port map (
            O => \N__67513\,
            I => \N__67505\
        );

    \I__16171\ : InMux
    port map (
            O => \N__67512\,
            I => \N__67501\
        );

    \I__16170\ : LocalMux
    port map (
            O => \N__67509\,
            I => \N__67498\
        );

    \I__16169\ : InMux
    port map (
            O => \N__67508\,
            I => \N__67495\
        );

    \I__16168\ : Span4Mux_v
    port map (
            O => \N__67505\,
            I => \N__67490\
        );

    \I__16167\ : InMux
    port map (
            O => \N__67504\,
            I => \N__67487\
        );

    \I__16166\ : LocalMux
    port map (
            O => \N__67501\,
            I => \N__67484\
        );

    \I__16165\ : Span4Mux_v
    port map (
            O => \N__67498\,
            I => \N__67479\
        );

    \I__16164\ : LocalMux
    port map (
            O => \N__67495\,
            I => \N__67479\
        );

    \I__16163\ : InMux
    port map (
            O => \N__67494\,
            I => \N__67476\
        );

    \I__16162\ : InMux
    port map (
            O => \N__67493\,
            I => \N__67473\
        );

    \I__16161\ : Odrv4
    port map (
            O => \N__67490\,
            I => \ALU.c_RNIO5N04A_0Z0Z_13\
        );

    \I__16160\ : LocalMux
    port map (
            O => \N__67487\,
            I => \ALU.c_RNIO5N04A_0Z0Z_13\
        );

    \I__16159\ : Odrv4
    port map (
            O => \N__67484\,
            I => \ALU.c_RNIO5N04A_0Z0Z_13\
        );

    \I__16158\ : Odrv4
    port map (
            O => \N__67479\,
            I => \ALU.c_RNIO5N04A_0Z0Z_13\
        );

    \I__16157\ : LocalMux
    port map (
            O => \N__67476\,
            I => \ALU.c_RNIO5N04A_0Z0Z_13\
        );

    \I__16156\ : LocalMux
    port map (
            O => \N__67473\,
            I => \ALU.c_RNIO5N04A_0Z0Z_13\
        );

    \I__16155\ : InMux
    port map (
            O => \N__67460\,
            I => \N__67456\
        );

    \I__16154\ : InMux
    port map (
            O => \N__67459\,
            I => \N__67452\
        );

    \I__16153\ : LocalMux
    port map (
            O => \N__67456\,
            I => \N__67446\
        );

    \I__16152\ : InMux
    port map (
            O => \N__67455\,
            I => \N__67443\
        );

    \I__16151\ : LocalMux
    port map (
            O => \N__67452\,
            I => \N__67439\
        );

    \I__16150\ : InMux
    port map (
            O => \N__67451\,
            I => \N__67436\
        );

    \I__16149\ : InMux
    port map (
            O => \N__67450\,
            I => \N__67433\
        );

    \I__16148\ : InMux
    port map (
            O => \N__67449\,
            I => \N__67429\
        );

    \I__16147\ : Span4Mux_h
    port map (
            O => \N__67446\,
            I => \N__67424\
        );

    \I__16146\ : LocalMux
    port map (
            O => \N__67443\,
            I => \N__67424\
        );

    \I__16145\ : InMux
    port map (
            O => \N__67442\,
            I => \N__67421\
        );

    \I__16144\ : Span4Mux_v
    port map (
            O => \N__67439\,
            I => \N__67414\
        );

    \I__16143\ : LocalMux
    port map (
            O => \N__67436\,
            I => \N__67414\
        );

    \I__16142\ : LocalMux
    port map (
            O => \N__67433\,
            I => \N__67414\
        );

    \I__16141\ : InMux
    port map (
            O => \N__67432\,
            I => \N__67411\
        );

    \I__16140\ : LocalMux
    port map (
            O => \N__67429\,
            I => \ALU.c_RNIO5N04AZ0Z_13\
        );

    \I__16139\ : Odrv4
    port map (
            O => \N__67424\,
            I => \ALU.c_RNIO5N04AZ0Z_13\
        );

    \I__16138\ : LocalMux
    port map (
            O => \N__67421\,
            I => \ALU.c_RNIO5N04AZ0Z_13\
        );

    \I__16137\ : Odrv4
    port map (
            O => \N__67414\,
            I => \ALU.c_RNIO5N04AZ0Z_13\
        );

    \I__16136\ : LocalMux
    port map (
            O => \N__67411\,
            I => \ALU.c_RNIO5N04AZ0Z_13\
        );

    \I__16135\ : InMux
    port map (
            O => \N__67400\,
            I => \N__67396\
        );

    \I__16134\ : InMux
    port map (
            O => \N__67399\,
            I => \N__67393\
        );

    \I__16133\ : LocalMux
    port map (
            O => \N__67396\,
            I => \N__67385\
        );

    \I__16132\ : LocalMux
    port map (
            O => \N__67393\,
            I => \N__67382\
        );

    \I__16131\ : InMux
    port map (
            O => \N__67392\,
            I => \N__67379\
        );

    \I__16130\ : InMux
    port map (
            O => \N__67391\,
            I => \N__67376\
        );

    \I__16129\ : InMux
    port map (
            O => \N__67390\,
            I => \N__67373\
        );

    \I__16128\ : InMux
    port map (
            O => \N__67389\,
            I => \N__67370\
        );

    \I__16127\ : InMux
    port map (
            O => \N__67388\,
            I => \N__67367\
        );

    \I__16126\ : Odrv4
    port map (
            O => \N__67385\,
            I => \ALU.mult_558_c_RNIB75F9GZ0\
        );

    \I__16125\ : Odrv4
    port map (
            O => \N__67382\,
            I => \ALU.mult_558_c_RNIB75F9GZ0\
        );

    \I__16124\ : LocalMux
    port map (
            O => \N__67379\,
            I => \ALU.mult_558_c_RNIB75F9GZ0\
        );

    \I__16123\ : LocalMux
    port map (
            O => \N__67376\,
            I => \ALU.mult_558_c_RNIB75F9GZ0\
        );

    \I__16122\ : LocalMux
    port map (
            O => \N__67373\,
            I => \ALU.mult_558_c_RNIB75F9GZ0\
        );

    \I__16121\ : LocalMux
    port map (
            O => \N__67370\,
            I => \ALU.mult_558_c_RNIB75F9GZ0\
        );

    \I__16120\ : LocalMux
    port map (
            O => \N__67367\,
            I => \ALU.mult_558_c_RNIB75F9GZ0\
        );

    \I__16119\ : InMux
    port map (
            O => \N__67352\,
            I => \N__67349\
        );

    \I__16118\ : LocalMux
    port map (
            O => \N__67349\,
            I => \N__67345\
        );

    \I__16117\ : InMux
    port map (
            O => \N__67348\,
            I => \N__67342\
        );

    \I__16116\ : Span4Mux_h
    port map (
            O => \N__67345\,
            I => \N__67339\
        );

    \I__16115\ : LocalMux
    port map (
            O => \N__67342\,
            I => \N__67336\
        );

    \I__16114\ : Span4Mux_v
    port map (
            O => \N__67339\,
            I => \N__67333\
        );

    \I__16113\ : Span4Mux_v
    port map (
            O => \N__67336\,
            I => \N__67330\
        );

    \I__16112\ : Span4Mux_h
    port map (
            O => \N__67333\,
            I => \N__67327\
        );

    \I__16111\ : Span4Mux_v
    port map (
            O => \N__67330\,
            I => \N__67324\
        );

    \I__16110\ : Span4Mux_h
    port map (
            O => \N__67327\,
            I => \N__67321\
        );

    \I__16109\ : Span4Mux_h
    port map (
            O => \N__67324\,
            I => \N__67316\
        );

    \I__16108\ : Span4Mux_v
    port map (
            O => \N__67321\,
            I => \N__67316\
        );

    \I__16107\ : Odrv4
    port map (
            O => \N__67316\,
            I => \ALU.cZ0Z_13\
        );

    \I__16106\ : InMux
    port map (
            O => \N__67313\,
            I => \N__67309\
        );

    \I__16105\ : InMux
    port map (
            O => \N__67312\,
            I => \N__67306\
        );

    \I__16104\ : LocalMux
    port map (
            O => \N__67309\,
            I => \N__67303\
        );

    \I__16103\ : LocalMux
    port map (
            O => \N__67306\,
            I => \N__67300\
        );

    \I__16102\ : Span4Mux_v
    port map (
            O => \N__67303\,
            I => \N__67297\
        );

    \I__16101\ : Span4Mux_v
    port map (
            O => \N__67300\,
            I => \N__67294\
        );

    \I__16100\ : Span4Mux_h
    port map (
            O => \N__67297\,
            I => \N__67289\
        );

    \I__16099\ : Span4Mux_h
    port map (
            O => \N__67294\,
            I => \N__67289\
        );

    \I__16098\ : Odrv4
    port map (
            O => \N__67289\,
            I => \ALU.cZ0Z_14\
        );

    \I__16097\ : CascadeMux
    port map (
            O => \N__67286\,
            I => \N__67283\
        );

    \I__16096\ : InMux
    port map (
            O => \N__67283\,
            I => \N__67277\
        );

    \I__16095\ : InMux
    port map (
            O => \N__67282\,
            I => \N__67277\
        );

    \I__16094\ : LocalMux
    port map (
            O => \N__67277\,
            I => \N__67274\
        );

    \I__16093\ : Span4Mux_v
    port map (
            O => \N__67274\,
            I => \N__67263\
        );

    \I__16092\ : InMux
    port map (
            O => \N__67273\,
            I => \N__67256\
        );

    \I__16091\ : InMux
    port map (
            O => \N__67272\,
            I => \N__67256\
        );

    \I__16090\ : InMux
    port map (
            O => \N__67271\,
            I => \N__67256\
        );

    \I__16089\ : CascadeMux
    port map (
            O => \N__67270\,
            I => \N__67245\
        );

    \I__16088\ : InMux
    port map (
            O => \N__67269\,
            I => \N__67239\
        );

    \I__16087\ : CascadeMux
    port map (
            O => \N__67268\,
            I => \N__67236\
        );

    \I__16086\ : CascadeMux
    port map (
            O => \N__67267\,
            I => \N__67233\
        );

    \I__16085\ : CascadeMux
    port map (
            O => \N__67266\,
            I => \N__67227\
        );

    \I__16084\ : Span4Mux_h
    port map (
            O => \N__67263\,
            I => \N__67220\
        );

    \I__16083\ : LocalMux
    port map (
            O => \N__67256\,
            I => \N__67220\
        );

    \I__16082\ : CascadeMux
    port map (
            O => \N__67255\,
            I => \N__67209\
        );

    \I__16081\ : InMux
    port map (
            O => \N__67254\,
            I => \N__67197\
        );

    \I__16080\ : InMux
    port map (
            O => \N__67253\,
            I => \N__67197\
        );

    \I__16079\ : InMux
    port map (
            O => \N__67252\,
            I => \N__67197\
        );

    \I__16078\ : InMux
    port map (
            O => \N__67251\,
            I => \N__67184\
        );

    \I__16077\ : InMux
    port map (
            O => \N__67250\,
            I => \N__67184\
        );

    \I__16076\ : InMux
    port map (
            O => \N__67249\,
            I => \N__67184\
        );

    \I__16075\ : InMux
    port map (
            O => \N__67248\,
            I => \N__67184\
        );

    \I__16074\ : InMux
    port map (
            O => \N__67245\,
            I => \N__67184\
        );

    \I__16073\ : InMux
    port map (
            O => \N__67244\,
            I => \N__67184\
        );

    \I__16072\ : CascadeMux
    port map (
            O => \N__67243\,
            I => \N__67180\
        );

    \I__16071\ : CascadeMux
    port map (
            O => \N__67242\,
            I => \N__67176\
        );

    \I__16070\ : LocalMux
    port map (
            O => \N__67239\,
            I => \N__67173\
        );

    \I__16069\ : InMux
    port map (
            O => \N__67236\,
            I => \N__67170\
        );

    \I__16068\ : InMux
    port map (
            O => \N__67233\,
            I => \N__67165\
        );

    \I__16067\ : InMux
    port map (
            O => \N__67232\,
            I => \N__67165\
        );

    \I__16066\ : InMux
    port map (
            O => \N__67231\,
            I => \N__67161\
        );

    \I__16065\ : InMux
    port map (
            O => \N__67230\,
            I => \N__67158\
        );

    \I__16064\ : InMux
    port map (
            O => \N__67227\,
            I => \N__67151\
        );

    \I__16063\ : InMux
    port map (
            O => \N__67226\,
            I => \N__67151\
        );

    \I__16062\ : InMux
    port map (
            O => \N__67225\,
            I => \N__67151\
        );

    \I__16061\ : Span4Mux_v
    port map (
            O => \N__67220\,
            I => \N__67148\
        );

    \I__16060\ : InMux
    port map (
            O => \N__67219\,
            I => \N__67145\
        );

    \I__16059\ : InMux
    port map (
            O => \N__67218\,
            I => \N__67138\
        );

    \I__16058\ : InMux
    port map (
            O => \N__67217\,
            I => \N__67138\
        );

    \I__16057\ : InMux
    port map (
            O => \N__67216\,
            I => \N__67138\
        );

    \I__16056\ : InMux
    port map (
            O => \N__67215\,
            I => \N__67135\
        );

    \I__16055\ : InMux
    port map (
            O => \N__67214\,
            I => \N__67130\
        );

    \I__16054\ : InMux
    port map (
            O => \N__67213\,
            I => \N__67130\
        );

    \I__16053\ : InMux
    port map (
            O => \N__67212\,
            I => \N__67123\
        );

    \I__16052\ : InMux
    port map (
            O => \N__67209\,
            I => \N__67123\
        );

    \I__16051\ : InMux
    port map (
            O => \N__67208\,
            I => \N__67123\
        );

    \I__16050\ : InMux
    port map (
            O => \N__67207\,
            I => \N__67116\
        );

    \I__16049\ : InMux
    port map (
            O => \N__67206\,
            I => \N__67116\
        );

    \I__16048\ : InMux
    port map (
            O => \N__67205\,
            I => \N__67116\
        );

    \I__16047\ : CascadeMux
    port map (
            O => \N__67204\,
            I => \N__67112\
        );

    \I__16046\ : LocalMux
    port map (
            O => \N__67197\,
            I => \N__67107\
        );

    \I__16045\ : LocalMux
    port map (
            O => \N__67184\,
            I => \N__67107\
        );

    \I__16044\ : InMux
    port map (
            O => \N__67183\,
            I => \N__67100\
        );

    \I__16043\ : InMux
    port map (
            O => \N__67180\,
            I => \N__67100\
        );

    \I__16042\ : InMux
    port map (
            O => \N__67179\,
            I => \N__67100\
        );

    \I__16041\ : InMux
    port map (
            O => \N__67176\,
            I => \N__67097\
        );

    \I__16040\ : Span4Mux_h
    port map (
            O => \N__67173\,
            I => \N__67090\
        );

    \I__16039\ : LocalMux
    port map (
            O => \N__67170\,
            I => \N__67090\
        );

    \I__16038\ : LocalMux
    port map (
            O => \N__67165\,
            I => \N__67090\
        );

    \I__16037\ : InMux
    port map (
            O => \N__67164\,
            I => \N__67087\
        );

    \I__16036\ : LocalMux
    port map (
            O => \N__67161\,
            I => \N__67066\
        );

    \I__16035\ : LocalMux
    port map (
            O => \N__67158\,
            I => \N__67066\
        );

    \I__16034\ : LocalMux
    port map (
            O => \N__67151\,
            I => \N__67066\
        );

    \I__16033\ : Span4Mux_v
    port map (
            O => \N__67148\,
            I => \N__67066\
        );

    \I__16032\ : LocalMux
    port map (
            O => \N__67145\,
            I => \N__67066\
        );

    \I__16031\ : LocalMux
    port map (
            O => \N__67138\,
            I => \N__67066\
        );

    \I__16030\ : LocalMux
    port map (
            O => \N__67135\,
            I => \N__67066\
        );

    \I__16029\ : LocalMux
    port map (
            O => \N__67130\,
            I => \N__67066\
        );

    \I__16028\ : LocalMux
    port map (
            O => \N__67123\,
            I => \N__67066\
        );

    \I__16027\ : LocalMux
    port map (
            O => \N__67116\,
            I => \N__67066\
        );

    \I__16026\ : CascadeMux
    port map (
            O => \N__67115\,
            I => \N__67061\
        );

    \I__16025\ : InMux
    port map (
            O => \N__67112\,
            I => \N__67057\
        );

    \I__16024\ : Span4Mux_v
    port map (
            O => \N__67107\,
            I => \N__67054\
        );

    \I__16023\ : LocalMux
    port map (
            O => \N__67100\,
            I => \N__67048\
        );

    \I__16022\ : LocalMux
    port map (
            O => \N__67097\,
            I => \N__67039\
        );

    \I__16021\ : Span4Mux_v
    port map (
            O => \N__67090\,
            I => \N__67036\
        );

    \I__16020\ : LocalMux
    port map (
            O => \N__67087\,
            I => \N__67033\
        );

    \I__16019\ : Span4Mux_v
    port map (
            O => \N__67066\,
            I => \N__67030\
        );

    \I__16018\ : InMux
    port map (
            O => \N__67065\,
            I => \N__67027\
        );

    \I__16017\ : InMux
    port map (
            O => \N__67064\,
            I => \N__67020\
        );

    \I__16016\ : InMux
    port map (
            O => \N__67061\,
            I => \N__67020\
        );

    \I__16015\ : InMux
    port map (
            O => \N__67060\,
            I => \N__67020\
        );

    \I__16014\ : LocalMux
    port map (
            O => \N__67057\,
            I => \N__67017\
        );

    \I__16013\ : Span4Mux_h
    port map (
            O => \N__67054\,
            I => \N__67014\
        );

    \I__16012\ : InMux
    port map (
            O => \N__67053\,
            I => \N__67007\
        );

    \I__16011\ : InMux
    port map (
            O => \N__67052\,
            I => \N__67007\
        );

    \I__16010\ : InMux
    port map (
            O => \N__67051\,
            I => \N__67007\
        );

    \I__16009\ : Span4Mux_v
    port map (
            O => \N__67048\,
            I => \N__67004\
        );

    \I__16008\ : InMux
    port map (
            O => \N__67047\,
            I => \N__66997\
        );

    \I__16007\ : InMux
    port map (
            O => \N__67046\,
            I => \N__66997\
        );

    \I__16006\ : InMux
    port map (
            O => \N__67045\,
            I => \N__66997\
        );

    \I__16005\ : InMux
    port map (
            O => \N__67044\,
            I => \N__66994\
        );

    \I__16004\ : InMux
    port map (
            O => \N__67043\,
            I => \N__66991\
        );

    \I__16003\ : InMux
    port map (
            O => \N__67042\,
            I => \N__66988\
        );

    \I__16002\ : Span4Mux_v
    port map (
            O => \N__67039\,
            I => \N__66985\
        );

    \I__16001\ : Span4Mux_h
    port map (
            O => \N__67036\,
            I => \N__66982\
        );

    \I__16000\ : Span4Mux_v
    port map (
            O => \N__67033\,
            I => \N__66977\
        );

    \I__15999\ : Span4Mux_h
    port map (
            O => \N__67030\,
            I => \N__66977\
        );

    \I__15998\ : LocalMux
    port map (
            O => \N__67027\,
            I => \N__66973\
        );

    \I__15997\ : LocalMux
    port map (
            O => \N__67020\,
            I => \N__66970\
        );

    \I__15996\ : Span4Mux_h
    port map (
            O => \N__67017\,
            I => \N__66963\
        );

    \I__15995\ : Span4Mux_h
    port map (
            O => \N__67014\,
            I => \N__66963\
        );

    \I__15994\ : LocalMux
    port map (
            O => \N__67007\,
            I => \N__66963\
        );

    \I__15993\ : Span4Mux_h
    port map (
            O => \N__67004\,
            I => \N__66958\
        );

    \I__15992\ : LocalMux
    port map (
            O => \N__66997\,
            I => \N__66958\
        );

    \I__15991\ : LocalMux
    port map (
            O => \N__66994\,
            I => \N__66951\
        );

    \I__15990\ : LocalMux
    port map (
            O => \N__66991\,
            I => \N__66951\
        );

    \I__15989\ : LocalMux
    port map (
            O => \N__66988\,
            I => \N__66951\
        );

    \I__15988\ : Span4Mux_h
    port map (
            O => \N__66985\,
            I => \N__66948\
        );

    \I__15987\ : Span4Mux_h
    port map (
            O => \N__66982\,
            I => \N__66945\
        );

    \I__15986\ : Span4Mux_v
    port map (
            O => \N__66977\,
            I => \N__66942\
        );

    \I__15985\ : InMux
    port map (
            O => \N__66976\,
            I => \N__66939\
        );

    \I__15984\ : Span4Mux_v
    port map (
            O => \N__66973\,
            I => \N__66930\
        );

    \I__15983\ : Span4Mux_v
    port map (
            O => \N__66970\,
            I => \N__66930\
        );

    \I__15982\ : Span4Mux_v
    port map (
            O => \N__66963\,
            I => \N__66930\
        );

    \I__15981\ : Span4Mux_h
    port map (
            O => \N__66958\,
            I => \N__66930\
        );

    \I__15980\ : Sp12to4
    port map (
            O => \N__66951\,
            I => \N__66927\
        );

    \I__15979\ : Sp12to4
    port map (
            O => \N__66948\,
            I => \N__66920\
        );

    \I__15978\ : Sp12to4
    port map (
            O => \N__66945\,
            I => \N__66920\
        );

    \I__15977\ : Sp12to4
    port map (
            O => \N__66942\,
            I => \N__66920\
        );

    \I__15976\ : LocalMux
    port map (
            O => \N__66939\,
            I => \N__66915\
        );

    \I__15975\ : Span4Mux_h
    port map (
            O => \N__66930\,
            I => \N__66915\
        );

    \I__15974\ : Span12Mux_v
    port map (
            O => \N__66927\,
            I => \N__66910\
        );

    \I__15973\ : Span12Mux_h
    port map (
            O => \N__66920\,
            I => \N__66910\
        );

    \I__15972\ : Span4Mux_v
    port map (
            O => \N__66915\,
            I => \N__66907\
        );

    \I__15971\ : Odrv12
    port map (
            O => \N__66910\,
            I => \aluOperation_0\
        );

    \I__15970\ : Odrv4
    port map (
            O => \N__66907\,
            I => \aluOperation_0\
        );

    \I__15969\ : CascadeMux
    port map (
            O => \N__66902\,
            I => \N__66898\
        );

    \I__15968\ : InMux
    port map (
            O => \N__66901\,
            I => \N__66891\
        );

    \I__15967\ : InMux
    port map (
            O => \N__66898\,
            I => \N__66891\
        );

    \I__15966\ : CascadeMux
    port map (
            O => \N__66897\,
            I => \N__66888\
        );

    \I__15965\ : InMux
    port map (
            O => \N__66896\,
            I => \N__66885\
        );

    \I__15964\ : LocalMux
    port map (
            O => \N__66891\,
            I => \N__66882\
        );

    \I__15963\ : InMux
    port map (
            O => \N__66888\,
            I => \N__66879\
        );

    \I__15962\ : LocalMux
    port map (
            O => \N__66885\,
            I => \N__66876\
        );

    \I__15961\ : Span4Mux_v
    port map (
            O => \N__66882\,
            I => \N__66873\
        );

    \I__15960\ : LocalMux
    port map (
            O => \N__66879\,
            I => \N__66870\
        );

    \I__15959\ : Span4Mux_v
    port map (
            O => \N__66876\,
            I => \N__66865\
        );

    \I__15958\ : Span4Mux_h
    port map (
            O => \N__66873\,
            I => \N__66865\
        );

    \I__15957\ : Odrv4
    port map (
            O => \N__66870\,
            I => \ALU.a_15_d_sZ0Z_10\
        );

    \I__15956\ : Odrv4
    port map (
            O => \N__66865\,
            I => \ALU.a_15_d_sZ0Z_10\
        );

    \I__15955\ : InMux
    port map (
            O => \N__66860\,
            I => \N__66857\
        );

    \I__15954\ : LocalMux
    port map (
            O => \N__66857\,
            I => \N__66853\
        );

    \I__15953\ : InMux
    port map (
            O => \N__66856\,
            I => \N__66850\
        );

    \I__15952\ : Odrv4
    port map (
            O => \N__66853\,
            I => \ALU.addsub_9\
        );

    \I__15951\ : LocalMux
    port map (
            O => \N__66850\,
            I => \ALU.addsub_9\
        );

    \I__15950\ : InMux
    port map (
            O => \N__66845\,
            I => \N__66840\
        );

    \I__15949\ : InMux
    port map (
            O => \N__66844\,
            I => \N__66837\
        );

    \I__15948\ : InMux
    port map (
            O => \N__66843\,
            I => \N__66834\
        );

    \I__15947\ : LocalMux
    port map (
            O => \N__66840\,
            I => \N__66828\
        );

    \I__15946\ : LocalMux
    port map (
            O => \N__66837\,
            I => \N__66822\
        );

    \I__15945\ : LocalMux
    port map (
            O => \N__66834\,
            I => \N__66822\
        );

    \I__15944\ : InMux
    port map (
            O => \N__66833\,
            I => \N__66819\
        );

    \I__15943\ : InMux
    port map (
            O => \N__66832\,
            I => \N__66816\
        );

    \I__15942\ : InMux
    port map (
            O => \N__66831\,
            I => \N__66813\
        );

    \I__15941\ : Span4Mux_v
    port map (
            O => \N__66828\,
            I => \N__66810\
        );

    \I__15940\ : InMux
    port map (
            O => \N__66827\,
            I => \N__66807\
        );

    \I__15939\ : Sp12to4
    port map (
            O => \N__66822\,
            I => \N__66801\
        );

    \I__15938\ : LocalMux
    port map (
            O => \N__66819\,
            I => \N__66801\
        );

    \I__15937\ : LocalMux
    port map (
            O => \N__66816\,
            I => \N__66796\
        );

    \I__15936\ : LocalMux
    port map (
            O => \N__66813\,
            I => \N__66796\
        );

    \I__15935\ : Span4Mux_v
    port map (
            O => \N__66810\,
            I => \N__66791\
        );

    \I__15934\ : LocalMux
    port map (
            O => \N__66807\,
            I => \N__66791\
        );

    \I__15933\ : InMux
    port map (
            O => \N__66806\,
            I => \N__66788\
        );

    \I__15932\ : Span12Mux_v
    port map (
            O => \N__66801\,
            I => \N__66785\
        );

    \I__15931\ : Span4Mux_v
    port map (
            O => \N__66796\,
            I => \N__66778\
        );

    \I__15930\ : Span4Mux_h
    port map (
            O => \N__66791\,
            I => \N__66778\
        );

    \I__15929\ : LocalMux
    port map (
            O => \N__66788\,
            I => \N__66778\
        );

    \I__15928\ : Odrv12
    port map (
            O => \N__66785\,
            I => \ALU.a_15_d_ns_sx_9\
        );

    \I__15927\ : Odrv4
    port map (
            O => \N__66778\,
            I => \ALU.a_15_d_ns_sx_9\
        );

    \I__15926\ : CascadeMux
    port map (
            O => \N__66773\,
            I => \N__66769\
        );

    \I__15925\ : InMux
    port map (
            O => \N__66772\,
            I => \N__66758\
        );

    \I__15924\ : InMux
    port map (
            O => \N__66769\,
            I => \N__66750\
        );

    \I__15923\ : InMux
    port map (
            O => \N__66768\,
            I => \N__66747\
        );

    \I__15922\ : CascadeMux
    port map (
            O => \N__66767\,
            I => \N__66743\
        );

    \I__15921\ : InMux
    port map (
            O => \N__66766\,
            I => \N__66737\
        );

    \I__15920\ : InMux
    port map (
            O => \N__66765\,
            I => \N__66737\
        );

    \I__15919\ : InMux
    port map (
            O => \N__66764\,
            I => \N__66730\
        );

    \I__15918\ : InMux
    port map (
            O => \N__66763\,
            I => \N__66727\
        );

    \I__15917\ : InMux
    port map (
            O => \N__66762\,
            I => \N__66722\
        );

    \I__15916\ : InMux
    port map (
            O => \N__66761\,
            I => \N__66722\
        );

    \I__15915\ : LocalMux
    port map (
            O => \N__66758\,
            I => \N__66710\
        );

    \I__15914\ : InMux
    port map (
            O => \N__66757\,
            I => \N__66705\
        );

    \I__15913\ : InMux
    port map (
            O => \N__66756\,
            I => \N__66705\
        );

    \I__15912\ : CascadeMux
    port map (
            O => \N__66755\,
            I => \N__66693\
        );

    \I__15911\ : InMux
    port map (
            O => \N__66754\,
            I => \N__66690\
        );

    \I__15910\ : InMux
    port map (
            O => \N__66753\,
            I => \N__66687\
        );

    \I__15909\ : LocalMux
    port map (
            O => \N__66750\,
            I => \N__66677\
        );

    \I__15908\ : LocalMux
    port map (
            O => \N__66747\,
            I => \N__66677\
        );

    \I__15907\ : InMux
    port map (
            O => \N__66746\,
            I => \N__66672\
        );

    \I__15906\ : InMux
    port map (
            O => \N__66743\,
            I => \N__66672\
        );

    \I__15905\ : InMux
    port map (
            O => \N__66742\,
            I => \N__66669\
        );

    \I__15904\ : LocalMux
    port map (
            O => \N__66737\,
            I => \N__66666\
        );

    \I__15903\ : InMux
    port map (
            O => \N__66736\,
            I => \N__66663\
        );

    \I__15902\ : InMux
    port map (
            O => \N__66735\,
            I => \N__66659\
        );

    \I__15901\ : InMux
    port map (
            O => \N__66734\,
            I => \N__66654\
        );

    \I__15900\ : InMux
    port map (
            O => \N__66733\,
            I => \N__66654\
        );

    \I__15899\ : LocalMux
    port map (
            O => \N__66730\,
            I => \N__66647\
        );

    \I__15898\ : LocalMux
    port map (
            O => \N__66727\,
            I => \N__66647\
        );

    \I__15897\ : LocalMux
    port map (
            O => \N__66722\,
            I => \N__66644\
        );

    \I__15896\ : InMux
    port map (
            O => \N__66721\,
            I => \N__66641\
        );

    \I__15895\ : InMux
    port map (
            O => \N__66720\,
            I => \N__66634\
        );

    \I__15894\ : InMux
    port map (
            O => \N__66719\,
            I => \N__66634\
        );

    \I__15893\ : InMux
    port map (
            O => \N__66718\,
            I => \N__66634\
        );

    \I__15892\ : CascadeMux
    port map (
            O => \N__66717\,
            I => \N__66631\
        );

    \I__15891\ : InMux
    port map (
            O => \N__66716\,
            I => \N__66626\
        );

    \I__15890\ : InMux
    port map (
            O => \N__66715\,
            I => \N__66623\
        );

    \I__15889\ : InMux
    port map (
            O => \N__66714\,
            I => \N__66618\
        );

    \I__15888\ : InMux
    port map (
            O => \N__66713\,
            I => \N__66618\
        );

    \I__15887\ : Span4Mux_h
    port map (
            O => \N__66710\,
            I => \N__66615\
        );

    \I__15886\ : LocalMux
    port map (
            O => \N__66705\,
            I => \N__66612\
        );

    \I__15885\ : InMux
    port map (
            O => \N__66704\,
            I => \N__66609\
        );

    \I__15884\ : InMux
    port map (
            O => \N__66703\,
            I => \N__66604\
        );

    \I__15883\ : InMux
    port map (
            O => \N__66702\,
            I => \N__66604\
        );

    \I__15882\ : InMux
    port map (
            O => \N__66701\,
            I => \N__66591\
        );

    \I__15881\ : InMux
    port map (
            O => \N__66700\,
            I => \N__66591\
        );

    \I__15880\ : InMux
    port map (
            O => \N__66699\,
            I => \N__66586\
        );

    \I__15879\ : InMux
    port map (
            O => \N__66698\,
            I => \N__66586\
        );

    \I__15878\ : InMux
    port map (
            O => \N__66697\,
            I => \N__66583\
        );

    \I__15877\ : CascadeMux
    port map (
            O => \N__66696\,
            I => \N__66574\
        );

    \I__15876\ : InMux
    port map (
            O => \N__66693\,
            I => \N__66571\
        );

    \I__15875\ : LocalMux
    port map (
            O => \N__66690\,
            I => \N__66564\
        );

    \I__15874\ : LocalMux
    port map (
            O => \N__66687\,
            I => \N__66564\
        );

    \I__15873\ : InMux
    port map (
            O => \N__66686\,
            I => \N__66559\
        );

    \I__15872\ : InMux
    port map (
            O => \N__66685\,
            I => \N__66559\
        );

    \I__15871\ : InMux
    port map (
            O => \N__66684\,
            I => \N__66552\
        );

    \I__15870\ : InMux
    port map (
            O => \N__66683\,
            I => \N__66552\
        );

    \I__15869\ : InMux
    port map (
            O => \N__66682\,
            I => \N__66552\
        );

    \I__15868\ : Span4Mux_v
    port map (
            O => \N__66677\,
            I => \N__66547\
        );

    \I__15867\ : LocalMux
    port map (
            O => \N__66672\,
            I => \N__66547\
        );

    \I__15866\ : LocalMux
    port map (
            O => \N__66669\,
            I => \N__66540\
        );

    \I__15865\ : Span4Mux_v
    port map (
            O => \N__66666\,
            I => \N__66540\
        );

    \I__15864\ : LocalMux
    port map (
            O => \N__66663\,
            I => \N__66540\
        );

    \I__15863\ : InMux
    port map (
            O => \N__66662\,
            I => \N__66537\
        );

    \I__15862\ : LocalMux
    port map (
            O => \N__66659\,
            I => \N__66532\
        );

    \I__15861\ : LocalMux
    port map (
            O => \N__66654\,
            I => \N__66532\
        );

    \I__15860\ : InMux
    port map (
            O => \N__66653\,
            I => \N__66529\
        );

    \I__15859\ : InMux
    port map (
            O => \N__66652\,
            I => \N__66526\
        );

    \I__15858\ : Span4Mux_h
    port map (
            O => \N__66647\,
            I => \N__66523\
        );

    \I__15857\ : Span4Mux_h
    port map (
            O => \N__66644\,
            I => \N__66516\
        );

    \I__15856\ : LocalMux
    port map (
            O => \N__66641\,
            I => \N__66516\
        );

    \I__15855\ : LocalMux
    port map (
            O => \N__66634\,
            I => \N__66516\
        );

    \I__15854\ : InMux
    port map (
            O => \N__66631\,
            I => \N__66513\
        );

    \I__15853\ : InMux
    port map (
            O => \N__66630\,
            I => \N__66508\
        );

    \I__15852\ : InMux
    port map (
            O => \N__66629\,
            I => \N__66508\
        );

    \I__15851\ : LocalMux
    port map (
            O => \N__66626\,
            I => \N__66501\
        );

    \I__15850\ : LocalMux
    port map (
            O => \N__66623\,
            I => \N__66501\
        );

    \I__15849\ : LocalMux
    port map (
            O => \N__66618\,
            I => \N__66501\
        );

    \I__15848\ : Span4Mux_v
    port map (
            O => \N__66615\,
            I => \N__66492\
        );

    \I__15847\ : Span4Mux_v
    port map (
            O => \N__66612\,
            I => \N__66492\
        );

    \I__15846\ : LocalMux
    port map (
            O => \N__66609\,
            I => \N__66492\
        );

    \I__15845\ : LocalMux
    port map (
            O => \N__66604\,
            I => \N__66492\
        );

    \I__15844\ : InMux
    port map (
            O => \N__66603\,
            I => \N__66487\
        );

    \I__15843\ : InMux
    port map (
            O => \N__66602\,
            I => \N__66487\
        );

    \I__15842\ : InMux
    port map (
            O => \N__66601\,
            I => \N__66482\
        );

    \I__15841\ : InMux
    port map (
            O => \N__66600\,
            I => \N__66482\
        );

    \I__15840\ : InMux
    port map (
            O => \N__66599\,
            I => \N__66473\
        );

    \I__15839\ : InMux
    port map (
            O => \N__66598\,
            I => \N__66473\
        );

    \I__15838\ : InMux
    port map (
            O => \N__66597\,
            I => \N__66473\
        );

    \I__15837\ : InMux
    port map (
            O => \N__66596\,
            I => \N__66473\
        );

    \I__15836\ : LocalMux
    port map (
            O => \N__66591\,
            I => \N__66468\
        );

    \I__15835\ : LocalMux
    port map (
            O => \N__66586\,
            I => \N__66468\
        );

    \I__15834\ : LocalMux
    port map (
            O => \N__66583\,
            I => \N__66465\
        );

    \I__15833\ : InMux
    port map (
            O => \N__66582\,
            I => \N__66462\
        );

    \I__15832\ : InMux
    port map (
            O => \N__66581\,
            I => \N__66451\
        );

    \I__15831\ : InMux
    port map (
            O => \N__66580\,
            I => \N__66451\
        );

    \I__15830\ : InMux
    port map (
            O => \N__66579\,
            I => \N__66451\
        );

    \I__15829\ : InMux
    port map (
            O => \N__66578\,
            I => \N__66451\
        );

    \I__15828\ : InMux
    port map (
            O => \N__66577\,
            I => \N__66451\
        );

    \I__15827\ : InMux
    port map (
            O => \N__66574\,
            I => \N__66448\
        );

    \I__15826\ : LocalMux
    port map (
            O => \N__66571\,
            I => \N__66445\
        );

    \I__15825\ : InMux
    port map (
            O => \N__66570\,
            I => \N__66442\
        );

    \I__15824\ : InMux
    port map (
            O => \N__66569\,
            I => \N__66438\
        );

    \I__15823\ : Span4Mux_v
    port map (
            O => \N__66564\,
            I => \N__66435\
        );

    \I__15822\ : LocalMux
    port map (
            O => \N__66559\,
            I => \N__66426\
        );

    \I__15821\ : LocalMux
    port map (
            O => \N__66552\,
            I => \N__66426\
        );

    \I__15820\ : Span4Mux_v
    port map (
            O => \N__66547\,
            I => \N__66426\
        );

    \I__15819\ : Span4Mux_h
    port map (
            O => \N__66540\,
            I => \N__66426\
        );

    \I__15818\ : LocalMux
    port map (
            O => \N__66537\,
            I => \N__66421\
        );

    \I__15817\ : Span4Mux_v
    port map (
            O => \N__66532\,
            I => \N__66421\
        );

    \I__15816\ : LocalMux
    port map (
            O => \N__66529\,
            I => \N__66418\
        );

    \I__15815\ : LocalMux
    port map (
            O => \N__66526\,
            I => \N__66415\
        );

    \I__15814\ : Span4Mux_v
    port map (
            O => \N__66523\,
            I => \N__66410\
        );

    \I__15813\ : Span4Mux_h
    port map (
            O => \N__66516\,
            I => \N__66410\
        );

    \I__15812\ : LocalMux
    port map (
            O => \N__66513\,
            I => \N__66401\
        );

    \I__15811\ : LocalMux
    port map (
            O => \N__66508\,
            I => \N__66401\
        );

    \I__15810\ : Span4Mux_v
    port map (
            O => \N__66501\,
            I => \N__66401\
        );

    \I__15809\ : Span4Mux_h
    port map (
            O => \N__66492\,
            I => \N__66401\
        );

    \I__15808\ : LocalMux
    port map (
            O => \N__66487\,
            I => \N__66394\
        );

    \I__15807\ : LocalMux
    port map (
            O => \N__66482\,
            I => \N__66394\
        );

    \I__15806\ : LocalMux
    port map (
            O => \N__66473\,
            I => \N__66394\
        );

    \I__15805\ : Span4Mux_h
    port map (
            O => \N__66468\,
            I => \N__66385\
        );

    \I__15804\ : Span4Mux_v
    port map (
            O => \N__66465\,
            I => \N__66385\
        );

    \I__15803\ : LocalMux
    port map (
            O => \N__66462\,
            I => \N__66385\
        );

    \I__15802\ : LocalMux
    port map (
            O => \N__66451\,
            I => \N__66385\
        );

    \I__15801\ : LocalMux
    port map (
            O => \N__66448\,
            I => \N__66378\
        );

    \I__15800\ : Span4Mux_h
    port map (
            O => \N__66445\,
            I => \N__66378\
        );

    \I__15799\ : LocalMux
    port map (
            O => \N__66442\,
            I => \N__66378\
        );

    \I__15798\ : InMux
    port map (
            O => \N__66441\,
            I => \N__66372\
        );

    \I__15797\ : LocalMux
    port map (
            O => \N__66438\,
            I => \N__66369\
        );

    \I__15796\ : Span4Mux_v
    port map (
            O => \N__66435\,
            I => \N__66362\
        );

    \I__15795\ : Span4Mux_h
    port map (
            O => \N__66426\,
            I => \N__66362\
        );

    \I__15794\ : Span4Mux_v
    port map (
            O => \N__66421\,
            I => \N__66362\
        );

    \I__15793\ : Span4Mux_v
    port map (
            O => \N__66418\,
            I => \N__66355\
        );

    \I__15792\ : Span4Mux_v
    port map (
            O => \N__66415\,
            I => \N__66355\
        );

    \I__15791\ : Span4Mux_h
    port map (
            O => \N__66410\,
            I => \N__66355\
        );

    \I__15790\ : Span4Mux_h
    port map (
            O => \N__66401\,
            I => \N__66350\
        );

    \I__15789\ : Span4Mux_v
    port map (
            O => \N__66394\,
            I => \N__66350\
        );

    \I__15788\ : Span4Mux_h
    port map (
            O => \N__66385\,
            I => \N__66345\
        );

    \I__15787\ : Span4Mux_v
    port map (
            O => \N__66378\,
            I => \N__66345\
        );

    \I__15786\ : InMux
    port map (
            O => \N__66377\,
            I => \N__66340\
        );

    \I__15785\ : InMux
    port map (
            O => \N__66376\,
            I => \N__66340\
        );

    \I__15784\ : InMux
    port map (
            O => \N__66375\,
            I => \N__66337\
        );

    \I__15783\ : LocalMux
    port map (
            O => \N__66372\,
            I => \ALU.status_19\
        );

    \I__15782\ : Odrv4
    port map (
            O => \N__66369\,
            I => \ALU.status_19\
        );

    \I__15781\ : Odrv4
    port map (
            O => \N__66362\,
            I => \ALU.status_19\
        );

    \I__15780\ : Odrv4
    port map (
            O => \N__66355\,
            I => \ALU.status_19\
        );

    \I__15779\ : Odrv4
    port map (
            O => \N__66350\,
            I => \ALU.status_19\
        );

    \I__15778\ : Odrv4
    port map (
            O => \N__66345\,
            I => \ALU.status_19\
        );

    \I__15777\ : LocalMux
    port map (
            O => \N__66340\,
            I => \ALU.status_19\
        );

    \I__15776\ : LocalMux
    port map (
            O => \N__66337\,
            I => \ALU.status_19\
        );

    \I__15775\ : InMux
    port map (
            O => \N__66320\,
            I => \N__66317\
        );

    \I__15774\ : LocalMux
    port map (
            O => \N__66317\,
            I => \N__66309\
        );

    \I__15773\ : InMux
    port map (
            O => \N__66316\,
            I => \N__66304\
        );

    \I__15772\ : InMux
    port map (
            O => \N__66315\,
            I => \N__66304\
        );

    \I__15771\ : InMux
    port map (
            O => \N__66314\,
            I => \N__66300\
        );

    \I__15770\ : InMux
    port map (
            O => \N__66313\,
            I => \N__66293\
        );

    \I__15769\ : InMux
    port map (
            O => \N__66312\,
            I => \N__66289\
        );

    \I__15768\ : Span4Mux_v
    port map (
            O => \N__66309\,
            I => \N__66284\
        );

    \I__15767\ : LocalMux
    port map (
            O => \N__66304\,
            I => \N__66281\
        );

    \I__15766\ : InMux
    port map (
            O => \N__66303\,
            I => \N__66278\
        );

    \I__15765\ : LocalMux
    port map (
            O => \N__66300\,
            I => \N__66275\
        );

    \I__15764\ : InMux
    port map (
            O => \N__66299\,
            I => \N__66272\
        );

    \I__15763\ : InMux
    port map (
            O => \N__66298\,
            I => \N__66266\
        );

    \I__15762\ : InMux
    port map (
            O => \N__66297\,
            I => \N__66263\
        );

    \I__15761\ : InMux
    port map (
            O => \N__66296\,
            I => \N__66260\
        );

    \I__15760\ : LocalMux
    port map (
            O => \N__66293\,
            I => \N__66257\
        );

    \I__15759\ : InMux
    port map (
            O => \N__66292\,
            I => \N__66254\
        );

    \I__15758\ : LocalMux
    port map (
            O => \N__66289\,
            I => \N__66245\
        );

    \I__15757\ : InMux
    port map (
            O => \N__66288\,
            I => \N__66242\
        );

    \I__15756\ : InMux
    port map (
            O => \N__66287\,
            I => \N__66237\
        );

    \I__15755\ : Span4Mux_v
    port map (
            O => \N__66284\,
            I => \N__66230\
        );

    \I__15754\ : Span4Mux_v
    port map (
            O => \N__66281\,
            I => \N__66230\
        );

    \I__15753\ : LocalMux
    port map (
            O => \N__66278\,
            I => \N__66230\
        );

    \I__15752\ : Span4Mux_v
    port map (
            O => \N__66275\,
            I => \N__66225\
        );

    \I__15751\ : LocalMux
    port map (
            O => \N__66272\,
            I => \N__66222\
        );

    \I__15750\ : InMux
    port map (
            O => \N__66271\,
            I => \N__66215\
        );

    \I__15749\ : InMux
    port map (
            O => \N__66270\,
            I => \N__66215\
        );

    \I__15748\ : InMux
    port map (
            O => \N__66269\,
            I => \N__66215\
        );

    \I__15747\ : LocalMux
    port map (
            O => \N__66266\,
            I => \N__66208\
        );

    \I__15746\ : LocalMux
    port map (
            O => \N__66263\,
            I => \N__66208\
        );

    \I__15745\ : LocalMux
    port map (
            O => \N__66260\,
            I => \N__66208\
        );

    \I__15744\ : Span4Mux_v
    port map (
            O => \N__66257\,
            I => \N__66203\
        );

    \I__15743\ : LocalMux
    port map (
            O => \N__66254\,
            I => \N__66203\
        );

    \I__15742\ : InMux
    port map (
            O => \N__66253\,
            I => \N__66198\
        );

    \I__15741\ : InMux
    port map (
            O => \N__66252\,
            I => \N__66198\
        );

    \I__15740\ : InMux
    port map (
            O => \N__66251\,
            I => \N__66195\
        );

    \I__15739\ : InMux
    port map (
            O => \N__66250\,
            I => \N__66188\
        );

    \I__15738\ : InMux
    port map (
            O => \N__66249\,
            I => \N__66188\
        );

    \I__15737\ : InMux
    port map (
            O => \N__66248\,
            I => \N__66188\
        );

    \I__15736\ : Span4Mux_h
    port map (
            O => \N__66245\,
            I => \N__66183\
        );

    \I__15735\ : LocalMux
    port map (
            O => \N__66242\,
            I => \N__66183\
        );

    \I__15734\ : InMux
    port map (
            O => \N__66241\,
            I => \N__66180\
        );

    \I__15733\ : InMux
    port map (
            O => \N__66240\,
            I => \N__66177\
        );

    \I__15732\ : LocalMux
    port map (
            O => \N__66237\,
            I => \N__66169\
        );

    \I__15731\ : Span4Mux_h
    port map (
            O => \N__66230\,
            I => \N__66169\
        );

    \I__15730\ : InMux
    port map (
            O => \N__66229\,
            I => \N__66164\
        );

    \I__15729\ : InMux
    port map (
            O => \N__66228\,
            I => \N__66164\
        );

    \I__15728\ : Span4Mux_h
    port map (
            O => \N__66225\,
            I => \N__66161\
        );

    \I__15727\ : Span4Mux_v
    port map (
            O => \N__66222\,
            I => \N__66154\
        );

    \I__15726\ : LocalMux
    port map (
            O => \N__66215\,
            I => \N__66154\
        );

    \I__15725\ : Span4Mux_v
    port map (
            O => \N__66208\,
            I => \N__66154\
        );

    \I__15724\ : Span4Mux_v
    port map (
            O => \N__66203\,
            I => \N__66151\
        );

    \I__15723\ : LocalMux
    port map (
            O => \N__66198\,
            I => \N__66140\
        );

    \I__15722\ : LocalMux
    port map (
            O => \N__66195\,
            I => \N__66140\
        );

    \I__15721\ : LocalMux
    port map (
            O => \N__66188\,
            I => \N__66140\
        );

    \I__15720\ : Span4Mux_v
    port map (
            O => \N__66183\,
            I => \N__66140\
        );

    \I__15719\ : LocalMux
    port map (
            O => \N__66180\,
            I => \N__66140\
        );

    \I__15718\ : LocalMux
    port map (
            O => \N__66177\,
            I => \N__66137\
        );

    \I__15717\ : InMux
    port map (
            O => \N__66176\,
            I => \N__66134\
        );

    \I__15716\ : InMux
    port map (
            O => \N__66175\,
            I => \N__66131\
        );

    \I__15715\ : InMux
    port map (
            O => \N__66174\,
            I => \N__66128\
        );

    \I__15714\ : Span4Mux_h
    port map (
            O => \N__66169\,
            I => \N__66124\
        );

    \I__15713\ : LocalMux
    port map (
            O => \N__66164\,
            I => \N__66117\
        );

    \I__15712\ : Span4Mux_h
    port map (
            O => \N__66161\,
            I => \N__66117\
        );

    \I__15711\ : Span4Mux_h
    port map (
            O => \N__66154\,
            I => \N__66117\
        );

    \I__15710\ : Span4Mux_h
    port map (
            O => \N__66151\,
            I => \N__66112\
        );

    \I__15709\ : Span4Mux_v
    port map (
            O => \N__66140\,
            I => \N__66112\
        );

    \I__15708\ : Span12Mux_h
    port map (
            O => \N__66137\,
            I => \N__66103\
        );

    \I__15707\ : LocalMux
    port map (
            O => \N__66134\,
            I => \N__66103\
        );

    \I__15706\ : LocalMux
    port map (
            O => \N__66131\,
            I => \N__66103\
        );

    \I__15705\ : LocalMux
    port map (
            O => \N__66128\,
            I => \N__66103\
        );

    \I__15704\ : InMux
    port map (
            O => \N__66127\,
            I => \N__66100\
        );

    \I__15703\ : Odrv4
    port map (
            O => \N__66124\,
            I => \aluOut_2\
        );

    \I__15702\ : Odrv4
    port map (
            O => \N__66117\,
            I => \aluOut_2\
        );

    \I__15701\ : Odrv4
    port map (
            O => \N__66112\,
            I => \aluOut_2\
        );

    \I__15700\ : Odrv12
    port map (
            O => \N__66103\,
            I => \aluOut_2\
        );

    \I__15699\ : LocalMux
    port map (
            O => \N__66100\,
            I => \aluOut_2\
        );

    \I__15698\ : CascadeMux
    port map (
            O => \N__66089\,
            I => \N__66086\
        );

    \I__15697\ : InMux
    port map (
            O => \N__66086\,
            I => \N__66068\
        );

    \I__15696\ : InMux
    port map (
            O => \N__66085\,
            I => \N__66068\
        );

    \I__15695\ : InMux
    port map (
            O => \N__66084\,
            I => \N__66055\
        );

    \I__15694\ : CascadeMux
    port map (
            O => \N__66083\,
            I => \N__66052\
        );

    \I__15693\ : InMux
    port map (
            O => \N__66082\,
            I => \N__66040\
        );

    \I__15692\ : InMux
    port map (
            O => \N__66081\,
            I => \N__66040\
        );

    \I__15691\ : InMux
    port map (
            O => \N__66080\,
            I => \N__66037\
        );

    \I__15690\ : InMux
    port map (
            O => \N__66079\,
            I => \N__66030\
        );

    \I__15689\ : InMux
    port map (
            O => \N__66078\,
            I => \N__66030\
        );

    \I__15688\ : InMux
    port map (
            O => \N__66077\,
            I => \N__66030\
        );

    \I__15687\ : InMux
    port map (
            O => \N__66076\,
            I => \N__66023\
        );

    \I__15686\ : InMux
    port map (
            O => \N__66075\,
            I => \N__66020\
        );

    \I__15685\ : InMux
    port map (
            O => \N__66074\,
            I => \N__66015\
        );

    \I__15684\ : InMux
    port map (
            O => \N__66073\,
            I => \N__66015\
        );

    \I__15683\ : LocalMux
    port map (
            O => \N__66068\,
            I => \N__66007\
        );

    \I__15682\ : InMux
    port map (
            O => \N__66067\,
            I => \N__66000\
        );

    \I__15681\ : InMux
    port map (
            O => \N__66066\,
            I => \N__66000\
        );

    \I__15680\ : InMux
    port map (
            O => \N__66065\,
            I => \N__66000\
        );

    \I__15679\ : InMux
    port map (
            O => \N__66064\,
            I => \N__65991\
        );

    \I__15678\ : InMux
    port map (
            O => \N__66063\,
            I => \N__65991\
        );

    \I__15677\ : InMux
    port map (
            O => \N__66062\,
            I => \N__65991\
        );

    \I__15676\ : InMux
    port map (
            O => \N__66061\,
            I => \N__65991\
        );

    \I__15675\ : InMux
    port map (
            O => \N__66060\,
            I => \N__65986\
        );

    \I__15674\ : InMux
    port map (
            O => \N__66059\,
            I => \N__65981\
        );

    \I__15673\ : InMux
    port map (
            O => \N__66058\,
            I => \N__65981\
        );

    \I__15672\ : LocalMux
    port map (
            O => \N__66055\,
            I => \N__65978\
        );

    \I__15671\ : InMux
    port map (
            O => \N__66052\,
            I => \N__65969\
        );

    \I__15670\ : InMux
    port map (
            O => \N__66051\,
            I => \N__65969\
        );

    \I__15669\ : InMux
    port map (
            O => \N__66050\,
            I => \N__65969\
        );

    \I__15668\ : InMux
    port map (
            O => \N__66049\,
            I => \N__65969\
        );

    \I__15667\ : InMux
    port map (
            O => \N__66048\,
            I => \N__65959\
        );

    \I__15666\ : InMux
    port map (
            O => \N__66047\,
            I => \N__65944\
        );

    \I__15665\ : InMux
    port map (
            O => \N__66046\,
            I => \N__65944\
        );

    \I__15664\ : InMux
    port map (
            O => \N__66045\,
            I => \N__65944\
        );

    \I__15663\ : LocalMux
    port map (
            O => \N__66040\,
            I => \N__65937\
        );

    \I__15662\ : LocalMux
    port map (
            O => \N__66037\,
            I => \N__65937\
        );

    \I__15661\ : LocalMux
    port map (
            O => \N__66030\,
            I => \N__65937\
        );

    \I__15660\ : CascadeMux
    port map (
            O => \N__66029\,
            I => \N__65932\
        );

    \I__15659\ : InMux
    port map (
            O => \N__66028\,
            I => \N__65921\
        );

    \I__15658\ : InMux
    port map (
            O => \N__66027\,
            I => \N__65921\
        );

    \I__15657\ : InMux
    port map (
            O => \N__66026\,
            I => \N__65918\
        );

    \I__15656\ : LocalMux
    port map (
            O => \N__66023\,
            I => \N__65911\
        );

    \I__15655\ : LocalMux
    port map (
            O => \N__66020\,
            I => \N__65911\
        );

    \I__15654\ : LocalMux
    port map (
            O => \N__66015\,
            I => \N__65911\
        );

    \I__15653\ : InMux
    port map (
            O => \N__66014\,
            I => \N__65906\
        );

    \I__15652\ : InMux
    port map (
            O => \N__66013\,
            I => \N__65906\
        );

    \I__15651\ : InMux
    port map (
            O => \N__66012\,
            I => \N__65899\
        );

    \I__15650\ : InMux
    port map (
            O => \N__66011\,
            I => \N__65896\
        );

    \I__15649\ : InMux
    port map (
            O => \N__66010\,
            I => \N__65893\
        );

    \I__15648\ : Span4Mux_v
    port map (
            O => \N__66007\,
            I => \N__65890\
        );

    \I__15647\ : LocalMux
    port map (
            O => \N__66000\,
            I => \N__65887\
        );

    \I__15646\ : LocalMux
    port map (
            O => \N__65991\,
            I => \N__65884\
        );

    \I__15645\ : InMux
    port map (
            O => \N__65990\,
            I => \N__65881\
        );

    \I__15644\ : InMux
    port map (
            O => \N__65989\,
            I => \N__65878\
        );

    \I__15643\ : LocalMux
    port map (
            O => \N__65986\,
            I => \N__65873\
        );

    \I__15642\ : LocalMux
    port map (
            O => \N__65981\,
            I => \N__65873\
        );

    \I__15641\ : Span4Mux_h
    port map (
            O => \N__65978\,
            I => \N__65868\
        );

    \I__15640\ : LocalMux
    port map (
            O => \N__65969\,
            I => \N__65868\
        );

    \I__15639\ : InMux
    port map (
            O => \N__65968\,
            I => \N__65861\
        );

    \I__15638\ : InMux
    port map (
            O => \N__65967\,
            I => \N__65861\
        );

    \I__15637\ : InMux
    port map (
            O => \N__65966\,
            I => \N__65861\
        );

    \I__15636\ : InMux
    port map (
            O => \N__65965\,
            I => \N__65852\
        );

    \I__15635\ : InMux
    port map (
            O => \N__65964\,
            I => \N__65852\
        );

    \I__15634\ : InMux
    port map (
            O => \N__65963\,
            I => \N__65852\
        );

    \I__15633\ : InMux
    port map (
            O => \N__65962\,
            I => \N__65852\
        );

    \I__15632\ : LocalMux
    port map (
            O => \N__65959\,
            I => \N__65849\
        );

    \I__15631\ : InMux
    port map (
            O => \N__65958\,
            I => \N__65840\
        );

    \I__15630\ : InMux
    port map (
            O => \N__65957\,
            I => \N__65840\
        );

    \I__15629\ : InMux
    port map (
            O => \N__65956\,
            I => \N__65840\
        );

    \I__15628\ : InMux
    port map (
            O => \N__65955\,
            I => \N__65840\
        );

    \I__15627\ : InMux
    port map (
            O => \N__65954\,
            I => \N__65837\
        );

    \I__15626\ : InMux
    port map (
            O => \N__65953\,
            I => \N__65834\
        );

    \I__15625\ : InMux
    port map (
            O => \N__65952\,
            I => \N__65829\
        );

    \I__15624\ : InMux
    port map (
            O => \N__65951\,
            I => \N__65829\
        );

    \I__15623\ : LocalMux
    port map (
            O => \N__65944\,
            I => \N__65823\
        );

    \I__15622\ : Span4Mux_v
    port map (
            O => \N__65937\,
            I => \N__65820\
        );

    \I__15621\ : InMux
    port map (
            O => \N__65936\,
            I => \N__65817\
        );

    \I__15620\ : InMux
    port map (
            O => \N__65935\,
            I => \N__65814\
        );

    \I__15619\ : InMux
    port map (
            O => \N__65932\,
            I => \N__65811\
        );

    \I__15618\ : InMux
    port map (
            O => \N__65931\,
            I => \N__65808\
        );

    \I__15617\ : InMux
    port map (
            O => \N__65930\,
            I => \N__65805\
        );

    \I__15616\ : InMux
    port map (
            O => \N__65929\,
            I => \N__65802\
        );

    \I__15615\ : CascadeMux
    port map (
            O => \N__65928\,
            I => \N__65799\
        );

    \I__15614\ : InMux
    port map (
            O => \N__65927\,
            I => \N__65794\
        );

    \I__15613\ : InMux
    port map (
            O => \N__65926\,
            I => \N__65794\
        );

    \I__15612\ : LocalMux
    port map (
            O => \N__65921\,
            I => \N__65789\
        );

    \I__15611\ : LocalMux
    port map (
            O => \N__65918\,
            I => \N__65789\
        );

    \I__15610\ : Span4Mux_v
    port map (
            O => \N__65911\,
            I => \N__65784\
        );

    \I__15609\ : LocalMux
    port map (
            O => \N__65906\,
            I => \N__65784\
        );

    \I__15608\ : InMux
    port map (
            O => \N__65905\,
            I => \N__65779\
        );

    \I__15607\ : InMux
    port map (
            O => \N__65904\,
            I => \N__65779\
        );

    \I__15606\ : InMux
    port map (
            O => \N__65903\,
            I => \N__65774\
        );

    \I__15605\ : InMux
    port map (
            O => \N__65902\,
            I => \N__65774\
        );

    \I__15604\ : LocalMux
    port map (
            O => \N__65899\,
            I => \N__65771\
        );

    \I__15603\ : LocalMux
    port map (
            O => \N__65896\,
            I => \N__65766\
        );

    \I__15602\ : LocalMux
    port map (
            O => \N__65893\,
            I => \N__65766\
        );

    \I__15601\ : Span4Mux_h
    port map (
            O => \N__65890\,
            I => \N__65759\
        );

    \I__15600\ : Span4Mux_v
    port map (
            O => \N__65887\,
            I => \N__65759\
        );

    \I__15599\ : Span4Mux_v
    port map (
            O => \N__65884\,
            I => \N__65759\
        );

    \I__15598\ : LocalMux
    port map (
            O => \N__65881\,
            I => \N__65756\
        );

    \I__15597\ : LocalMux
    port map (
            O => \N__65878\,
            I => \N__65750\
        );

    \I__15596\ : Span4Mux_h
    port map (
            O => \N__65873\,
            I => \N__65743\
        );

    \I__15595\ : Span4Mux_v
    port map (
            O => \N__65868\,
            I => \N__65743\
        );

    \I__15594\ : LocalMux
    port map (
            O => \N__65861\,
            I => \N__65743\
        );

    \I__15593\ : LocalMux
    port map (
            O => \N__65852\,
            I => \N__65740\
        );

    \I__15592\ : Span4Mux_h
    port map (
            O => \N__65849\,
            I => \N__65737\
        );

    \I__15591\ : LocalMux
    port map (
            O => \N__65840\,
            I => \N__65734\
        );

    \I__15590\ : LocalMux
    port map (
            O => \N__65837\,
            I => \N__65727\
        );

    \I__15589\ : LocalMux
    port map (
            O => \N__65834\,
            I => \N__65727\
        );

    \I__15588\ : LocalMux
    port map (
            O => \N__65829\,
            I => \N__65727\
        );

    \I__15587\ : InMux
    port map (
            O => \N__65828\,
            I => \N__65724\
        );

    \I__15586\ : CascadeMux
    port map (
            O => \N__65827\,
            I => \N__65721\
        );

    \I__15585\ : CascadeMux
    port map (
            O => \N__65826\,
            I => \N__65712\
        );

    \I__15584\ : Span4Mux_v
    port map (
            O => \N__65823\,
            I => \N__65701\
        );

    \I__15583\ : Span4Mux_h
    port map (
            O => \N__65820\,
            I => \N__65701\
        );

    \I__15582\ : LocalMux
    port map (
            O => \N__65817\,
            I => \N__65701\
        );

    \I__15581\ : LocalMux
    port map (
            O => \N__65814\,
            I => \N__65701\
        );

    \I__15580\ : LocalMux
    port map (
            O => \N__65811\,
            I => \N__65698\
        );

    \I__15579\ : LocalMux
    port map (
            O => \N__65808\,
            I => \N__65695\
        );

    \I__15578\ : LocalMux
    port map (
            O => \N__65805\,
            I => \N__65690\
        );

    \I__15577\ : LocalMux
    port map (
            O => \N__65802\,
            I => \N__65690\
        );

    \I__15576\ : InMux
    port map (
            O => \N__65799\,
            I => \N__65687\
        );

    \I__15575\ : LocalMux
    port map (
            O => \N__65794\,
            I => \N__65676\
        );

    \I__15574\ : Span4Mux_v
    port map (
            O => \N__65789\,
            I => \N__65676\
        );

    \I__15573\ : Span4Mux_h
    port map (
            O => \N__65784\,
            I => \N__65676\
        );

    \I__15572\ : LocalMux
    port map (
            O => \N__65779\,
            I => \N__65676\
        );

    \I__15571\ : LocalMux
    port map (
            O => \N__65774\,
            I => \N__65676\
        );

    \I__15570\ : Span4Mux_v
    port map (
            O => \N__65771\,
            I => \N__65667\
        );

    \I__15569\ : Span4Mux_v
    port map (
            O => \N__65766\,
            I => \N__65667\
        );

    \I__15568\ : Span4Mux_h
    port map (
            O => \N__65759\,
            I => \N__65667\
        );

    \I__15567\ : Span4Mux_v
    port map (
            O => \N__65756\,
            I => \N__65667\
        );

    \I__15566\ : InMux
    port map (
            O => \N__65755\,
            I => \N__65660\
        );

    \I__15565\ : InMux
    port map (
            O => \N__65754\,
            I => \N__65660\
        );

    \I__15564\ : InMux
    port map (
            O => \N__65753\,
            I => \N__65660\
        );

    \I__15563\ : Span4Mux_v
    port map (
            O => \N__65750\,
            I => \N__65655\
        );

    \I__15562\ : Span4Mux_h
    port map (
            O => \N__65743\,
            I => \N__65655\
        );

    \I__15561\ : Span4Mux_v
    port map (
            O => \N__65740\,
            I => \N__65652\
        );

    \I__15560\ : Span4Mux_h
    port map (
            O => \N__65737\,
            I => \N__65647\
        );

    \I__15559\ : Span4Mux_h
    port map (
            O => \N__65734\,
            I => \N__65647\
        );

    \I__15558\ : Span4Mux_h
    port map (
            O => \N__65727\,
            I => \N__65642\
        );

    \I__15557\ : LocalMux
    port map (
            O => \N__65724\,
            I => \N__65642\
        );

    \I__15556\ : InMux
    port map (
            O => \N__65721\,
            I => \N__65635\
        );

    \I__15555\ : InMux
    port map (
            O => \N__65720\,
            I => \N__65635\
        );

    \I__15554\ : InMux
    port map (
            O => \N__65719\,
            I => \N__65635\
        );

    \I__15553\ : InMux
    port map (
            O => \N__65718\,
            I => \N__65628\
        );

    \I__15552\ : InMux
    port map (
            O => \N__65717\,
            I => \N__65628\
        );

    \I__15551\ : InMux
    port map (
            O => \N__65716\,
            I => \N__65628\
        );

    \I__15550\ : InMux
    port map (
            O => \N__65715\,
            I => \N__65619\
        );

    \I__15549\ : InMux
    port map (
            O => \N__65712\,
            I => \N__65619\
        );

    \I__15548\ : InMux
    port map (
            O => \N__65711\,
            I => \N__65619\
        );

    \I__15547\ : InMux
    port map (
            O => \N__65710\,
            I => \N__65619\
        );

    \I__15546\ : Span4Mux_h
    port map (
            O => \N__65701\,
            I => \N__65610\
        );

    \I__15545\ : Span4Mux_v
    port map (
            O => \N__65698\,
            I => \N__65610\
        );

    \I__15544\ : Span4Mux_v
    port map (
            O => \N__65695\,
            I => \N__65610\
        );

    \I__15543\ : Span4Mux_h
    port map (
            O => \N__65690\,
            I => \N__65610\
        );

    \I__15542\ : LocalMux
    port map (
            O => \N__65687\,
            I => \ALU.status_19_0\
        );

    \I__15541\ : Odrv4
    port map (
            O => \N__65676\,
            I => \ALU.status_19_0\
        );

    \I__15540\ : Odrv4
    port map (
            O => \N__65667\,
            I => \ALU.status_19_0\
        );

    \I__15539\ : LocalMux
    port map (
            O => \N__65660\,
            I => \ALU.status_19_0\
        );

    \I__15538\ : Odrv4
    port map (
            O => \N__65655\,
            I => \ALU.status_19_0\
        );

    \I__15537\ : Odrv4
    port map (
            O => \N__65652\,
            I => \ALU.status_19_0\
        );

    \I__15536\ : Odrv4
    port map (
            O => \N__65647\,
            I => \ALU.status_19_0\
        );

    \I__15535\ : Odrv4
    port map (
            O => \N__65642\,
            I => \ALU.status_19_0\
        );

    \I__15534\ : LocalMux
    port map (
            O => \N__65635\,
            I => \ALU.status_19_0\
        );

    \I__15533\ : LocalMux
    port map (
            O => \N__65628\,
            I => \ALU.status_19_0\
        );

    \I__15532\ : LocalMux
    port map (
            O => \N__65619\,
            I => \ALU.status_19_0\
        );

    \I__15531\ : Odrv4
    port map (
            O => \N__65610\,
            I => \ALU.status_19_0\
        );

    \I__15530\ : CascadeMux
    port map (
            O => \N__65585\,
            I => \N__65581\
        );

    \I__15529\ : InMux
    port map (
            O => \N__65584\,
            I => \N__65576\
        );

    \I__15528\ : InMux
    port map (
            O => \N__65581\,
            I => \N__65576\
        );

    \I__15527\ : LocalMux
    port map (
            O => \N__65576\,
            I => \N__65571\
        );

    \I__15526\ : CascadeMux
    port map (
            O => \N__65575\,
            I => \N__65566\
        );

    \I__15525\ : CascadeMux
    port map (
            O => \N__65574\,
            I => \N__65559\
        );

    \I__15524\ : Span4Mux_v
    port map (
            O => \N__65571\,
            I => \N__65553\
        );

    \I__15523\ : InMux
    port map (
            O => \N__65570\,
            I => \N__65547\
        );

    \I__15522\ : InMux
    port map (
            O => \N__65569\,
            I => \N__65531\
        );

    \I__15521\ : InMux
    port map (
            O => \N__65566\,
            I => \N__65531\
        );

    \I__15520\ : InMux
    port map (
            O => \N__65565\,
            I => \N__65528\
        );

    \I__15519\ : CascadeMux
    port map (
            O => \N__65564\,
            I => \N__65523\
        );

    \I__15518\ : InMux
    port map (
            O => \N__65563\,
            I => \N__65517\
        );

    \I__15517\ : InMux
    port map (
            O => \N__65562\,
            I => \N__65514\
        );

    \I__15516\ : InMux
    port map (
            O => \N__65559\,
            I => \N__65511\
        );

    \I__15515\ : InMux
    port map (
            O => \N__65558\,
            I => \N__65508\
        );

    \I__15514\ : InMux
    port map (
            O => \N__65557\,
            I => \N__65505\
        );

    \I__15513\ : InMux
    port map (
            O => \N__65556\,
            I => \N__65502\
        );

    \I__15512\ : Span4Mux_h
    port map (
            O => \N__65553\,
            I => \N__65499\
        );

    \I__15511\ : InMux
    port map (
            O => \N__65552\,
            I => \N__65494\
        );

    \I__15510\ : InMux
    port map (
            O => \N__65551\,
            I => \N__65494\
        );

    \I__15509\ : InMux
    port map (
            O => \N__65550\,
            I => \N__65490\
        );

    \I__15508\ : LocalMux
    port map (
            O => \N__65547\,
            I => \N__65487\
        );

    \I__15507\ : CascadeMux
    port map (
            O => \N__65546\,
            I => \N__65484\
        );

    \I__15506\ : InMux
    port map (
            O => \N__65545\,
            I => \N__65474\
        );

    \I__15505\ : InMux
    port map (
            O => \N__65544\,
            I => \N__65474\
        );

    \I__15504\ : InMux
    port map (
            O => \N__65543\,
            I => \N__65469\
        );

    \I__15503\ : InMux
    port map (
            O => \N__65542\,
            I => \N__65469\
        );

    \I__15502\ : InMux
    port map (
            O => \N__65541\,
            I => \N__65464\
        );

    \I__15501\ : InMux
    port map (
            O => \N__65540\,
            I => \N__65464\
        );

    \I__15500\ : InMux
    port map (
            O => \N__65539\,
            I => \N__65461\
        );

    \I__15499\ : InMux
    port map (
            O => \N__65538\,
            I => \N__65458\
        );

    \I__15498\ : InMux
    port map (
            O => \N__65537\,
            I => \N__65455\
        );

    \I__15497\ : InMux
    port map (
            O => \N__65536\,
            I => \N__65452\
        );

    \I__15496\ : LocalMux
    port map (
            O => \N__65531\,
            I => \N__65447\
        );

    \I__15495\ : LocalMux
    port map (
            O => \N__65528\,
            I => \N__65447\
        );

    \I__15494\ : InMux
    port map (
            O => \N__65527\,
            I => \N__65439\
        );

    \I__15493\ : InMux
    port map (
            O => \N__65526\,
            I => \N__65439\
        );

    \I__15492\ : InMux
    port map (
            O => \N__65523\,
            I => \N__65434\
        );

    \I__15491\ : InMux
    port map (
            O => \N__65522\,
            I => \N__65434\
        );

    \I__15490\ : InMux
    port map (
            O => \N__65521\,
            I => \N__65431\
        );

    \I__15489\ : InMux
    port map (
            O => \N__65520\,
            I => \N__65428\
        );

    \I__15488\ : LocalMux
    port map (
            O => \N__65517\,
            I => \N__65423\
        );

    \I__15487\ : LocalMux
    port map (
            O => \N__65514\,
            I => \N__65423\
        );

    \I__15486\ : LocalMux
    port map (
            O => \N__65511\,
            I => \N__65418\
        );

    \I__15485\ : LocalMux
    port map (
            O => \N__65508\,
            I => \N__65418\
        );

    \I__15484\ : LocalMux
    port map (
            O => \N__65505\,
            I => \N__65409\
        );

    \I__15483\ : LocalMux
    port map (
            O => \N__65502\,
            I => \N__65409\
        );

    \I__15482\ : Span4Mux_v
    port map (
            O => \N__65499\,
            I => \N__65409\
        );

    \I__15481\ : LocalMux
    port map (
            O => \N__65494\,
            I => \N__65409\
        );

    \I__15480\ : InMux
    port map (
            O => \N__65493\,
            I => \N__65404\
        );

    \I__15479\ : LocalMux
    port map (
            O => \N__65490\,
            I => \N__65399\
        );

    \I__15478\ : Span4Mux_h
    port map (
            O => \N__65487\,
            I => \N__65399\
        );

    \I__15477\ : InMux
    port map (
            O => \N__65484\,
            I => \N__65386\
        );

    \I__15476\ : InMux
    port map (
            O => \N__65483\,
            I => \N__65386\
        );

    \I__15475\ : InMux
    port map (
            O => \N__65482\,
            I => \N__65386\
        );

    \I__15474\ : InMux
    port map (
            O => \N__65481\,
            I => \N__65386\
        );

    \I__15473\ : InMux
    port map (
            O => \N__65480\,
            I => \N__65386\
        );

    \I__15472\ : InMux
    port map (
            O => \N__65479\,
            I => \N__65386\
        );

    \I__15471\ : LocalMux
    port map (
            O => \N__65474\,
            I => \N__65379\
        );

    \I__15470\ : LocalMux
    port map (
            O => \N__65469\,
            I => \N__65379\
        );

    \I__15469\ : LocalMux
    port map (
            O => \N__65464\,
            I => \N__65379\
        );

    \I__15468\ : LocalMux
    port map (
            O => \N__65461\,
            I => \N__65374\
        );

    \I__15467\ : LocalMux
    port map (
            O => \N__65458\,
            I => \N__65374\
        );

    \I__15466\ : LocalMux
    port map (
            O => \N__65455\,
            I => \N__65369\
        );

    \I__15465\ : LocalMux
    port map (
            O => \N__65452\,
            I => \N__65369\
        );

    \I__15464\ : Span4Mux_v
    port map (
            O => \N__65447\,
            I => \N__65366\
        );

    \I__15463\ : InMux
    port map (
            O => \N__65446\,
            I => \N__65359\
        );

    \I__15462\ : InMux
    port map (
            O => \N__65445\,
            I => \N__65359\
        );

    \I__15461\ : InMux
    port map (
            O => \N__65444\,
            I => \N__65359\
        );

    \I__15460\ : LocalMux
    port map (
            O => \N__65439\,
            I => \N__65352\
        );

    \I__15459\ : LocalMux
    port map (
            O => \N__65434\,
            I => \N__65352\
        );

    \I__15458\ : LocalMux
    port map (
            O => \N__65431\,
            I => \N__65352\
        );

    \I__15457\ : LocalMux
    port map (
            O => \N__65428\,
            I => \N__65348\
        );

    \I__15456\ : Span4Mux_v
    port map (
            O => \N__65423\,
            I => \N__65343\
        );

    \I__15455\ : Span4Mux_v
    port map (
            O => \N__65418\,
            I => \N__65343\
        );

    \I__15454\ : Span4Mux_h
    port map (
            O => \N__65409\,
            I => \N__65340\
        );

    \I__15453\ : InMux
    port map (
            O => \N__65408\,
            I => \N__65335\
        );

    \I__15452\ : InMux
    port map (
            O => \N__65407\,
            I => \N__65335\
        );

    \I__15451\ : LocalMux
    port map (
            O => \N__65404\,
            I => \N__65326\
        );

    \I__15450\ : Span4Mux_v
    port map (
            O => \N__65399\,
            I => \N__65326\
        );

    \I__15449\ : LocalMux
    port map (
            O => \N__65386\,
            I => \N__65326\
        );

    \I__15448\ : Span4Mux_h
    port map (
            O => \N__65379\,
            I => \N__65326\
        );

    \I__15447\ : Span12Mux_v
    port map (
            O => \N__65374\,
            I => \N__65319\
        );

    \I__15446\ : Span12Mux_v
    port map (
            O => \N__65369\,
            I => \N__65319\
        );

    \I__15445\ : Sp12to4
    port map (
            O => \N__65366\,
            I => \N__65319\
        );

    \I__15444\ : LocalMux
    port map (
            O => \N__65359\,
            I => \N__65316\
        );

    \I__15443\ : Span4Mux_v
    port map (
            O => \N__65352\,
            I => \N__65313\
        );

    \I__15442\ : InMux
    port map (
            O => \N__65351\,
            I => \N__65310\
        );

    \I__15441\ : Span4Mux_v
    port map (
            O => \N__65348\,
            I => \N__65305\
        );

    \I__15440\ : Span4Mux_h
    port map (
            O => \N__65343\,
            I => \N__65305\
        );

    \I__15439\ : Span4Mux_v
    port map (
            O => \N__65340\,
            I => \N__65298\
        );

    \I__15438\ : LocalMux
    port map (
            O => \N__65335\,
            I => \N__65298\
        );

    \I__15437\ : Span4Mux_v
    port map (
            O => \N__65326\,
            I => \N__65298\
        );

    \I__15436\ : Odrv12
    port map (
            O => \N__65319\,
            I => \aluOut_1\
        );

    \I__15435\ : Odrv12
    port map (
            O => \N__65316\,
            I => \aluOut_1\
        );

    \I__15434\ : Odrv4
    port map (
            O => \N__65313\,
            I => \aluOut_1\
        );

    \I__15433\ : LocalMux
    port map (
            O => \N__65310\,
            I => \aluOut_1\
        );

    \I__15432\ : Odrv4
    port map (
            O => \N__65305\,
            I => \aluOut_1\
        );

    \I__15431\ : Odrv4
    port map (
            O => \N__65298\,
            I => \aluOut_1\
        );

    \I__15430\ : InMux
    port map (
            O => \N__65285\,
            I => \N__65282\
        );

    \I__15429\ : LocalMux
    port map (
            O => \N__65282\,
            I => \ALU.d_RNIMGKJC1_0Z0Z_2\
        );

    \I__15428\ : CascadeMux
    port map (
            O => \N__65279\,
            I => \ALU.d_RNIMGKJC1Z0Z_2_cascade_\
        );

    \I__15427\ : InMux
    port map (
            O => \N__65276\,
            I => \N__65273\
        );

    \I__15426\ : LocalMux
    port map (
            O => \N__65273\,
            I => \N__65269\
        );

    \I__15425\ : InMux
    port map (
            O => \N__65272\,
            I => \N__65266\
        );

    \I__15424\ : Span4Mux_v
    port map (
            O => \N__65269\,
            I => \N__65263\
        );

    \I__15423\ : LocalMux
    port map (
            O => \N__65266\,
            I => \N__65260\
        );

    \I__15422\ : Sp12to4
    port map (
            O => \N__65263\,
            I => \N__65255\
        );

    \I__15421\ : Span12Mux_s9_h
    port map (
            O => \N__65260\,
            I => \N__65255\
        );

    \I__15420\ : Span12Mux_h
    port map (
            O => \N__65255\,
            I => \N__65252\
        );

    \I__15419\ : Odrv12
    port map (
            O => \N__65252\,
            I => \ALU.N_831\
        );

    \I__15418\ : InMux
    port map (
            O => \N__65249\,
            I => \N__65246\
        );

    \I__15417\ : LocalMux
    port map (
            O => \N__65246\,
            I => \N__65243\
        );

    \I__15416\ : Odrv4
    port map (
            O => \N__65243\,
            I => \PROM.ROMDATA.m427_bm\
        );

    \I__15415\ : CascadeMux
    port map (
            O => \N__65240\,
            I => \PROM.ROMDATA.m427_am_cascade_\
        );

    \I__15414\ : CascadeMux
    port map (
            O => \N__65237\,
            I => \N__65233\
        );

    \I__15413\ : InMux
    port map (
            O => \N__65236\,
            I => \N__65228\
        );

    \I__15412\ : InMux
    port map (
            O => \N__65233\,
            I => \N__65228\
        );

    \I__15411\ : LocalMux
    port map (
            O => \N__65228\,
            I => \N__65225\
        );

    \I__15410\ : Span4Mux_v
    port map (
            O => \N__65225\,
            I => \N__65222\
        );

    \I__15409\ : Sp12to4
    port map (
            O => \N__65222\,
            I => \N__65219\
        );

    \I__15408\ : Span12Mux_h
    port map (
            O => \N__65219\,
            I => \N__65216\
        );

    \I__15407\ : Odrv12
    port map (
            O => \N__65216\,
            I => \PROM.ROMDATA.m427_ns\
        );

    \I__15406\ : InMux
    port map (
            O => \N__65213\,
            I => \N__65210\
        );

    \I__15405\ : LocalMux
    port map (
            O => \N__65210\,
            I => \N__65207\
        );

    \I__15404\ : Span4Mux_h
    port map (
            O => \N__65207\,
            I => \N__65204\
        );

    \I__15403\ : Odrv4
    port map (
            O => \N__65204\,
            I => \PROM.ROMDATA.m492_am\
        );

    \I__15402\ : CascadeMux
    port map (
            O => \N__65201\,
            I => \N__65198\
        );

    \I__15401\ : InMux
    port map (
            O => \N__65198\,
            I => \N__65195\
        );

    \I__15400\ : LocalMux
    port map (
            O => \N__65195\,
            I => \PROM.ROMDATA.m492_bm\
        );

    \I__15399\ : InMux
    port map (
            O => \N__65192\,
            I => \N__65189\
        );

    \I__15398\ : LocalMux
    port map (
            O => \N__65189\,
            I => \N__65186\
        );

    \I__15397\ : Odrv12
    port map (
            O => \N__65186\,
            I => \PROM.ROMDATA.m494_ns_1\
        );

    \I__15396\ : InMux
    port map (
            O => \N__65183\,
            I => \N__65180\
        );

    \I__15395\ : LocalMux
    port map (
            O => \N__65180\,
            I => \N__65177\
        );

    \I__15394\ : Span4Mux_h
    port map (
            O => \N__65177\,
            I => \N__65174\
        );

    \I__15393\ : Odrv4
    port map (
            O => \N__65174\,
            I => \PROM.ROMDATA.m88\
        );

    \I__15392\ : InMux
    port map (
            O => \N__65171\,
            I => \N__65168\
        );

    \I__15391\ : LocalMux
    port map (
            O => \N__65168\,
            I => \N__65165\
        );

    \I__15390\ : Span4Mux_v
    port map (
            O => \N__65165\,
            I => \N__65162\
        );

    \I__15389\ : Sp12to4
    port map (
            O => \N__65162\,
            I => \N__65159\
        );

    \I__15388\ : Span12Mux_h
    port map (
            O => \N__65159\,
            I => \N__65156\
        );

    \I__15387\ : Odrv12
    port map (
            O => \N__65156\,
            I => \PROM.ROMDATA.m514_ns_1\
        );

    \I__15386\ : CascadeMux
    port map (
            O => \N__65153\,
            I => \PROM.ROMDATA.m181_cascade_\
        );

    \I__15385\ : InMux
    port map (
            O => \N__65150\,
            I => \N__65146\
        );

    \I__15384\ : CascadeMux
    port map (
            O => \N__65149\,
            I => \N__65143\
        );

    \I__15383\ : LocalMux
    port map (
            O => \N__65146\,
            I => \N__65140\
        );

    \I__15382\ : InMux
    port map (
            O => \N__65143\,
            I => \N__65137\
        );

    \I__15381\ : Span4Mux_v
    port map (
            O => \N__65140\,
            I => \N__65134\
        );

    \I__15380\ : LocalMux
    port map (
            O => \N__65137\,
            I => \N__65131\
        );

    \I__15379\ : Span4Mux_v
    port map (
            O => \N__65134\,
            I => \N__65126\
        );

    \I__15378\ : Span4Mux_h
    port map (
            O => \N__65131\,
            I => \N__65126\
        );

    \I__15377\ : Span4Mux_h
    port map (
            O => \N__65126\,
            I => \N__65123\
        );

    \I__15376\ : Span4Mux_v
    port map (
            O => \N__65123\,
            I => \N__65120\
        );

    \I__15375\ : Span4Mux_h
    port map (
            O => \N__65120\,
            I => \N__65117\
        );

    \I__15374\ : Odrv4
    port map (
            O => \N__65117\,
            I => \PROM.ROMDATA.m514_ns\
        );

    \I__15373\ : InMux
    port map (
            O => \N__65114\,
            I => \N__65111\
        );

    \I__15372\ : LocalMux
    port map (
            O => \N__65111\,
            I => \PROM.ROMDATA.N_525_mux\
        );

    \I__15371\ : InMux
    port map (
            O => \N__65108\,
            I => \N__65105\
        );

    \I__15370\ : LocalMux
    port map (
            O => \N__65105\,
            I => \PROM.ROMDATA.m164\
        );

    \I__15369\ : InMux
    port map (
            O => \N__65102\,
            I => \N__65099\
        );

    \I__15368\ : LocalMux
    port map (
            O => \N__65099\,
            I => \PROM.ROMDATA.m171_am\
        );

    \I__15367\ : InMux
    port map (
            O => \N__65096\,
            I => \N__65093\
        );

    \I__15366\ : LocalMux
    port map (
            O => \N__65093\,
            I => \N__65090\
        );

    \I__15365\ : Span4Mux_v
    port map (
            O => \N__65090\,
            I => \N__65086\
        );

    \I__15364\ : InMux
    port map (
            O => \N__65089\,
            I => \N__65083\
        );

    \I__15363\ : Span4Mux_h
    port map (
            O => \N__65086\,
            I => \N__65078\
        );

    \I__15362\ : LocalMux
    port map (
            O => \N__65083\,
            I => \N__65078\
        );

    \I__15361\ : Span4Mux_v
    port map (
            O => \N__65078\,
            I => \N__65075\
        );

    \I__15360\ : Span4Mux_h
    port map (
            O => \N__65075\,
            I => \N__65072\
        );

    \I__15359\ : Span4Mux_h
    port map (
            O => \N__65072\,
            I => \N__65069\
        );

    \I__15358\ : Span4Mux_h
    port map (
            O => \N__65069\,
            I => \N__65066\
        );

    \I__15357\ : Span4Mux_v
    port map (
            O => \N__65066\,
            I => \N__65063\
        );

    \I__15356\ : Odrv4
    port map (
            O => \N__65063\,
            I => \ALU.dZ0Z_12\
        );

    \I__15355\ : InMux
    port map (
            O => \N__65060\,
            I => \N__65057\
        );

    \I__15354\ : LocalMux
    port map (
            O => \N__65057\,
            I => \N__65053\
        );

    \I__15353\ : InMux
    port map (
            O => \N__65056\,
            I => \N__65050\
        );

    \I__15352\ : Span4Mux_v
    port map (
            O => \N__65053\,
            I => \N__65047\
        );

    \I__15351\ : LocalMux
    port map (
            O => \N__65050\,
            I => \N__65044\
        );

    \I__15350\ : Span4Mux_h
    port map (
            O => \N__65047\,
            I => \N__65041\
        );

    \I__15349\ : Span12Mux_h
    port map (
            O => \N__65044\,
            I => \N__65038\
        );

    \I__15348\ : Odrv4
    port map (
            O => \N__65041\,
            I => \ALU.dZ0Z_13\
        );

    \I__15347\ : Odrv12
    port map (
            O => \N__65038\,
            I => \ALU.dZ0Z_13\
        );

    \I__15346\ : CascadeMux
    port map (
            O => \N__65033\,
            I => \N__65030\
        );

    \I__15345\ : InMux
    port map (
            O => \N__65030\,
            I => \N__65026\
        );

    \I__15344\ : CascadeMux
    port map (
            O => \N__65029\,
            I => \N__65023\
        );

    \I__15343\ : LocalMux
    port map (
            O => \N__65026\,
            I => \N__65020\
        );

    \I__15342\ : InMux
    port map (
            O => \N__65023\,
            I => \N__65017\
        );

    \I__15341\ : Span4Mux_v
    port map (
            O => \N__65020\,
            I => \N__65014\
        );

    \I__15340\ : LocalMux
    port map (
            O => \N__65017\,
            I => \N__65010\
        );

    \I__15339\ : Span4Mux_h
    port map (
            O => \N__65014\,
            I => \N__65007\
        );

    \I__15338\ : InMux
    port map (
            O => \N__65013\,
            I => \N__65004\
        );

    \I__15337\ : Span4Mux_v
    port map (
            O => \N__65010\,
            I => \N__65001\
        );

    \I__15336\ : Span4Mux_h
    port map (
            O => \N__65007\,
            I => \N__64998\
        );

    \I__15335\ : LocalMux
    port map (
            O => \N__65004\,
            I => \N__64995\
        );

    \I__15334\ : Span4Mux_h
    port map (
            O => \N__65001\,
            I => \N__64992\
        );

    \I__15333\ : Span4Mux_h
    port map (
            O => \N__64998\,
            I => \N__64989\
        );

    \I__15332\ : Span4Mux_v
    port map (
            O => \N__64995\,
            I => \N__64984\
        );

    \I__15331\ : Span4Mux_h
    port map (
            O => \N__64992\,
            I => \N__64984\
        );

    \I__15330\ : Span4Mux_h
    port map (
            O => \N__64989\,
            I => \N__64981\
        );

    \I__15329\ : Odrv4
    port map (
            O => \N__64984\,
            I => \PROM.ROMDATA.m83\
        );

    \I__15328\ : Odrv4
    port map (
            O => \N__64981\,
            I => \PROM.ROMDATA.m83\
        );

    \I__15327\ : CascadeMux
    port map (
            O => \N__64976\,
            I => \PROM.ROMDATA.m83_cascade_\
        );

    \I__15326\ : InMux
    port map (
            O => \N__64973\,
            I => \N__64970\
        );

    \I__15325\ : LocalMux
    port map (
            O => \N__64970\,
            I => \N__64967\
        );

    \I__15324\ : Span4Mux_h
    port map (
            O => \N__64967\,
            I => \N__64961\
        );

    \I__15323\ : InMux
    port map (
            O => \N__64966\,
            I => \N__64958\
        );

    \I__15322\ : InMux
    port map (
            O => \N__64965\,
            I => \N__64955\
        );

    \I__15321\ : InMux
    port map (
            O => \N__64964\,
            I => \N__64952\
        );

    \I__15320\ : Span4Mux_h
    port map (
            O => \N__64961\,
            I => \N__64949\
        );

    \I__15319\ : LocalMux
    port map (
            O => \N__64958\,
            I => \N__64946\
        );

    \I__15318\ : LocalMux
    port map (
            O => \N__64955\,
            I => \N__64941\
        );

    \I__15317\ : LocalMux
    port map (
            O => \N__64952\,
            I => \N__64941\
        );

    \I__15316\ : Span4Mux_h
    port map (
            O => \N__64949\,
            I => \N__64933\
        );

    \I__15315\ : Span4Mux_h
    port map (
            O => \N__64946\,
            I => \N__64933\
        );

    \I__15314\ : Span4Mux_h
    port map (
            O => \N__64941\,
            I => \N__64933\
        );

    \I__15313\ : InMux
    port map (
            O => \N__64940\,
            I => \N__64930\
        );

    \I__15312\ : Odrv4
    port map (
            O => \N__64933\,
            I => \PROM.ROMDATA.m133\
        );

    \I__15311\ : LocalMux
    port map (
            O => \N__64930\,
            I => \PROM.ROMDATA.m133\
        );

    \I__15310\ : InMux
    port map (
            O => \N__64925\,
            I => \N__64922\
        );

    \I__15309\ : LocalMux
    port map (
            O => \N__64922\,
            I => \PROM.ROMDATA.m161\
        );

    \I__15308\ : InMux
    port map (
            O => \N__64919\,
            I => \N__64916\
        );

    \I__15307\ : LocalMux
    port map (
            O => \N__64916\,
            I => \PROM.ROMDATA.m15\
        );

    \I__15306\ : CascadeMux
    port map (
            O => \N__64913\,
            I => \PROM.ROMDATA.m171_ns_cascade_\
        );

    \I__15305\ : InMux
    port map (
            O => \N__64910\,
            I => \N__64907\
        );

    \I__15304\ : LocalMux
    port map (
            O => \N__64907\,
            I => \PROM.ROMDATA.m162\
        );

    \I__15303\ : InMux
    port map (
            O => \N__64904\,
            I => \N__64901\
        );

    \I__15302\ : LocalMux
    port map (
            O => \N__64901\,
            I => \N__64897\
        );

    \I__15301\ : InMux
    port map (
            O => \N__64900\,
            I => \N__64894\
        );

    \I__15300\ : Span4Mux_h
    port map (
            O => \N__64897\,
            I => \N__64891\
        );

    \I__15299\ : LocalMux
    port map (
            O => \N__64894\,
            I => \N__64888\
        );

    \I__15298\ : Span4Mux_h
    port map (
            O => \N__64891\,
            I => \N__64885\
        );

    \I__15297\ : Span4Mux_h
    port map (
            O => \N__64888\,
            I => \N__64882\
        );

    \I__15296\ : Odrv4
    port map (
            O => \N__64885\,
            I => \PROM.ROMDATA.m172\
        );

    \I__15295\ : Odrv4
    port map (
            O => \N__64882\,
            I => \PROM.ROMDATA.m172\
        );

    \I__15294\ : InMux
    port map (
            O => \N__64877\,
            I => \N__64872\
        );

    \I__15293\ : CascadeMux
    port map (
            O => \N__64876\,
            I => \N__64867\
        );

    \I__15292\ : CascadeMux
    port map (
            O => \N__64875\,
            I => \N__64864\
        );

    \I__15291\ : LocalMux
    port map (
            O => \N__64872\,
            I => \N__64858\
        );

    \I__15290\ : CascadeMux
    port map (
            O => \N__64871\,
            I => \N__64855\
        );

    \I__15289\ : InMux
    port map (
            O => \N__64870\,
            I => \N__64852\
        );

    \I__15288\ : InMux
    port map (
            O => \N__64867\,
            I => \N__64849\
        );

    \I__15287\ : InMux
    port map (
            O => \N__64864\,
            I => \N__64844\
        );

    \I__15286\ : InMux
    port map (
            O => \N__64863\,
            I => \N__64844\
        );

    \I__15285\ : InMux
    port map (
            O => \N__64862\,
            I => \N__64841\
        );

    \I__15284\ : CascadeMux
    port map (
            O => \N__64861\,
            I => \N__64838\
        );

    \I__15283\ : Span4Mux_v
    port map (
            O => \N__64858\,
            I => \N__64834\
        );

    \I__15282\ : InMux
    port map (
            O => \N__64855\,
            I => \N__64831\
        );

    \I__15281\ : LocalMux
    port map (
            O => \N__64852\,
            I => \N__64828\
        );

    \I__15280\ : LocalMux
    port map (
            O => \N__64849\,
            I => \N__64825\
        );

    \I__15279\ : LocalMux
    port map (
            O => \N__64844\,
            I => \N__64822\
        );

    \I__15278\ : LocalMux
    port map (
            O => \N__64841\,
            I => \N__64819\
        );

    \I__15277\ : InMux
    port map (
            O => \N__64838\,
            I => \N__64814\
        );

    \I__15276\ : InMux
    port map (
            O => \N__64837\,
            I => \N__64814\
        );

    \I__15275\ : Span4Mux_h
    port map (
            O => \N__64834\,
            I => \N__64809\
        );

    \I__15274\ : LocalMux
    port map (
            O => \N__64831\,
            I => \N__64809\
        );

    \I__15273\ : Span4Mux_v
    port map (
            O => \N__64828\,
            I => \N__64804\
        );

    \I__15272\ : Span4Mux_h
    port map (
            O => \N__64825\,
            I => \N__64804\
        );

    \I__15271\ : Odrv12
    port map (
            O => \N__64822\,
            I => \PROM.ROMDATA.m20\
        );

    \I__15270\ : Odrv12
    port map (
            O => \N__64819\,
            I => \PROM.ROMDATA.m20\
        );

    \I__15269\ : LocalMux
    port map (
            O => \N__64814\,
            I => \PROM.ROMDATA.m20\
        );

    \I__15268\ : Odrv4
    port map (
            O => \N__64809\,
            I => \PROM.ROMDATA.m20\
        );

    \I__15267\ : Odrv4
    port map (
            O => \N__64804\,
            I => \PROM.ROMDATA.m20\
        );

    \I__15266\ : InMux
    port map (
            O => \N__64793\,
            I => \N__64790\
        );

    \I__15265\ : LocalMux
    port map (
            O => \N__64790\,
            I => \N__64786\
        );

    \I__15264\ : InMux
    port map (
            O => \N__64789\,
            I => \N__64783\
        );

    \I__15263\ : Odrv4
    port map (
            O => \N__64786\,
            I => \PROM.ROMDATA.m156\
        );

    \I__15262\ : LocalMux
    port map (
            O => \N__64783\,
            I => \PROM.ROMDATA.m156\
        );

    \I__15261\ : InMux
    port map (
            O => \N__64778\,
            I => \N__64775\
        );

    \I__15260\ : LocalMux
    port map (
            O => \N__64775\,
            I => \PROM.ROMDATA.m171_bm\
        );

    \I__15259\ : CascadeMux
    port map (
            O => \N__64772\,
            I => \PROM.ROMDATA.m383_cascade_\
        );

    \I__15258\ : InMux
    port map (
            O => \N__64769\,
            I => \N__64766\
        );

    \I__15257\ : LocalMux
    port map (
            O => \N__64766\,
            I => \PROM.ROMDATA.m140\
        );

    \I__15256\ : CascadeMux
    port map (
            O => \N__64763\,
            I => \PROM.ROMDATA.m138_cascade_\
        );

    \I__15255\ : CascadeMux
    port map (
            O => \N__64760\,
            I => \PROM.ROMDATA.m80_bm_1_cascade_\
        );

    \I__15254\ : InMux
    port map (
            O => \N__64757\,
            I => \N__64754\
        );

    \I__15253\ : LocalMux
    port map (
            O => \N__64754\,
            I => \N__64751\
        );

    \I__15252\ : Odrv4
    port map (
            O => \N__64751\,
            I => \PROM.ROMDATA.m80_bm\
        );

    \I__15251\ : InMux
    port map (
            O => \N__64748\,
            I => \N__64742\
        );

    \I__15250\ : InMux
    port map (
            O => \N__64747\,
            I => \N__64742\
        );

    \I__15249\ : LocalMux
    port map (
            O => \N__64742\,
            I => \N__64737\
        );

    \I__15248\ : InMux
    port map (
            O => \N__64741\,
            I => \N__64734\
        );

    \I__15247\ : InMux
    port map (
            O => \N__64740\,
            I => \N__64731\
        );

    \I__15246\ : Span4Mux_h
    port map (
            O => \N__64737\,
            I => \N__64728\
        );

    \I__15245\ : LocalMux
    port map (
            O => \N__64734\,
            I => \N__64725\
        );

    \I__15244\ : LocalMux
    port map (
            O => \N__64731\,
            I => \N__64722\
        );

    \I__15243\ : Odrv4
    port map (
            O => \N__64728\,
            I => \N_417\
        );

    \I__15242\ : Odrv4
    port map (
            O => \N__64725\,
            I => \N_417\
        );

    \I__15241\ : Odrv12
    port map (
            O => \N__64722\,
            I => \N_417\
        );

    \I__15240\ : CascadeMux
    port map (
            O => \N__64715\,
            I => \N__64712\
        );

    \I__15239\ : InMux
    port map (
            O => \N__64712\,
            I => \N__64705\
        );

    \I__15238\ : InMux
    port map (
            O => \N__64711\,
            I => \N__64705\
        );

    \I__15237\ : InMux
    port map (
            O => \N__64710\,
            I => \N__64702\
        );

    \I__15236\ : LocalMux
    port map (
            O => \N__64705\,
            I => \N__64699\
        );

    \I__15235\ : LocalMux
    port map (
            O => \N__64702\,
            I => \N__64695\
        );

    \I__15234\ : Span4Mux_h
    port map (
            O => \N__64699\,
            I => \N__64689\
        );

    \I__15233\ : InMux
    port map (
            O => \N__64698\,
            I => \N__64686\
        );

    \I__15232\ : Span4Mux_v
    port map (
            O => \N__64695\,
            I => \N__64683\
        );

    \I__15231\ : InMux
    port map (
            O => \N__64694\,
            I => \N__64680\
        );

    \I__15230\ : InMux
    port map (
            O => \N__64693\,
            I => \N__64675\
        );

    \I__15229\ : InMux
    port map (
            O => \N__64692\,
            I => \N__64675\
        );

    \I__15228\ : Odrv4
    port map (
            O => \N__64689\,
            I => \CONTROL_addrstack_reto_2\
        );

    \I__15227\ : LocalMux
    port map (
            O => \N__64686\,
            I => \CONTROL_addrstack_reto_2\
        );

    \I__15226\ : Odrv4
    port map (
            O => \N__64683\,
            I => \CONTROL_addrstack_reto_2\
        );

    \I__15225\ : LocalMux
    port map (
            O => \N__64680\,
            I => \CONTROL_addrstack_reto_2\
        );

    \I__15224\ : LocalMux
    port map (
            O => \N__64675\,
            I => \CONTROL_addrstack_reto_2\
        );

    \I__15223\ : InMux
    port map (
            O => \N__64664\,
            I => \N__64659\
        );

    \I__15222\ : InMux
    port map (
            O => \N__64663\,
            I => \N__64656\
        );

    \I__15221\ : CascadeMux
    port map (
            O => \N__64662\,
            I => \N__64652\
        );

    \I__15220\ : LocalMux
    port map (
            O => \N__64659\,
            I => \N__64649\
        );

    \I__15219\ : LocalMux
    port map (
            O => \N__64656\,
            I => \N__64646\
        );

    \I__15218\ : InMux
    port map (
            O => \N__64655\,
            I => \N__64643\
        );

    \I__15217\ : InMux
    port map (
            O => \N__64652\,
            I => \N__64638\
        );

    \I__15216\ : Span4Mux_v
    port map (
            O => \N__64649\,
            I => \N__64635\
        );

    \I__15215\ : Span4Mux_v
    port map (
            O => \N__64646\,
            I => \N__64632\
        );

    \I__15214\ : LocalMux
    port map (
            O => \N__64643\,
            I => \N__64629\
        );

    \I__15213\ : InMux
    port map (
            O => \N__64642\,
            I => \N__64626\
        );

    \I__15212\ : CascadeMux
    port map (
            O => \N__64641\,
            I => \N__64623\
        );

    \I__15211\ : LocalMux
    port map (
            O => \N__64638\,
            I => \N__64620\
        );

    \I__15210\ : Span4Mux_v
    port map (
            O => \N__64635\,
            I => \N__64616\
        );

    \I__15209\ : Span4Mux_v
    port map (
            O => \N__64632\,
            I => \N__64611\
        );

    \I__15208\ : Span4Mux_v
    port map (
            O => \N__64629\,
            I => \N__64611\
        );

    \I__15207\ : LocalMux
    port map (
            O => \N__64626\,
            I => \N__64608\
        );

    \I__15206\ : InMux
    port map (
            O => \N__64623\,
            I => \N__64605\
        );

    \I__15205\ : Span4Mux_h
    port map (
            O => \N__64620\,
            I => \N__64602\
        );

    \I__15204\ : InMux
    port map (
            O => \N__64619\,
            I => \N__64599\
        );

    \I__15203\ : Span4Mux_h
    port map (
            O => \N__64616\,
            I => \N__64591\
        );

    \I__15202\ : Span4Mux_h
    port map (
            O => \N__64611\,
            I => \N__64588\
        );

    \I__15201\ : Span4Mux_h
    port map (
            O => \N__64608\,
            I => \N__64583\
        );

    \I__15200\ : LocalMux
    port map (
            O => \N__64605\,
            I => \N__64583\
        );

    \I__15199\ : Span4Mux_h
    port map (
            O => \N__64602\,
            I => \N__64580\
        );

    \I__15198\ : LocalMux
    port map (
            O => \N__64599\,
            I => \N__64577\
        );

    \I__15197\ : InMux
    port map (
            O => \N__64598\,
            I => \N__64574\
        );

    \I__15196\ : InMux
    port map (
            O => \N__64597\,
            I => \N__64569\
        );

    \I__15195\ : InMux
    port map (
            O => \N__64596\,
            I => \N__64569\
        );

    \I__15194\ : InMux
    port map (
            O => \N__64595\,
            I => \N__64566\
        );

    \I__15193\ : InMux
    port map (
            O => \N__64594\,
            I => \N__64563\
        );

    \I__15192\ : Odrv4
    port map (
            O => \N__64591\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15191\ : Odrv4
    port map (
            O => \N__64588\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15190\ : Odrv4
    port map (
            O => \N__64583\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15189\ : Odrv4
    port map (
            O => \N__64580\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15188\ : Odrv12
    port map (
            O => \N__64577\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15187\ : LocalMux
    port map (
            O => \N__64574\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15186\ : LocalMux
    port map (
            O => \N__64569\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15185\ : LocalMux
    port map (
            O => \N__64566\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15184\ : LocalMux
    port map (
            O => \N__64563\,
            I => \CONTROL_programCounter11_reto_rep2\
        );

    \I__15183\ : InMux
    port map (
            O => \N__64544\,
            I => \N__64541\
        );

    \I__15182\ : LocalMux
    port map (
            O => \N__64541\,
            I => \PROM.ROMDATA.m135\
        );

    \I__15181\ : InMux
    port map (
            O => \N__64538\,
            I => \N__64535\
        );

    \I__15180\ : LocalMux
    port map (
            O => \N__64535\,
            I => \PROM.ROMDATA.m132\
        );

    \I__15179\ : InMux
    port map (
            O => \N__64532\,
            I => \N__64528\
        );

    \I__15178\ : CascadeMux
    port map (
            O => \N__64531\,
            I => \N__64525\
        );

    \I__15177\ : LocalMux
    port map (
            O => \N__64528\,
            I => \N__64521\
        );

    \I__15176\ : InMux
    port map (
            O => \N__64525\,
            I => \N__64518\
        );

    \I__15175\ : InMux
    port map (
            O => \N__64524\,
            I => \N__64515\
        );

    \I__15174\ : Span4Mux_v
    port map (
            O => \N__64521\,
            I => \N__64512\
        );

    \I__15173\ : LocalMux
    port map (
            O => \N__64518\,
            I => \N__64509\
        );

    \I__15172\ : LocalMux
    port map (
            O => \N__64515\,
            I => \N__64506\
        );

    \I__15171\ : Span4Mux_h
    port map (
            O => \N__64512\,
            I => \N__64503\
        );

    \I__15170\ : Span4Mux_v
    port map (
            O => \N__64509\,
            I => \N__64500\
        );

    \I__15169\ : Span4Mux_h
    port map (
            O => \N__64506\,
            I => \N__64497\
        );

    \I__15168\ : Span4Mux_h
    port map (
            O => \N__64503\,
            I => \N__64492\
        );

    \I__15167\ : Span4Mux_h
    port map (
            O => \N__64500\,
            I => \N__64492\
        );

    \I__15166\ : Odrv4
    port map (
            O => \N__64497\,
            I => \N_418\
        );

    \I__15165\ : Odrv4
    port map (
            O => \N__64492\,
            I => \N_418\
        );

    \I__15164\ : InMux
    port map (
            O => \N__64487\,
            I => \N__64482\
        );

    \I__15163\ : InMux
    port map (
            O => \N__64486\,
            I => \N__64479\
        );

    \I__15162\ : InMux
    port map (
            O => \N__64485\,
            I => \N__64476\
        );

    \I__15161\ : LocalMux
    port map (
            O => \N__64482\,
            I => \N__64473\
        );

    \I__15160\ : LocalMux
    port map (
            O => \N__64479\,
            I => \N__64470\
        );

    \I__15159\ : LocalMux
    port map (
            O => \N__64476\,
            I => \N__64467\
        );

    \I__15158\ : Span12Mux_s11_v
    port map (
            O => \N__64473\,
            I => \N__64462\
        );

    \I__15157\ : Span4Mux_h
    port map (
            O => \N__64470\,
            I => \N__64459\
        );

    \I__15156\ : Span4Mux_h
    port map (
            O => \N__64467\,
            I => \N__64456\
        );

    \I__15155\ : InMux
    port map (
            O => \N__64466\,
            I => \N__64451\
        );

    \I__15154\ : InMux
    port map (
            O => \N__64465\,
            I => \N__64451\
        );

    \I__15153\ : Odrv12
    port map (
            O => \N__64462\,
            I => \CONTROL_addrstack_reto_3\
        );

    \I__15152\ : Odrv4
    port map (
            O => \N__64459\,
            I => \CONTROL_addrstack_reto_3\
        );

    \I__15151\ : Odrv4
    port map (
            O => \N__64456\,
            I => \CONTROL_addrstack_reto_3\
        );

    \I__15150\ : LocalMux
    port map (
            O => \N__64451\,
            I => \CONTROL_addrstack_reto_3\
        );

    \I__15149\ : CascadeMux
    port map (
            O => \N__64442\,
            I => \N__64439\
        );

    \I__15148\ : InMux
    port map (
            O => \N__64439\,
            I => \N__64436\
        );

    \I__15147\ : LocalMux
    port map (
            O => \N__64436\,
            I => \PROM.ROMDATA.m166_e\
        );

    \I__15146\ : InMux
    port map (
            O => \N__64433\,
            I => \N__64430\
        );

    \I__15145\ : LocalMux
    port map (
            O => \N__64430\,
            I => \N__64427\
        );

    \I__15144\ : Odrv4
    port map (
            O => \N__64427\,
            I => \PROM.ROMDATA.m104_ns_1\
        );

    \I__15143\ : InMux
    port map (
            O => \N__64424\,
            I => \N__64421\
        );

    \I__15142\ : LocalMux
    port map (
            O => \N__64421\,
            I => \PROM.ROMDATA.m107\
        );

    \I__15141\ : CascadeMux
    port map (
            O => \N__64418\,
            I => \PROM.ROMDATA.m104_ns_cascade_\
        );

    \I__15140\ : InMux
    port map (
            O => \N__64415\,
            I => \N__64412\
        );

    \I__15139\ : LocalMux
    port map (
            O => \N__64412\,
            I => \N__64409\
        );

    \I__15138\ : Span4Mux_v
    port map (
            O => \N__64409\,
            I => \N__64406\
        );

    \I__15137\ : Span4Mux_h
    port map (
            O => \N__64406\,
            I => \N__64403\
        );

    \I__15136\ : Odrv4
    port map (
            O => \N__64403\,
            I => \PROM.ROMDATA.m109_am\
        );

    \I__15135\ : CascadeMux
    port map (
            O => \N__64400\,
            I => \PROM.ROMDATA.m109_bm_cascade_\
        );

    \I__15134\ : InMux
    port map (
            O => \N__64397\,
            I => \N__64393\
        );

    \I__15133\ : InMux
    port map (
            O => \N__64396\,
            I => \N__64390\
        );

    \I__15132\ : LocalMux
    port map (
            O => \N__64393\,
            I => \N__64387\
        );

    \I__15131\ : LocalMux
    port map (
            O => \N__64390\,
            I => \N__64382\
        );

    \I__15130\ : Span4Mux_v
    port map (
            O => \N__64387\,
            I => \N__64382\
        );

    \I__15129\ : Span4Mux_h
    port map (
            O => \N__64382\,
            I => \N__64379\
        );

    \I__15128\ : Odrv4
    port map (
            O => \N__64379\,
            I => \PROM.ROMDATA.m121_ns\
        );

    \I__15127\ : InMux
    port map (
            O => \N__64376\,
            I => \N__64373\
        );

    \I__15126\ : LocalMux
    port map (
            O => \N__64373\,
            I => \PROM.ROMDATA.m114\
        );

    \I__15125\ : InMux
    port map (
            O => \N__64370\,
            I => \N__64367\
        );

    \I__15124\ : LocalMux
    port map (
            O => \N__64367\,
            I => \PROM.ROMDATA.m111\
        );

    \I__15123\ : CascadeMux
    port map (
            O => \N__64364\,
            I => \PROM.ROMDATA.m120_am_cascade_\
        );

    \I__15122\ : InMux
    port map (
            O => \N__64361\,
            I => \N__64358\
        );

    \I__15121\ : LocalMux
    port map (
            O => \N__64358\,
            I => \PROM.ROMDATA.m120_bm\
        );

    \I__15120\ : InMux
    port map (
            O => \N__64355\,
            I => \N__64352\
        );

    \I__15119\ : LocalMux
    port map (
            O => \N__64352\,
            I => \PROM.ROMDATA.m121_ns_1\
        );

    \I__15118\ : CascadeMux
    port map (
            O => \N__64349\,
            I => \PROM.ROMDATA.m287_cascade_\
        );

    \I__15117\ : InMux
    port map (
            O => \N__64346\,
            I => \N__64343\
        );

    \I__15116\ : LocalMux
    port map (
            O => \N__64343\,
            I => \PROM.ROMDATA.m410_bm\
        );

    \I__15115\ : InMux
    port map (
            O => \N__64340\,
            I => \N__64337\
        );

    \I__15114\ : LocalMux
    port map (
            O => \N__64337\,
            I => \N__64334\
        );

    \I__15113\ : Span12Mux_v
    port map (
            O => \N__64334\,
            I => \N__64331\
        );

    \I__15112\ : Odrv12
    port map (
            O => \N__64331\,
            I => \PROM.ROMDATA.m66\
        );

    \I__15111\ : CascadeMux
    port map (
            O => \N__64328\,
            I => \N__64325\
        );

    \I__15110\ : InMux
    port map (
            O => \N__64325\,
            I => \N__64320\
        );

    \I__15109\ : CascadeMux
    port map (
            O => \N__64324\,
            I => \N__64317\
        );

    \I__15108\ : InMux
    port map (
            O => \N__64323\,
            I => \N__64314\
        );

    \I__15107\ : LocalMux
    port map (
            O => \N__64320\,
            I => \N__64311\
        );

    \I__15106\ : InMux
    port map (
            O => \N__64317\,
            I => \N__64308\
        );

    \I__15105\ : LocalMux
    port map (
            O => \N__64314\,
            I => \N__64305\
        );

    \I__15104\ : Odrv4
    port map (
            O => \N__64311\,
            I => \PROM.ROMDATA.m163\
        );

    \I__15103\ : LocalMux
    port map (
            O => \N__64308\,
            I => \PROM.ROMDATA.m163\
        );

    \I__15102\ : Odrv4
    port map (
            O => \N__64305\,
            I => \PROM.ROMDATA.m163\
        );

    \I__15101\ : InMux
    port map (
            O => \N__64298\,
            I => \N__64295\
        );

    \I__15100\ : LocalMux
    port map (
            O => \N__64295\,
            I => \N__64292\
        );

    \I__15099\ : Span12Mux_v
    port map (
            O => \N__64292\,
            I => \N__64289\
        );

    \I__15098\ : Odrv12
    port map (
            O => \N__64289\,
            I => \PROM.ROMDATA.m490\
        );

    \I__15097\ : CascadeMux
    port map (
            O => \N__64286\,
            I => \N__64283\
        );

    \I__15096\ : InMux
    port map (
            O => \N__64283\,
            I => \N__64280\
        );

    \I__15095\ : LocalMux
    port map (
            O => \N__64280\,
            I => \PROM.ROMDATA.m149\
        );

    \I__15094\ : InMux
    port map (
            O => \N__64277\,
            I => \N__64274\
        );

    \I__15093\ : LocalMux
    port map (
            O => \N__64274\,
            I => \PROM.ROMDATA.m118\
        );

    \I__15092\ : InMux
    port map (
            O => \N__64271\,
            I => \N__64268\
        );

    \I__15091\ : LocalMux
    port map (
            O => \N__64268\,
            I => \PROM.ROMDATA.m117\
        );

    \I__15090\ : CascadeMux
    port map (
            O => \N__64265\,
            I => \N__64262\
        );

    \I__15089\ : InMux
    port map (
            O => \N__64262\,
            I => \N__64258\
        );

    \I__15088\ : InMux
    port map (
            O => \N__64261\,
            I => \N__64255\
        );

    \I__15087\ : LocalMux
    port map (
            O => \N__64258\,
            I => \N__64251\
        );

    \I__15086\ : LocalMux
    port map (
            O => \N__64255\,
            I => \N__64247\
        );

    \I__15085\ : InMux
    port map (
            O => \N__64254\,
            I => \N__64242\
        );

    \I__15084\ : Span4Mux_v
    port map (
            O => \N__64251\,
            I => \N__64239\
        );

    \I__15083\ : InMux
    port map (
            O => \N__64250\,
            I => \N__64236\
        );

    \I__15082\ : Span4Mux_v
    port map (
            O => \N__64247\,
            I => \N__64232\
        );

    \I__15081\ : InMux
    port map (
            O => \N__64246\,
            I => \N__64229\
        );

    \I__15080\ : InMux
    port map (
            O => \N__64245\,
            I => \N__64226\
        );

    \I__15079\ : LocalMux
    port map (
            O => \N__64242\,
            I => \N__64223\
        );

    \I__15078\ : Sp12to4
    port map (
            O => \N__64239\,
            I => \N__64218\
        );

    \I__15077\ : LocalMux
    port map (
            O => \N__64236\,
            I => \N__64218\
        );

    \I__15076\ : InMux
    port map (
            O => \N__64235\,
            I => \N__64215\
        );

    \I__15075\ : Odrv4
    port map (
            O => \N__64232\,
            I => \PROM.ROMDATA.m157\
        );

    \I__15074\ : LocalMux
    port map (
            O => \N__64229\,
            I => \PROM.ROMDATA.m157\
        );

    \I__15073\ : LocalMux
    port map (
            O => \N__64226\,
            I => \PROM.ROMDATA.m157\
        );

    \I__15072\ : Odrv4
    port map (
            O => \N__64223\,
            I => \PROM.ROMDATA.m157\
        );

    \I__15071\ : Odrv12
    port map (
            O => \N__64218\,
            I => \PROM.ROMDATA.m157\
        );

    \I__15070\ : LocalMux
    port map (
            O => \N__64215\,
            I => \PROM.ROMDATA.m157\
        );

    \I__15069\ : CascadeMux
    port map (
            O => \N__64202\,
            I => \PROM.ROMDATA.m456_ns_1_cascade_\
        );

    \I__15068\ : InMux
    port map (
            O => \N__64199\,
            I => \N__64196\
        );

    \I__15067\ : LocalMux
    port map (
            O => \N__64196\,
            I => \N__64193\
        );

    \I__15066\ : Span4Mux_v
    port map (
            O => \N__64193\,
            I => \N__64190\
        );

    \I__15065\ : Odrv4
    port map (
            O => \N__64190\,
            I => \PROM.ROMDATA.m456_ns\
        );

    \I__15064\ : InMux
    port map (
            O => \N__64187\,
            I => \N__64184\
        );

    \I__15063\ : LocalMux
    port map (
            O => \N__64184\,
            I => \PROM.ROMDATA.m414_ns_1\
        );

    \I__15062\ : CascadeMux
    port map (
            O => \N__64181\,
            I => \N__64178\
        );

    \I__15061\ : InMux
    port map (
            O => \N__64178\,
            I => \N__64175\
        );

    \I__15060\ : LocalMux
    port map (
            O => \N__64175\,
            I => \N__64172\
        );

    \I__15059\ : Odrv12
    port map (
            O => \N__64172\,
            I => \PROM.ROMDATA.m413_bm\
        );

    \I__15058\ : InMux
    port map (
            O => \N__64169\,
            I => \N__64166\
        );

    \I__15057\ : LocalMux
    port map (
            O => \N__64166\,
            I => \N__64163\
        );

    \I__15056\ : Span4Mux_h
    port map (
            O => \N__64163\,
            I => \N__64160\
        );

    \I__15055\ : Odrv4
    port map (
            O => \N__64160\,
            I => \PROM.ROMDATA.m414_ns\
        );

    \I__15054\ : CascadeMux
    port map (
            O => \N__64157\,
            I => \N__64154\
        );

    \I__15053\ : InMux
    port map (
            O => \N__64154\,
            I => \N__64151\
        );

    \I__15052\ : LocalMux
    port map (
            O => \N__64151\,
            I => \N__64148\
        );

    \I__15051\ : Odrv4
    port map (
            O => \N__64148\,
            I => \PROM.ROMDATA.m304\
        );

    \I__15050\ : CascadeMux
    port map (
            O => \N__64145\,
            I => \PROM_ROMDATA_dintern_13ro_cascade_\
        );

    \I__15049\ : CascadeMux
    port map (
            O => \N__64142\,
            I => \N__64139\
        );

    \I__15048\ : InMux
    port map (
            O => \N__64139\,
            I => \N__64136\
        );

    \I__15047\ : LocalMux
    port map (
            O => \N__64136\,
            I => \N__64133\
        );

    \I__15046\ : Span4Mux_h
    port map (
            O => \N__64133\,
            I => \N__64130\
        );

    \I__15045\ : Span4Mux_v
    port map (
            O => \N__64130\,
            I => \N__64127\
        );

    \I__15044\ : Odrv4
    port map (
            O => \N__64127\,
            I => \PROM.ROMDATA.m198\
        );

    \I__15043\ : InMux
    port map (
            O => \N__64124\,
            I => \N__64120\
        );

    \I__15042\ : InMux
    port map (
            O => \N__64123\,
            I => \N__64117\
        );

    \I__15041\ : LocalMux
    port map (
            O => \N__64120\,
            I => \N__64112\
        );

    \I__15040\ : LocalMux
    port map (
            O => \N__64117\,
            I => \N__64112\
        );

    \I__15039\ : Span4Mux_v
    port map (
            O => \N__64112\,
            I => \N__64109\
        );

    \I__15038\ : Span4Mux_h
    port map (
            O => \N__64109\,
            I => \N__64102\
        );

    \I__15037\ : InMux
    port map (
            O => \N__64108\,
            I => \N__64099\
        );

    \I__15036\ : InMux
    port map (
            O => \N__64107\,
            I => \N__64092\
        );

    \I__15035\ : InMux
    port map (
            O => \N__64106\,
            I => \N__64092\
        );

    \I__15034\ : InMux
    port map (
            O => \N__64105\,
            I => \N__64092\
        );

    \I__15033\ : Odrv4
    port map (
            O => \N__64102\,
            I => \PROM.ROMDATA.m16\
        );

    \I__15032\ : LocalMux
    port map (
            O => \N__64099\,
            I => \PROM.ROMDATA.m16\
        );

    \I__15031\ : LocalMux
    port map (
            O => \N__64092\,
            I => \PROM.ROMDATA.m16\
        );

    \I__15030\ : InMux
    port map (
            O => \N__64085\,
            I => \N__64080\
        );

    \I__15029\ : InMux
    port map (
            O => \N__64084\,
            I => \N__64075\
        );

    \I__15028\ : InMux
    port map (
            O => \N__64083\,
            I => \N__64075\
        );

    \I__15027\ : LocalMux
    port map (
            O => \N__64080\,
            I => \CONTROL.N_45_0\
        );

    \I__15026\ : LocalMux
    port map (
            O => \N__64075\,
            I => \CONTROL.N_45_0\
        );

    \I__15025\ : CascadeMux
    port map (
            O => \N__64070\,
            I => \PROM_ROMDATA_dintern_15ro_cascade_\
        );

    \I__15024\ : CascadeMux
    port map (
            O => \N__64067\,
            I => \N__64064\
        );

    \I__15023\ : InMux
    port map (
            O => \N__64064\,
            I => \N__64061\
        );

    \I__15022\ : LocalMux
    port map (
            O => \N__64061\,
            I => \PROM.ROMDATA.m139\
        );

    \I__15021\ : CascadeMux
    port map (
            O => \N__64058\,
            I => \N__64054\
        );

    \I__15020\ : InMux
    port map (
            O => \N__64057\,
            I => \N__64049\
        );

    \I__15019\ : InMux
    port map (
            O => \N__64054\,
            I => \N__64049\
        );

    \I__15018\ : LocalMux
    port map (
            O => \N__64049\,
            I => \N__64046\
        );

    \I__15017\ : Span4Mux_v
    port map (
            O => \N__64046\,
            I => \N__64043\
        );

    \I__15016\ : Span4Mux_h
    port map (
            O => \N__64043\,
            I => \N__64040\
        );

    \I__15015\ : Span4Mux_h
    port map (
            O => \N__64040\,
            I => \N__64037\
        );

    \I__15014\ : Span4Mux_v
    port map (
            O => \N__64037\,
            I => \N__64034\
        );

    \I__15013\ : Odrv4
    port map (
            O => \N__64034\,
            I => \PROM.ROMDATA.N_564_mux\
        );

    \I__15012\ : InMux
    port map (
            O => \N__64031\,
            I => \N__64028\
        );

    \I__15011\ : LocalMux
    port map (
            O => \N__64028\,
            I => \N__64025\
        );

    \I__15010\ : Odrv4
    port map (
            O => \N__64025\,
            I => \PROM.ROMDATA.m298_bm\
        );

    \I__15009\ : InMux
    port map (
            O => \N__64022\,
            I => \N__64019\
        );

    \I__15008\ : LocalMux
    port map (
            O => \N__64019\,
            I => \N__64014\
        );

    \I__15007\ : CascadeMux
    port map (
            O => \N__64018\,
            I => \N__64011\
        );

    \I__15006\ : InMux
    port map (
            O => \N__64017\,
            I => \N__64008\
        );

    \I__15005\ : Span4Mux_h
    port map (
            O => \N__64014\,
            I => \N__64004\
        );

    \I__15004\ : InMux
    port map (
            O => \N__64011\,
            I => \N__64001\
        );

    \I__15003\ : LocalMux
    port map (
            O => \N__64008\,
            I => \N__63998\
        );

    \I__15002\ : InMux
    port map (
            O => \N__64007\,
            I => \N__63995\
        );

    \I__15001\ : Span4Mux_v
    port map (
            O => \N__64004\,
            I => \N__63992\
        );

    \I__15000\ : LocalMux
    port map (
            O => \N__64001\,
            I => \N__63987\
        );

    \I__14999\ : Span4Mux_v
    port map (
            O => \N__63998\,
            I => \N__63987\
        );

    \I__14998\ : LocalMux
    port map (
            O => \N__63995\,
            I => \N__63984\
        );

    \I__14997\ : Sp12to4
    port map (
            O => \N__63992\,
            I => \N__63981\
        );

    \I__14996\ : Span4Mux_v
    port map (
            O => \N__63987\,
            I => \N__63978\
        );

    \I__14995\ : Span4Mux_h
    port map (
            O => \N__63984\,
            I => \N__63975\
        );

    \I__14994\ : Odrv12
    port map (
            O => \N__63981\,
            I => \PROM.ROMDATA.N_72_i\
        );

    \I__14993\ : Odrv4
    port map (
            O => \N__63978\,
            I => \PROM.ROMDATA.N_72_i\
        );

    \I__14992\ : Odrv4
    port map (
            O => \N__63975\,
            I => \PROM.ROMDATA.N_72_i\
        );

    \I__14991\ : CascadeMux
    port map (
            O => \N__63968\,
            I => \N__63964\
        );

    \I__14990\ : InMux
    port map (
            O => \N__63967\,
            I => \N__63959\
        );

    \I__14989\ : InMux
    port map (
            O => \N__63964\,
            I => \N__63959\
        );

    \I__14988\ : LocalMux
    port map (
            O => \N__63959\,
            I => \N__63956\
        );

    \I__14987\ : Span12Mux_v
    port map (
            O => \N__63956\,
            I => \N__63953\
        );

    \I__14986\ : Odrv12
    port map (
            O => \N__63953\,
            I => \PROM.ROMDATA.N_565_mux\
        );

    \I__14985\ : InMux
    port map (
            O => \N__63950\,
            I => \N__63947\
        );

    \I__14984\ : LocalMux
    port map (
            O => \N__63947\,
            I => \N__63944\
        );

    \I__14983\ : Span4Mux_h
    port map (
            O => \N__63944\,
            I => \N__63941\
        );

    \I__14982\ : Odrv4
    port map (
            O => \N__63941\,
            I => \PROM.ROMDATA.m498_bm\
        );

    \I__14981\ : CascadeMux
    port map (
            O => \N__63938\,
            I => \PROM.ROMDATA.m498_am_cascade_\
        );

    \I__14980\ : CascadeMux
    port map (
            O => \N__63935\,
            I => \N__63932\
        );

    \I__14979\ : InMux
    port map (
            O => \N__63932\,
            I => \N__63929\
        );

    \I__14978\ : LocalMux
    port map (
            O => \N__63929\,
            I => \PROM.ROMDATA.m498_ns\
        );

    \I__14977\ : InMux
    port map (
            O => \N__63926\,
            I => \N__63923\
        );

    \I__14976\ : LocalMux
    port map (
            O => \N__63923\,
            I => \N__63920\
        );

    \I__14975\ : Span12Mux_v
    port map (
            O => \N__63920\,
            I => \N__63917\
        );

    \I__14974\ : Odrv12
    port map (
            O => \N__63917\,
            I => \PROM.ROMDATA.m317_am\
        );

    \I__14973\ : CascadeMux
    port map (
            O => \N__63914\,
            I => \PROM.ROMDATA.m317_bm_cascade_\
        );

    \I__14972\ : InMux
    port map (
            O => \N__63911\,
            I => \N__63908\
        );

    \I__14971\ : LocalMux
    port map (
            O => \N__63908\,
            I => \N__63905\
        );

    \I__14970\ : Span4Mux_v
    port map (
            O => \N__63905\,
            I => \N__63902\
        );

    \I__14969\ : Odrv4
    port map (
            O => \N__63902\,
            I => \PROM.ROMDATA.m312_ns\
        );

    \I__14968\ : CascadeMux
    port map (
            O => \N__63899\,
            I => \PROM.ROMDATA.m317_ns_cascade_\
        );

    \I__14967\ : CascadeMux
    port map (
            O => \N__63896\,
            I => \PROM.ROMDATA.m325_ns_1_cascade_\
        );

    \I__14966\ : InMux
    port map (
            O => \N__63893\,
            I => \N__63890\
        );

    \I__14965\ : LocalMux
    port map (
            O => \N__63890\,
            I => \N__63887\
        );

    \I__14964\ : Odrv4
    port map (
            O => \N__63887\,
            I => \PROM.ROMDATA.m320_ns\
        );

    \I__14963\ : CascadeMux
    port map (
            O => \N__63884\,
            I => \N__63881\
        );

    \I__14962\ : InMux
    port map (
            O => \N__63881\,
            I => \N__63878\
        );

    \I__14961\ : LocalMux
    port map (
            O => \N__63878\,
            I => \N__63875\
        );

    \I__14960\ : Odrv4
    port map (
            O => \N__63875\,
            I => \PROM.ROMDATA.m325_ns\
        );

    \I__14959\ : CascadeMux
    port map (
            O => \N__63872\,
            I => \PROM_ROMDATA_dintern_14ro_cascade_\
        );

    \I__14958\ : InMux
    port map (
            O => \N__63869\,
            I => \N__63866\
        );

    \I__14957\ : LocalMux
    port map (
            O => \N__63866\,
            I => \PROM.ROMDATA.m494_ns\
        );

    \I__14956\ : InMux
    port map (
            O => \N__63863\,
            I => \ALU.addsub_cry_12\
        );

    \I__14955\ : InMux
    port map (
            O => \N__63860\,
            I => \N__63857\
        );

    \I__14954\ : LocalMux
    port map (
            O => \N__63857\,
            I => \ALU.c_RNIDDGOIZ0Z_14\
        );

    \I__14953\ : CascadeMux
    port map (
            O => \N__63854\,
            I => \N__63849\
        );

    \I__14952\ : CascadeMux
    port map (
            O => \N__63853\,
            I => \N__63844\
        );

    \I__14951\ : InMux
    port map (
            O => \N__63852\,
            I => \N__63839\
        );

    \I__14950\ : InMux
    port map (
            O => \N__63849\,
            I => \N__63836\
        );

    \I__14949\ : CascadeMux
    port map (
            O => \N__63848\,
            I => \N__63832\
        );

    \I__14948\ : InMux
    port map (
            O => \N__63847\,
            I => \N__63829\
        );

    \I__14947\ : InMux
    port map (
            O => \N__63844\,
            I => \N__63826\
        );

    \I__14946\ : InMux
    port map (
            O => \N__63843\,
            I => \N__63823\
        );

    \I__14945\ : CascadeMux
    port map (
            O => \N__63842\,
            I => \N__63820\
        );

    \I__14944\ : LocalMux
    port map (
            O => \N__63839\,
            I => \N__63816\
        );

    \I__14943\ : LocalMux
    port map (
            O => \N__63836\,
            I => \N__63813\
        );

    \I__14942\ : InMux
    port map (
            O => \N__63835\,
            I => \N__63810\
        );

    \I__14941\ : InMux
    port map (
            O => \N__63832\,
            I => \N__63806\
        );

    \I__14940\ : LocalMux
    port map (
            O => \N__63829\,
            I => \N__63803\
        );

    \I__14939\ : LocalMux
    port map (
            O => \N__63826\,
            I => \N__63797\
        );

    \I__14938\ : LocalMux
    port map (
            O => \N__63823\,
            I => \N__63797\
        );

    \I__14937\ : InMux
    port map (
            O => \N__63820\,
            I => \N__63794\
        );

    \I__14936\ : CascadeMux
    port map (
            O => \N__63819\,
            I => \N__63791\
        );

    \I__14935\ : Span4Mux_v
    port map (
            O => \N__63816\,
            I => \N__63788\
        );

    \I__14934\ : Span4Mux_v
    port map (
            O => \N__63813\,
            I => \N__63783\
        );

    \I__14933\ : LocalMux
    port map (
            O => \N__63810\,
            I => \N__63783\
        );

    \I__14932\ : InMux
    port map (
            O => \N__63809\,
            I => \N__63780\
        );

    \I__14931\ : LocalMux
    port map (
            O => \N__63806\,
            I => \N__63775\
        );

    \I__14930\ : Span4Mux_v
    port map (
            O => \N__63803\,
            I => \N__63771\
        );

    \I__14929\ : InMux
    port map (
            O => \N__63802\,
            I => \N__63768\
        );

    \I__14928\ : Span4Mux_v
    port map (
            O => \N__63797\,
            I => \N__63763\
        );

    \I__14927\ : LocalMux
    port map (
            O => \N__63794\,
            I => \N__63763\
        );

    \I__14926\ : InMux
    port map (
            O => \N__63791\,
            I => \N__63760\
        );

    \I__14925\ : Span4Mux_h
    port map (
            O => \N__63788\,
            I => \N__63753\
        );

    \I__14924\ : Span4Mux_h
    port map (
            O => \N__63783\,
            I => \N__63753\
        );

    \I__14923\ : LocalMux
    port map (
            O => \N__63780\,
            I => \N__63753\
        );

    \I__14922\ : InMux
    port map (
            O => \N__63779\,
            I => \N__63748\
        );

    \I__14921\ : InMux
    port map (
            O => \N__63778\,
            I => \N__63748\
        );

    \I__14920\ : Span4Mux_v
    port map (
            O => \N__63775\,
            I => \N__63745\
        );

    \I__14919\ : InMux
    port map (
            O => \N__63774\,
            I => \N__63742\
        );

    \I__14918\ : Span4Mux_v
    port map (
            O => \N__63771\,
            I => \N__63739\
        );

    \I__14917\ : LocalMux
    port map (
            O => \N__63768\,
            I => \N__63734\
        );

    \I__14916\ : Span4Mux_v
    port map (
            O => \N__63763\,
            I => \N__63734\
        );

    \I__14915\ : LocalMux
    port map (
            O => \N__63760\,
            I => \N__63731\
        );

    \I__14914\ : Span4Mux_v
    port map (
            O => \N__63753\,
            I => \N__63728\
        );

    \I__14913\ : LocalMux
    port map (
            O => \N__63748\,
            I => \N__63721\
        );

    \I__14912\ : Span4Mux_v
    port map (
            O => \N__63745\,
            I => \N__63721\
        );

    \I__14911\ : LocalMux
    port map (
            O => \N__63742\,
            I => \N__63721\
        );

    \I__14910\ : Span4Mux_h
    port map (
            O => \N__63739\,
            I => \N__63716\
        );

    \I__14909\ : Span4Mux_v
    port map (
            O => \N__63734\,
            I => \N__63716\
        );

    \I__14908\ : Span4Mux_v
    port map (
            O => \N__63731\,
            I => \N__63711\
        );

    \I__14907\ : Span4Mux_v
    port map (
            O => \N__63728\,
            I => \N__63711\
        );

    \I__14906\ : Span4Mux_v
    port map (
            O => \N__63721\,
            I => \N__63706\
        );

    \I__14905\ : Span4Mux_h
    port map (
            O => \N__63716\,
            I => \N__63706\
        );

    \I__14904\ : Odrv4
    port map (
            O => \N__63711\,
            I => \aluOut_14\
        );

    \I__14903\ : Odrv4
    port map (
            O => \N__63706\,
            I => \aluOut_14\
        );

    \I__14902\ : InMux
    port map (
            O => \N__63701\,
            I => \N__63694\
        );

    \I__14901\ : InMux
    port map (
            O => \N__63700\,
            I => \N__63694\
        );

    \I__14900\ : InMux
    port map (
            O => \N__63699\,
            I => \N__63691\
        );

    \I__14899\ : LocalMux
    port map (
            O => \N__63694\,
            I => \N__63688\
        );

    \I__14898\ : LocalMux
    port map (
            O => \N__63691\,
            I => \ALU.addsub_14\
        );

    \I__14897\ : Odrv12
    port map (
            O => \N__63688\,
            I => \ALU.addsub_14\
        );

    \I__14896\ : InMux
    port map (
            O => \N__63683\,
            I => \ALU.addsub_cry_13\
        );

    \I__14895\ : InMux
    port map (
            O => \N__63680\,
            I => \N__63677\
        );

    \I__14894\ : LocalMux
    port map (
            O => \N__63677\,
            I => \ALU.c_RNI0NMSHZ0Z_15\
        );

    \I__14893\ : InMux
    port map (
            O => \N__63674\,
            I => \N__63671\
        );

    \I__14892\ : LocalMux
    port map (
            O => \N__63671\,
            I => \N__63665\
        );

    \I__14891\ : CascadeMux
    port map (
            O => \N__63670\,
            I => \N__63662\
        );

    \I__14890\ : InMux
    port map (
            O => \N__63669\,
            I => \N__63659\
        );

    \I__14889\ : InMux
    port map (
            O => \N__63668\,
            I => \N__63655\
        );

    \I__14888\ : Span4Mux_h
    port map (
            O => \N__63665\,
            I => \N__63652\
        );

    \I__14887\ : InMux
    port map (
            O => \N__63662\,
            I => \N__63649\
        );

    \I__14886\ : LocalMux
    port map (
            O => \N__63659\,
            I => \N__63646\
        );

    \I__14885\ : InMux
    port map (
            O => \N__63658\,
            I => \N__63641\
        );

    \I__14884\ : LocalMux
    port map (
            O => \N__63655\,
            I => \N__63635\
        );

    \I__14883\ : Span4Mux_h
    port map (
            O => \N__63652\,
            I => \N__63628\
        );

    \I__14882\ : LocalMux
    port map (
            O => \N__63649\,
            I => \N__63628\
        );

    \I__14881\ : Span4Mux_v
    port map (
            O => \N__63646\,
            I => \N__63628\
        );

    \I__14880\ : InMux
    port map (
            O => \N__63645\,
            I => \N__63625\
        );

    \I__14879\ : InMux
    port map (
            O => \N__63644\,
            I => \N__63622\
        );

    \I__14878\ : LocalMux
    port map (
            O => \N__63641\,
            I => \N__63619\
        );

    \I__14877\ : InMux
    port map (
            O => \N__63640\,
            I => \N__63616\
        );

    \I__14876\ : InMux
    port map (
            O => \N__63639\,
            I => \N__63607\
        );

    \I__14875\ : InMux
    port map (
            O => \N__63638\,
            I => \N__63607\
        );

    \I__14874\ : Span4Mux_v
    port map (
            O => \N__63635\,
            I => \N__63598\
        );

    \I__14873\ : Span4Mux_h
    port map (
            O => \N__63628\,
            I => \N__63598\
        );

    \I__14872\ : LocalMux
    port map (
            O => \N__63625\,
            I => \N__63598\
        );

    \I__14871\ : LocalMux
    port map (
            O => \N__63622\,
            I => \N__63598\
        );

    \I__14870\ : Span4Mux_h
    port map (
            O => \N__63619\,
            I => \N__63595\
        );

    \I__14869\ : LocalMux
    port map (
            O => \N__63616\,
            I => \N__63589\
        );

    \I__14868\ : InMux
    port map (
            O => \N__63615\,
            I => \N__63586\
        );

    \I__14867\ : CascadeMux
    port map (
            O => \N__63614\,
            I => \N__63583\
        );

    \I__14866\ : CascadeMux
    port map (
            O => \N__63613\,
            I => \N__63579\
        );

    \I__14865\ : CascadeMux
    port map (
            O => \N__63612\,
            I => \N__63576\
        );

    \I__14864\ : LocalMux
    port map (
            O => \N__63607\,
            I => \N__63571\
        );

    \I__14863\ : Span4Mux_h
    port map (
            O => \N__63598\,
            I => \N__63571\
        );

    \I__14862\ : Span4Mux_h
    port map (
            O => \N__63595\,
            I => \N__63568\
        );

    \I__14861\ : InMux
    port map (
            O => \N__63594\,
            I => \N__63561\
        );

    \I__14860\ : InMux
    port map (
            O => \N__63593\,
            I => \N__63561\
        );

    \I__14859\ : InMux
    port map (
            O => \N__63592\,
            I => \N__63561\
        );

    \I__14858\ : Span12Mux_s10_h
    port map (
            O => \N__63589\,
            I => \N__63558\
        );

    \I__14857\ : LocalMux
    port map (
            O => \N__63586\,
            I => \N__63555\
        );

    \I__14856\ : InMux
    port map (
            O => \N__63583\,
            I => \N__63548\
        );

    \I__14855\ : InMux
    port map (
            O => \N__63582\,
            I => \N__63548\
        );

    \I__14854\ : InMux
    port map (
            O => \N__63579\,
            I => \N__63548\
        );

    \I__14853\ : InMux
    port map (
            O => \N__63576\,
            I => \N__63545\
        );

    \I__14852\ : Span4Mux_v
    port map (
            O => \N__63571\,
            I => \N__63542\
        );

    \I__14851\ : Span4Mux_v
    port map (
            O => \N__63568\,
            I => \N__63537\
        );

    \I__14850\ : LocalMux
    port map (
            O => \N__63561\,
            I => \N__63537\
        );

    \I__14849\ : Odrv12
    port map (
            O => \N__63558\,
            I => \aluOut_15\
        );

    \I__14848\ : Odrv12
    port map (
            O => \N__63555\,
            I => \aluOut_15\
        );

    \I__14847\ : LocalMux
    port map (
            O => \N__63548\,
            I => \aluOut_15\
        );

    \I__14846\ : LocalMux
    port map (
            O => \N__63545\,
            I => \aluOut_15\
        );

    \I__14845\ : Odrv4
    port map (
            O => \N__63542\,
            I => \aluOut_15\
        );

    \I__14844\ : Odrv4
    port map (
            O => \N__63537\,
            I => \aluOut_15\
        );

    \I__14843\ : InMux
    port map (
            O => \N__63524\,
            I => \N__63520\
        );

    \I__14842\ : InMux
    port map (
            O => \N__63523\,
            I => \N__63517\
        );

    \I__14841\ : LocalMux
    port map (
            O => \N__63520\,
            I => \N__63513\
        );

    \I__14840\ : LocalMux
    port map (
            O => \N__63517\,
            I => \N__63509\
        );

    \I__14839\ : InMux
    port map (
            O => \N__63516\,
            I => \N__63506\
        );

    \I__14838\ : Span4Mux_h
    port map (
            O => \N__63513\,
            I => \N__63503\
        );

    \I__14837\ : InMux
    port map (
            O => \N__63512\,
            I => \N__63500\
        );

    \I__14836\ : Span4Mux_h
    port map (
            O => \N__63509\,
            I => \N__63497\
        );

    \I__14835\ : LocalMux
    port map (
            O => \N__63506\,
            I => \ALU.addsub_15\
        );

    \I__14834\ : Odrv4
    port map (
            O => \N__63503\,
            I => \ALU.addsub_15\
        );

    \I__14833\ : LocalMux
    port map (
            O => \N__63500\,
            I => \ALU.addsub_15\
        );

    \I__14832\ : Odrv4
    port map (
            O => \N__63497\,
            I => \ALU.addsub_15\
        );

    \I__14831\ : InMux
    port map (
            O => \N__63488\,
            I => \bfn_23_16_0_\
        );

    \I__14830\ : CascadeMux
    port map (
            O => \N__63485\,
            I => \N__63482\
        );

    \I__14829\ : InMux
    port map (
            O => \N__63482\,
            I => \N__63478\
        );

    \I__14828\ : CascadeMux
    port map (
            O => \N__63481\,
            I => \N__63475\
        );

    \I__14827\ : LocalMux
    port map (
            O => \N__63478\,
            I => \N__63472\
        );

    \I__14826\ : InMux
    port map (
            O => \N__63475\,
            I => \N__63469\
        );

    \I__14825\ : Span4Mux_h
    port map (
            O => \N__63472\,
            I => \N__63464\
        );

    \I__14824\ : LocalMux
    port map (
            O => \N__63469\,
            I => \N__63464\
        );

    \I__14823\ : Span4Mux_h
    port map (
            O => \N__63464\,
            I => \N__63456\
        );

    \I__14822\ : InMux
    port map (
            O => \N__63463\,
            I => \N__63453\
        );

    \I__14821\ : InMux
    port map (
            O => \N__63462\,
            I => \N__63448\
        );

    \I__14820\ : InMux
    port map (
            O => \N__63461\,
            I => \N__63448\
        );

    \I__14819\ : InMux
    port map (
            O => \N__63460\,
            I => \N__63443\
        );

    \I__14818\ : InMux
    port map (
            O => \N__63459\,
            I => \N__63443\
        );

    \I__14817\ : Span4Mux_v
    port map (
            O => \N__63456\,
            I => \N__63435\
        );

    \I__14816\ : LocalMux
    port map (
            O => \N__63453\,
            I => \N__63435\
        );

    \I__14815\ : LocalMux
    port map (
            O => \N__63448\,
            I => \N__63435\
        );

    \I__14814\ : LocalMux
    port map (
            O => \N__63443\,
            I => \N__63432\
        );

    \I__14813\ : InMux
    port map (
            O => \N__63442\,
            I => \N__63429\
        );

    \I__14812\ : Span4Mux_h
    port map (
            O => \N__63435\,
            I => \N__63426\
        );

    \I__14811\ : Span4Mux_v
    port map (
            O => \N__63432\,
            I => \N__63423\
        );

    \I__14810\ : LocalMux
    port map (
            O => \N__63429\,
            I => \N__63418\
        );

    \I__14809\ : Span4Mux_h
    port map (
            O => \N__63426\,
            I => \N__63418\
        );

    \I__14808\ : Span4Mux_h
    port map (
            O => \N__63423\,
            I => \N__63415\
        );

    \I__14807\ : Span4Mux_v
    port map (
            O => \N__63418\,
            I => \N__63411\
        );

    \I__14806\ : Span4Mux_v
    port map (
            O => \N__63415\,
            I => \N__63408\
        );

    \I__14805\ : InMux
    port map (
            O => \N__63414\,
            I => \N__63405\
        );

    \I__14804\ : Span4Mux_v
    port map (
            O => \N__63411\,
            I => \N__63402\
        );

    \I__14803\ : Span4Mux_v
    port map (
            O => \N__63408\,
            I => \N__63399\
        );

    \I__14802\ : LocalMux
    port map (
            O => \N__63405\,
            I => \aluStatus_1\
        );

    \I__14801\ : Odrv4
    port map (
            O => \N__63402\,
            I => \aluStatus_1\
        );

    \I__14800\ : Odrv4
    port map (
            O => \N__63399\,
            I => \aluStatus_1\
        );

    \I__14799\ : InMux
    port map (
            O => \N__63392\,
            I => \ALU.addsub_cry_15\
        );

    \I__14798\ : InMux
    port map (
            O => \N__63389\,
            I => \N__63386\
        );

    \I__14797\ : LocalMux
    port map (
            O => \N__63386\,
            I => \N__63383\
        );

    \I__14796\ : Odrv12
    port map (
            O => \N__63383\,
            I => \ALU.N_545\
        );

    \I__14795\ : IoInMux
    port map (
            O => \N__63380\,
            I => \N__63377\
        );

    \I__14794\ : LocalMux
    port map (
            O => \N__63377\,
            I => \N__63374\
        );

    \I__14793\ : Span4Mux_s1_h
    port map (
            O => \N__63374\,
            I => \N__63371\
        );

    \I__14792\ : Span4Mux_v
    port map (
            O => \N__63371\,
            I => \N__63367\
        );

    \I__14791\ : IoInMux
    port map (
            O => \N__63370\,
            I => \N__63364\
        );

    \I__14790\ : Span4Mux_v
    port map (
            O => \N__63367\,
            I => \N__63361\
        );

    \I__14789\ : LocalMux
    port map (
            O => \N__63364\,
            I => \N__63357\
        );

    \I__14788\ : Span4Mux_h
    port map (
            O => \N__63361\,
            I => \N__63354\
        );

    \I__14787\ : InMux
    port map (
            O => \N__63360\,
            I => \N__63351\
        );

    \I__14786\ : IoSpan4Mux
    port map (
            O => \N__63357\,
            I => \N__63348\
        );

    \I__14785\ : Span4Mux_h
    port map (
            O => \N__63354\,
            I => \N__63343\
        );

    \I__14784\ : LocalMux
    port map (
            O => \N__63351\,
            I => \N__63343\
        );

    \I__14783\ : Span4Mux_s3_h
    port map (
            O => \N__63348\,
            I => \N__63340\
        );

    \I__14782\ : Span4Mux_v
    port map (
            O => \N__63343\,
            I => \N__63337\
        );

    \I__14781\ : Sp12to4
    port map (
            O => \N__63340\,
            I => \N__63334\
        );

    \I__14780\ : Sp12to4
    port map (
            O => \N__63337\,
            I => \N__63331\
        );

    \I__14779\ : Span12Mux_v
    port map (
            O => \N__63334\,
            I => \N__63328\
        );

    \I__14778\ : Span12Mux_h
    port map (
            O => \N__63331\,
            I => \N__63325\
        );

    \I__14777\ : Odrv12
    port map (
            O => \N__63328\,
            I => bus_6
        );

    \I__14776\ : Odrv12
    port map (
            O => \N__63325\,
            I => bus_6
        );

    \I__14775\ : InMux
    port map (
            O => \N__63320\,
            I => \N__63314\
        );

    \I__14774\ : InMux
    port map (
            O => \N__63319\,
            I => \N__63314\
        );

    \I__14773\ : LocalMux
    port map (
            O => \N__63314\,
            I => \N__63311\
        );

    \I__14772\ : Span4Mux_h
    port map (
            O => \N__63311\,
            I => \N__63308\
        );

    \I__14771\ : Span4Mux_h
    port map (
            O => \N__63308\,
            I => \N__63305\
        );

    \I__14770\ : Odrv4
    port map (
            O => \N__63305\,
            I => \ALU.c_RNIPBAG72Z0Z_14\
        );

    \I__14769\ : CascadeMux
    port map (
            O => \N__63302\,
            I => \N__63294\
        );

    \I__14768\ : InMux
    port map (
            O => \N__63301\,
            I => \N__63280\
        );

    \I__14767\ : InMux
    port map (
            O => \N__63300\,
            I => \N__63280\
        );

    \I__14766\ : InMux
    port map (
            O => \N__63299\,
            I => \N__63280\
        );

    \I__14765\ : InMux
    port map (
            O => \N__63298\,
            I => \N__63280\
        );

    \I__14764\ : CascadeMux
    port map (
            O => \N__63297\,
            I => \N__63277\
        );

    \I__14763\ : InMux
    port map (
            O => \N__63294\,
            I => \N__63270\
        );

    \I__14762\ : CascadeMux
    port map (
            O => \N__63293\,
            I => \N__63266\
        );

    \I__14761\ : CascadeMux
    port map (
            O => \N__63292\,
            I => \N__63262\
        );

    \I__14760\ : InMux
    port map (
            O => \N__63291\,
            I => \N__63257\
        );

    \I__14759\ : CascadeMux
    port map (
            O => \N__63290\,
            I => \N__63250\
        );

    \I__14758\ : InMux
    port map (
            O => \N__63289\,
            I => \N__63243\
        );

    \I__14757\ : LocalMux
    port map (
            O => \N__63280\,
            I => \N__63235\
        );

    \I__14756\ : InMux
    port map (
            O => \N__63277\,
            I => \N__63232\
        );

    \I__14755\ : InMux
    port map (
            O => \N__63276\,
            I => \N__63229\
        );

    \I__14754\ : CascadeMux
    port map (
            O => \N__63275\,
            I => \N__63226\
        );

    \I__14753\ : CascadeMux
    port map (
            O => \N__63274\,
            I => \N__63222\
        );

    \I__14752\ : CascadeMux
    port map (
            O => \N__63273\,
            I => \N__63219\
        );

    \I__14751\ : LocalMux
    port map (
            O => \N__63270\,
            I => \N__63214\
        );

    \I__14750\ : InMux
    port map (
            O => \N__63269\,
            I => \N__63209\
        );

    \I__14749\ : InMux
    port map (
            O => \N__63266\,
            I => \N__63209\
        );

    \I__14748\ : InMux
    port map (
            O => \N__63265\,
            I => \N__63204\
        );

    \I__14747\ : InMux
    port map (
            O => \N__63262\,
            I => \N__63204\
        );

    \I__14746\ : InMux
    port map (
            O => \N__63261\,
            I => \N__63199\
        );

    \I__14745\ : InMux
    port map (
            O => \N__63260\,
            I => \N__63199\
        );

    \I__14744\ : LocalMux
    port map (
            O => \N__63257\,
            I => \N__63196\
        );

    \I__14743\ : InMux
    port map (
            O => \N__63256\,
            I => \N__63193\
        );

    \I__14742\ : InMux
    port map (
            O => \N__63255\,
            I => \N__63188\
        );

    \I__14741\ : InMux
    port map (
            O => \N__63254\,
            I => \N__63188\
        );

    \I__14740\ : InMux
    port map (
            O => \N__63253\,
            I => \N__63185\
        );

    \I__14739\ : InMux
    port map (
            O => \N__63250\,
            I => \N__63178\
        );

    \I__14738\ : InMux
    port map (
            O => \N__63249\,
            I => \N__63178\
        );

    \I__14737\ : InMux
    port map (
            O => \N__63248\,
            I => \N__63178\
        );

    \I__14736\ : InMux
    port map (
            O => \N__63247\,
            I => \N__63173\
        );

    \I__14735\ : InMux
    port map (
            O => \N__63246\,
            I => \N__63173\
        );

    \I__14734\ : LocalMux
    port map (
            O => \N__63243\,
            I => \N__63170\
        );

    \I__14733\ : InMux
    port map (
            O => \N__63242\,
            I => \N__63163\
        );

    \I__14732\ : InMux
    port map (
            O => \N__63241\,
            I => \N__63163\
        );

    \I__14731\ : InMux
    port map (
            O => \N__63240\,
            I => \N__63163\
        );

    \I__14730\ : InMux
    port map (
            O => \N__63239\,
            I => \N__63158\
        );

    \I__14729\ : InMux
    port map (
            O => \N__63238\,
            I => \N__63158\
        );

    \I__14728\ : Span4Mux_v
    port map (
            O => \N__63235\,
            I => \N__63151\
        );

    \I__14727\ : LocalMux
    port map (
            O => \N__63232\,
            I => \N__63151\
        );

    \I__14726\ : LocalMux
    port map (
            O => \N__63229\,
            I => \N__63151\
        );

    \I__14725\ : InMux
    port map (
            O => \N__63226\,
            I => \N__63147\
        );

    \I__14724\ : InMux
    port map (
            O => \N__63225\,
            I => \N__63142\
        );

    \I__14723\ : InMux
    port map (
            O => \N__63222\,
            I => \N__63142\
        );

    \I__14722\ : InMux
    port map (
            O => \N__63219\,
            I => \N__63135\
        );

    \I__14721\ : InMux
    port map (
            O => \N__63218\,
            I => \N__63135\
        );

    \I__14720\ : InMux
    port map (
            O => \N__63217\,
            I => \N__63135\
        );

    \I__14719\ : Span4Mux_v
    port map (
            O => \N__63214\,
            I => \N__63132\
        );

    \I__14718\ : LocalMux
    port map (
            O => \N__63209\,
            I => \N__63125\
        );

    \I__14717\ : LocalMux
    port map (
            O => \N__63204\,
            I => \N__63125\
        );

    \I__14716\ : LocalMux
    port map (
            O => \N__63199\,
            I => \N__63125\
        );

    \I__14715\ : Span4Mux_v
    port map (
            O => \N__63196\,
            I => \N__63122\
        );

    \I__14714\ : LocalMux
    port map (
            O => \N__63193\,
            I => \N__63117\
        );

    \I__14713\ : LocalMux
    port map (
            O => \N__63188\,
            I => \N__63117\
        );

    \I__14712\ : LocalMux
    port map (
            O => \N__63185\,
            I => \N__63109\
        );

    \I__14711\ : LocalMux
    port map (
            O => \N__63178\,
            I => \N__63106\
        );

    \I__14710\ : LocalMux
    port map (
            O => \N__63173\,
            I => \N__63103\
        );

    \I__14709\ : Span4Mux_v
    port map (
            O => \N__63170\,
            I => \N__63100\
        );

    \I__14708\ : LocalMux
    port map (
            O => \N__63163\,
            I => \N__63093\
        );

    \I__14707\ : LocalMux
    port map (
            O => \N__63158\,
            I => \N__63093\
        );

    \I__14706\ : Span4Mux_v
    port map (
            O => \N__63151\,
            I => \N__63093\
        );

    \I__14705\ : InMux
    port map (
            O => \N__63150\,
            I => \N__63090\
        );

    \I__14704\ : LocalMux
    port map (
            O => \N__63147\,
            I => \N__63087\
        );

    \I__14703\ : LocalMux
    port map (
            O => \N__63142\,
            I => \N__63082\
        );

    \I__14702\ : LocalMux
    port map (
            O => \N__63135\,
            I => \N__63082\
        );

    \I__14701\ : Span4Mux_v
    port map (
            O => \N__63132\,
            I => \N__63077\
        );

    \I__14700\ : Span4Mux_v
    port map (
            O => \N__63125\,
            I => \N__63077\
        );

    \I__14699\ : Span4Mux_v
    port map (
            O => \N__63122\,
            I => \N__63070\
        );

    \I__14698\ : Span4Mux_v
    port map (
            O => \N__63117\,
            I => \N__63070\
        );

    \I__14697\ : InMux
    port map (
            O => \N__63116\,
            I => \N__63067\
        );

    \I__14696\ : InMux
    port map (
            O => \N__63115\,
            I => \N__63062\
        );

    \I__14695\ : InMux
    port map (
            O => \N__63114\,
            I => \N__63062\
        );

    \I__14694\ : InMux
    port map (
            O => \N__63113\,
            I => \N__63059\
        );

    \I__14693\ : InMux
    port map (
            O => \N__63112\,
            I => \N__63056\
        );

    \I__14692\ : Span4Mux_v
    port map (
            O => \N__63109\,
            I => \N__63053\
        );

    \I__14691\ : Span4Mux_v
    port map (
            O => \N__63106\,
            I => \N__63050\
        );

    \I__14690\ : Span4Mux_v
    port map (
            O => \N__63103\,
            I => \N__63047\
        );

    \I__14689\ : Span4Mux_h
    port map (
            O => \N__63100\,
            I => \N__63044\
        );

    \I__14688\ : Span4Mux_v
    port map (
            O => \N__63093\,
            I => \N__63041\
        );

    \I__14687\ : LocalMux
    port map (
            O => \N__63090\,
            I => \N__63036\
        );

    \I__14686\ : Span4Mux_v
    port map (
            O => \N__63087\,
            I => \N__63036\
        );

    \I__14685\ : Span4Mux_h
    port map (
            O => \N__63082\,
            I => \N__63031\
        );

    \I__14684\ : Span4Mux_h
    port map (
            O => \N__63077\,
            I => \N__63031\
        );

    \I__14683\ : CascadeMux
    port map (
            O => \N__63076\,
            I => \N__63027\
        );

    \I__14682\ : CascadeMux
    port map (
            O => \N__63075\,
            I => \N__63023\
        );

    \I__14681\ : Sp12to4
    port map (
            O => \N__63070\,
            I => \N__63009\
        );

    \I__14680\ : LocalMux
    port map (
            O => \N__63067\,
            I => \N__63009\
        );

    \I__14679\ : LocalMux
    port map (
            O => \N__63062\,
            I => \N__63009\
        );

    \I__14678\ : LocalMux
    port map (
            O => \N__63059\,
            I => \N__63009\
        );

    \I__14677\ : LocalMux
    port map (
            O => \N__63056\,
            I => \N__63009\
        );

    \I__14676\ : Sp12to4
    port map (
            O => \N__63053\,
            I => \N__63009\
        );

    \I__14675\ : Sp12to4
    port map (
            O => \N__63050\,
            I => \N__63004\
        );

    \I__14674\ : Sp12to4
    port map (
            O => \N__63047\,
            I => \N__63004\
        );

    \I__14673\ : Sp12to4
    port map (
            O => \N__63044\,
            I => \N__63001\
        );

    \I__14672\ : Span4Mux_h
    port map (
            O => \N__63041\,
            I => \N__62998\
        );

    \I__14671\ : Span4Mux_v
    port map (
            O => \N__63036\,
            I => \N__62993\
        );

    \I__14670\ : Span4Mux_h
    port map (
            O => \N__63031\,
            I => \N__62993\
        );

    \I__14669\ : InMux
    port map (
            O => \N__63030\,
            I => \N__62986\
        );

    \I__14668\ : InMux
    port map (
            O => \N__63027\,
            I => \N__62986\
        );

    \I__14667\ : InMux
    port map (
            O => \N__63026\,
            I => \N__62986\
        );

    \I__14666\ : InMux
    port map (
            O => \N__63023\,
            I => \N__62981\
        );

    \I__14665\ : InMux
    port map (
            O => \N__63022\,
            I => \N__62981\
        );

    \I__14664\ : Span12Mux_h
    port map (
            O => \N__63009\,
            I => \N__62978\
        );

    \I__14663\ : Span12Mux_h
    port map (
            O => \N__63004\,
            I => \N__62973\
        );

    \I__14662\ : Span12Mux_v
    port map (
            O => \N__63001\,
            I => \N__62973\
        );

    \I__14661\ : Span4Mux_h
    port map (
            O => \N__62998\,
            I => \N__62968\
        );

    \I__14660\ : Span4Mux_v
    port map (
            O => \N__62993\,
            I => \N__62968\
        );

    \I__14659\ : LocalMux
    port map (
            O => \N__62986\,
            I => \aluParams_0\
        );

    \I__14658\ : LocalMux
    port map (
            O => \N__62981\,
            I => \aluParams_0\
        );

    \I__14657\ : Odrv12
    port map (
            O => \N__62978\,
            I => \aluParams_0\
        );

    \I__14656\ : Odrv12
    port map (
            O => \N__62973\,
            I => \aluParams_0\
        );

    \I__14655\ : Odrv4
    port map (
            O => \N__62968\,
            I => \aluParams_0\
        );

    \I__14654\ : CascadeMux
    port map (
            O => \N__62957\,
            I => \N__62953\
        );

    \I__14653\ : CascadeMux
    port map (
            O => \N__62956\,
            I => \N__62950\
        );

    \I__14652\ : InMux
    port map (
            O => \N__62953\,
            I => \N__62946\
        );

    \I__14651\ : InMux
    port map (
            O => \N__62950\,
            I => \N__62943\
        );

    \I__14650\ : CascadeMux
    port map (
            O => \N__62949\,
            I => \N__62940\
        );

    \I__14649\ : LocalMux
    port map (
            O => \N__62946\,
            I => \N__62936\
        );

    \I__14648\ : LocalMux
    port map (
            O => \N__62943\,
            I => \N__62933\
        );

    \I__14647\ : InMux
    port map (
            O => \N__62940\,
            I => \N__62928\
        );

    \I__14646\ : InMux
    port map (
            O => \N__62939\,
            I => \N__62928\
        );

    \I__14645\ : Span4Mux_h
    port map (
            O => \N__62936\,
            I => \N__62922\
        );

    \I__14644\ : Span4Mux_v
    port map (
            O => \N__62933\,
            I => \N__62922\
        );

    \I__14643\ : LocalMux
    port map (
            O => \N__62928\,
            I => \N__62919\
        );

    \I__14642\ : InMux
    port map (
            O => \N__62927\,
            I => \N__62916\
        );

    \I__14641\ : Span4Mux_h
    port map (
            O => \N__62922\,
            I => \N__62913\
        );

    \I__14640\ : Span4Mux_v
    port map (
            O => \N__62919\,
            I => \N__62910\
        );

    \I__14639\ : LocalMux
    port map (
            O => \N__62916\,
            I => \N__62907\
        );

    \I__14638\ : Span4Mux_h
    port map (
            O => \N__62913\,
            I => \N__62904\
        );

    \I__14637\ : Span4Mux_v
    port map (
            O => \N__62910\,
            I => \N__62899\
        );

    \I__14636\ : Span4Mux_h
    port map (
            O => \N__62907\,
            I => \N__62899\
        );

    \I__14635\ : Span4Mux_v
    port map (
            O => \N__62904\,
            I => \N__62894\
        );

    \I__14634\ : Span4Mux_h
    port map (
            O => \N__62899\,
            I => \N__62894\
        );

    \I__14633\ : Odrv4
    port map (
            O => \N__62894\,
            I => \ALU.combOperand2_0_9\
        );

    \I__14632\ : InMux
    port map (
            O => \N__62891\,
            I => \N__62878\
        );

    \I__14631\ : InMux
    port map (
            O => \N__62890\,
            I => \N__62875\
        );

    \I__14630\ : InMux
    port map (
            O => \N__62889\,
            I => \N__62868\
        );

    \I__14629\ : InMux
    port map (
            O => \N__62888\,
            I => \N__62863\
        );

    \I__14628\ : InMux
    port map (
            O => \N__62887\,
            I => \N__62863\
        );

    \I__14627\ : CascadeMux
    port map (
            O => \N__62886\,
            I => \N__62860\
        );

    \I__14626\ : InMux
    port map (
            O => \N__62885\,
            I => \N__62856\
        );

    \I__14625\ : InMux
    port map (
            O => \N__62884\,
            I => \N__62849\
        );

    \I__14624\ : InMux
    port map (
            O => \N__62883\,
            I => \N__62849\
        );

    \I__14623\ : InMux
    port map (
            O => \N__62882\,
            I => \N__62849\
        );

    \I__14622\ : InMux
    port map (
            O => \N__62881\,
            I => \N__62846\
        );

    \I__14621\ : LocalMux
    port map (
            O => \N__62878\,
            I => \N__62842\
        );

    \I__14620\ : LocalMux
    port map (
            O => \N__62875\,
            I => \N__62839\
        );

    \I__14619\ : InMux
    port map (
            O => \N__62874\,
            I => \N__62836\
        );

    \I__14618\ : InMux
    port map (
            O => \N__62873\,
            I => \N__62833\
        );

    \I__14617\ : InMux
    port map (
            O => \N__62872\,
            I => \N__62830\
        );

    \I__14616\ : InMux
    port map (
            O => \N__62871\,
            I => \N__62826\
        );

    \I__14615\ : LocalMux
    port map (
            O => \N__62868\,
            I => \N__62821\
        );

    \I__14614\ : LocalMux
    port map (
            O => \N__62863\,
            I => \N__62821\
        );

    \I__14613\ : InMux
    port map (
            O => \N__62860\,
            I => \N__62815\
        );

    \I__14612\ : InMux
    port map (
            O => \N__62859\,
            I => \N__62812\
        );

    \I__14611\ : LocalMux
    port map (
            O => \N__62856\,
            I => \N__62806\
        );

    \I__14610\ : LocalMux
    port map (
            O => \N__62849\,
            I => \N__62806\
        );

    \I__14609\ : LocalMux
    port map (
            O => \N__62846\,
            I => \N__62802\
        );

    \I__14608\ : InMux
    port map (
            O => \N__62845\,
            I => \N__62798\
        );

    \I__14607\ : Span4Mux_v
    port map (
            O => \N__62842\,
            I => \N__62793\
        );

    \I__14606\ : Span4Mux_v
    port map (
            O => \N__62839\,
            I => \N__62793\
        );

    \I__14605\ : LocalMux
    port map (
            O => \N__62836\,
            I => \N__62786\
        );

    \I__14604\ : LocalMux
    port map (
            O => \N__62833\,
            I => \N__62786\
        );

    \I__14603\ : LocalMux
    port map (
            O => \N__62830\,
            I => \N__62786\
        );

    \I__14602\ : InMux
    port map (
            O => \N__62829\,
            I => \N__62782\
        );

    \I__14601\ : LocalMux
    port map (
            O => \N__62826\,
            I => \N__62777\
        );

    \I__14600\ : Span4Mux_v
    port map (
            O => \N__62821\,
            I => \N__62777\
        );

    \I__14599\ : InMux
    port map (
            O => \N__62820\,
            I => \N__62774\
        );

    \I__14598\ : InMux
    port map (
            O => \N__62819\,
            I => \N__62769\
        );

    \I__14597\ : InMux
    port map (
            O => \N__62818\,
            I => \N__62769\
        );

    \I__14596\ : LocalMux
    port map (
            O => \N__62815\,
            I => \N__62766\
        );

    \I__14595\ : LocalMux
    port map (
            O => \N__62812\,
            I => \N__62761\
        );

    \I__14594\ : InMux
    port map (
            O => \N__62811\,
            I => \N__62758\
        );

    \I__14593\ : Span4Mux_h
    port map (
            O => \N__62806\,
            I => \N__62755\
        );

    \I__14592\ : InMux
    port map (
            O => \N__62805\,
            I => \N__62752\
        );

    \I__14591\ : Span4Mux_v
    port map (
            O => \N__62802\,
            I => \N__62749\
        );

    \I__14590\ : InMux
    port map (
            O => \N__62801\,
            I => \N__62746\
        );

    \I__14589\ : LocalMux
    port map (
            O => \N__62798\,
            I => \N__62739\
        );

    \I__14588\ : Span4Mux_h
    port map (
            O => \N__62793\,
            I => \N__62739\
        );

    \I__14587\ : Span4Mux_v
    port map (
            O => \N__62786\,
            I => \N__62739\
        );

    \I__14586\ : InMux
    port map (
            O => \N__62785\,
            I => \N__62736\
        );

    \I__14585\ : LocalMux
    port map (
            O => \N__62782\,
            I => \N__62733\
        );

    \I__14584\ : Span4Mux_h
    port map (
            O => \N__62777\,
            I => \N__62726\
        );

    \I__14583\ : LocalMux
    port map (
            O => \N__62774\,
            I => \N__62726\
        );

    \I__14582\ : LocalMux
    port map (
            O => \N__62769\,
            I => \N__62726\
        );

    \I__14581\ : Span4Mux_v
    port map (
            O => \N__62766\,
            I => \N__62723\
        );

    \I__14580\ : InMux
    port map (
            O => \N__62765\,
            I => \N__62718\
        );

    \I__14579\ : InMux
    port map (
            O => \N__62764\,
            I => \N__62718\
        );

    \I__14578\ : Span4Mux_v
    port map (
            O => \N__62761\,
            I => \N__62709\
        );

    \I__14577\ : LocalMux
    port map (
            O => \N__62758\,
            I => \N__62709\
        );

    \I__14576\ : Span4Mux_v
    port map (
            O => \N__62755\,
            I => \N__62709\
        );

    \I__14575\ : LocalMux
    port map (
            O => \N__62752\,
            I => \N__62709\
        );

    \I__14574\ : Sp12to4
    port map (
            O => \N__62749\,
            I => \N__62704\
        );

    \I__14573\ : LocalMux
    port map (
            O => \N__62746\,
            I => \N__62704\
        );

    \I__14572\ : Span4Mux_v
    port map (
            O => \N__62739\,
            I => \N__62701\
        );

    \I__14571\ : LocalMux
    port map (
            O => \N__62736\,
            I => \N__62698\
        );

    \I__14570\ : Span4Mux_h
    port map (
            O => \N__62733\,
            I => \N__62693\
        );

    \I__14569\ : Span4Mux_h
    port map (
            O => \N__62726\,
            I => \N__62693\
        );

    \I__14568\ : Span4Mux_v
    port map (
            O => \N__62723\,
            I => \N__62688\
        );

    \I__14567\ : LocalMux
    port map (
            O => \N__62718\,
            I => \N__62688\
        );

    \I__14566\ : Span4Mux_h
    port map (
            O => \N__62709\,
            I => \N__62685\
        );

    \I__14565\ : Odrv12
    port map (
            O => \N__62704\,
            I => \aluOut_9\
        );

    \I__14564\ : Odrv4
    port map (
            O => \N__62701\,
            I => \aluOut_9\
        );

    \I__14563\ : Odrv12
    port map (
            O => \N__62698\,
            I => \aluOut_9\
        );

    \I__14562\ : Odrv4
    port map (
            O => \N__62693\,
            I => \aluOut_9\
        );

    \I__14561\ : Odrv4
    port map (
            O => \N__62688\,
            I => \aluOut_9\
        );

    \I__14560\ : Odrv4
    port map (
            O => \N__62685\,
            I => \aluOut_9\
        );

    \I__14559\ : CascadeMux
    port map (
            O => \N__62672\,
            I => \N__62669\
        );

    \I__14558\ : InMux
    port map (
            O => \N__62669\,
            I => \N__62666\
        );

    \I__14557\ : LocalMux
    port map (
            O => \N__62666\,
            I => \ALU.d_RNI70I1IZ0Z_9\
        );

    \I__14556\ : InMux
    port map (
            O => \N__62663\,
            I => \N__62660\
        );

    \I__14555\ : LocalMux
    port map (
            O => \N__62660\,
            I => \N__62657\
        );

    \I__14554\ : Span4Mux_h
    port map (
            O => \N__62657\,
            I => \N__62652\
        );

    \I__14553\ : CascadeMux
    port map (
            O => \N__62656\,
            I => \N__62649\
        );

    \I__14552\ : InMux
    port map (
            O => \N__62655\,
            I => \N__62645\
        );

    \I__14551\ : Span4Mux_v
    port map (
            O => \N__62652\,
            I => \N__62642\
        );

    \I__14550\ : InMux
    port map (
            O => \N__62649\,
            I => \N__62639\
        );

    \I__14549\ : InMux
    port map (
            O => \N__62648\,
            I => \N__62636\
        );

    \I__14548\ : LocalMux
    port map (
            O => \N__62645\,
            I => \ALU.N_980\
        );

    \I__14547\ : Odrv4
    port map (
            O => \N__62642\,
            I => \ALU.N_980\
        );

    \I__14546\ : LocalMux
    port map (
            O => \N__62639\,
            I => \ALU.N_980\
        );

    \I__14545\ : LocalMux
    port map (
            O => \N__62636\,
            I => \ALU.N_980\
        );

    \I__14544\ : InMux
    port map (
            O => \N__62627\,
            I => \N__62624\
        );

    \I__14543\ : LocalMux
    port map (
            O => \N__62624\,
            I => \ALU.N_1029\
        );

    \I__14542\ : InMux
    port map (
            O => \N__62621\,
            I => \N__62618\
        );

    \I__14541\ : LocalMux
    port map (
            O => \N__62618\,
            I => \N__62615\
        );

    \I__14540\ : Span4Mux_h
    port map (
            O => \N__62615\,
            I => \N__62612\
        );

    \I__14539\ : Odrv4
    port map (
            O => \N__62612\,
            I => \PROM.ROMDATA.m500_ns_1\
        );

    \I__14538\ : InMux
    port map (
            O => \N__62609\,
            I => \N__62603\
        );

    \I__14537\ : InMux
    port map (
            O => \N__62608\,
            I => \N__62603\
        );

    \I__14536\ : LocalMux
    port map (
            O => \N__62603\,
            I => \N__62600\
        );

    \I__14535\ : Span4Mux_h
    port map (
            O => \N__62600\,
            I => \N__62597\
        );

    \I__14534\ : Span4Mux_h
    port map (
            O => \N__62597\,
            I => \N__62594\
        );

    \I__14533\ : Span4Mux_v
    port map (
            O => \N__62594\,
            I => \N__62591\
        );

    \I__14532\ : Odrv4
    port map (
            O => \N__62591\,
            I => \PROM.ROMDATA.m500_ns\
        );

    \I__14531\ : CascadeMux
    port map (
            O => \N__62588\,
            I => \N__62580\
        );

    \I__14530\ : InMux
    port map (
            O => \N__62587\,
            I => \N__62576\
        );

    \I__14529\ : InMux
    port map (
            O => \N__62586\,
            I => \N__62573\
        );

    \I__14528\ : CascadeMux
    port map (
            O => \N__62585\,
            I => \N__62567\
        );

    \I__14527\ : CascadeMux
    port map (
            O => \N__62584\,
            I => \N__62564\
        );

    \I__14526\ : InMux
    port map (
            O => \N__62583\,
            I => \N__62559\
        );

    \I__14525\ : InMux
    port map (
            O => \N__62580\,
            I => \N__62559\
        );

    \I__14524\ : CascadeMux
    port map (
            O => \N__62579\,
            I => \N__62553\
        );

    \I__14523\ : LocalMux
    port map (
            O => \N__62576\,
            I => \N__62547\
        );

    \I__14522\ : LocalMux
    port map (
            O => \N__62573\,
            I => \N__62544\
        );

    \I__14521\ : CascadeMux
    port map (
            O => \N__62572\,
            I => \N__62541\
        );

    \I__14520\ : InMux
    port map (
            O => \N__62571\,
            I => \N__62538\
        );

    \I__14519\ : InMux
    port map (
            O => \N__62570\,
            I => \N__62535\
        );

    \I__14518\ : InMux
    port map (
            O => \N__62567\,
            I => \N__62530\
        );

    \I__14517\ : InMux
    port map (
            O => \N__62564\,
            I => \N__62530\
        );

    \I__14516\ : LocalMux
    port map (
            O => \N__62559\,
            I => \N__62527\
        );

    \I__14515\ : InMux
    port map (
            O => \N__62558\,
            I => \N__62524\
        );

    \I__14514\ : CascadeMux
    port map (
            O => \N__62557\,
            I => \N__62520\
        );

    \I__14513\ : InMux
    port map (
            O => \N__62556\,
            I => \N__62515\
        );

    \I__14512\ : InMux
    port map (
            O => \N__62553\,
            I => \N__62512\
        );

    \I__14511\ : InMux
    port map (
            O => \N__62552\,
            I => \N__62507\
        );

    \I__14510\ : InMux
    port map (
            O => \N__62551\,
            I => \N__62507\
        );

    \I__14509\ : InMux
    port map (
            O => \N__62550\,
            I => \N__62499\
        );

    \I__14508\ : Span4Mux_v
    port map (
            O => \N__62547\,
            I => \N__62496\
        );

    \I__14507\ : Span4Mux_v
    port map (
            O => \N__62544\,
            I => \N__62493\
        );

    \I__14506\ : InMux
    port map (
            O => \N__62541\,
            I => \N__62490\
        );

    \I__14505\ : LocalMux
    port map (
            O => \N__62538\,
            I => \N__62487\
        );

    \I__14504\ : LocalMux
    port map (
            O => \N__62535\,
            I => \N__62482\
        );

    \I__14503\ : LocalMux
    port map (
            O => \N__62530\,
            I => \N__62482\
        );

    \I__14502\ : Span4Mux_v
    port map (
            O => \N__62527\,
            I => \N__62479\
        );

    \I__14501\ : LocalMux
    port map (
            O => \N__62524\,
            I => \N__62476\
        );

    \I__14500\ : InMux
    port map (
            O => \N__62523\,
            I => \N__62473\
        );

    \I__14499\ : InMux
    port map (
            O => \N__62520\,
            I => \N__62468\
        );

    \I__14498\ : InMux
    port map (
            O => \N__62519\,
            I => \N__62468\
        );

    \I__14497\ : InMux
    port map (
            O => \N__62518\,
            I => \N__62465\
        );

    \I__14496\ : LocalMux
    port map (
            O => \N__62515\,
            I => \N__62462\
        );

    \I__14495\ : LocalMux
    port map (
            O => \N__62512\,
            I => \N__62459\
        );

    \I__14494\ : LocalMux
    port map (
            O => \N__62507\,
            I => \N__62456\
        );

    \I__14493\ : InMux
    port map (
            O => \N__62506\,
            I => \N__62447\
        );

    \I__14492\ : InMux
    port map (
            O => \N__62505\,
            I => \N__62447\
        );

    \I__14491\ : InMux
    port map (
            O => \N__62504\,
            I => \N__62447\
        );

    \I__14490\ : InMux
    port map (
            O => \N__62503\,
            I => \N__62447\
        );

    \I__14489\ : InMux
    port map (
            O => \N__62502\,
            I => \N__62444\
        );

    \I__14488\ : LocalMux
    port map (
            O => \N__62499\,
            I => \N__62441\
        );

    \I__14487\ : Span4Mux_v
    port map (
            O => \N__62496\,
            I => \N__62436\
        );

    \I__14486\ : Span4Mux_h
    port map (
            O => \N__62493\,
            I => \N__62436\
        );

    \I__14485\ : LocalMux
    port map (
            O => \N__62490\,
            I => \N__62433\
        );

    \I__14484\ : Span4Mux_v
    port map (
            O => \N__62487\,
            I => \N__62430\
        );

    \I__14483\ : Span4Mux_h
    port map (
            O => \N__62482\,
            I => \N__62427\
        );

    \I__14482\ : Span4Mux_h
    port map (
            O => \N__62479\,
            I => \N__62422\
        );

    \I__14481\ : Span4Mux_v
    port map (
            O => \N__62476\,
            I => \N__62422\
        );

    \I__14480\ : LocalMux
    port map (
            O => \N__62473\,
            I => \N__62417\
        );

    \I__14479\ : LocalMux
    port map (
            O => \N__62468\,
            I => \N__62417\
        );

    \I__14478\ : LocalMux
    port map (
            O => \N__62465\,
            I => \N__62414\
        );

    \I__14477\ : Span4Mux_v
    port map (
            O => \N__62462\,
            I => \N__62411\
        );

    \I__14476\ : Span4Mux_h
    port map (
            O => \N__62459\,
            I => \N__62402\
        );

    \I__14475\ : Span4Mux_v
    port map (
            O => \N__62456\,
            I => \N__62402\
        );

    \I__14474\ : LocalMux
    port map (
            O => \N__62447\,
            I => \N__62402\
        );

    \I__14473\ : LocalMux
    port map (
            O => \N__62444\,
            I => \N__62402\
        );

    \I__14472\ : Span12Mux_h
    port map (
            O => \N__62441\,
            I => \N__62399\
        );

    \I__14471\ : Span4Mux_h
    port map (
            O => \N__62436\,
            I => \N__62392\
        );

    \I__14470\ : Span4Mux_h
    port map (
            O => \N__62433\,
            I => \N__62392\
        );

    \I__14469\ : Span4Mux_v
    port map (
            O => \N__62430\,
            I => \N__62392\
        );

    \I__14468\ : Span4Mux_v
    port map (
            O => \N__62427\,
            I => \N__62389\
        );

    \I__14467\ : Span4Mux_h
    port map (
            O => \N__62422\,
            I => \N__62382\
        );

    \I__14466\ : Span4Mux_v
    port map (
            O => \N__62417\,
            I => \N__62382\
        );

    \I__14465\ : Span4Mux_h
    port map (
            O => \N__62414\,
            I => \N__62382\
        );

    \I__14464\ : Span4Mux_v
    port map (
            O => \N__62411\,
            I => \N__62377\
        );

    \I__14463\ : Span4Mux_v
    port map (
            O => \N__62402\,
            I => \N__62377\
        );

    \I__14462\ : Odrv12
    port map (
            O => \N__62399\,
            I => \aluOut_6\
        );

    \I__14461\ : Odrv4
    port map (
            O => \N__62392\,
            I => \aluOut_6\
        );

    \I__14460\ : Odrv4
    port map (
            O => \N__62389\,
            I => \aluOut_6\
        );

    \I__14459\ : Odrv4
    port map (
            O => \N__62382\,
            I => \aluOut_6\
        );

    \I__14458\ : Odrv4
    port map (
            O => \N__62377\,
            I => \aluOut_6\
        );

    \I__14457\ : CascadeMux
    port map (
            O => \N__62366\,
            I => \N__62363\
        );

    \I__14456\ : InMux
    port map (
            O => \N__62363\,
            I => \N__62360\
        );

    \I__14455\ : LocalMux
    port map (
            O => \N__62360\,
            I => \N__62357\
        );

    \I__14454\ : Span4Mux_v
    port map (
            O => \N__62357\,
            I => \N__62354\
        );

    \I__14453\ : Span4Mux_h
    port map (
            O => \N__62354\,
            I => \N__62351\
        );

    \I__14452\ : Sp12to4
    port map (
            O => \N__62351\,
            I => \N__62348\
        );

    \I__14451\ : Odrv12
    port map (
            O => \N__62348\,
            I => \ALU.d_RNIALE3IZ0Z_6\
        );

    \I__14450\ : InMux
    port map (
            O => \N__62345\,
            I => \N__62342\
        );

    \I__14449\ : LocalMux
    port map (
            O => \N__62342\,
            I => \N__62339\
        );

    \I__14448\ : Span4Mux_h
    port map (
            O => \N__62339\,
            I => \N__62335\
        );

    \I__14447\ : InMux
    port map (
            O => \N__62338\,
            I => \N__62332\
        );

    \I__14446\ : Odrv4
    port map (
            O => \N__62335\,
            I => \ALU.addsub_6\
        );

    \I__14445\ : LocalMux
    port map (
            O => \N__62332\,
            I => \ALU.addsub_6\
        );

    \I__14444\ : InMux
    port map (
            O => \N__62327\,
            I => \ALU.addsub_cry_5\
        );

    \I__14443\ : CascadeMux
    port map (
            O => \N__62324\,
            I => \N__62321\
        );

    \I__14442\ : InMux
    port map (
            O => \N__62321\,
            I => \N__62317\
        );

    \I__14441\ : CascadeMux
    port map (
            O => \N__62320\,
            I => \N__62311\
        );

    \I__14440\ : LocalMux
    port map (
            O => \N__62317\,
            I => \N__62308\
        );

    \I__14439\ : CascadeMux
    port map (
            O => \N__62316\,
            I => \N__62303\
        );

    \I__14438\ : CascadeMux
    port map (
            O => \N__62315\,
            I => \N__62299\
        );

    \I__14437\ : InMux
    port map (
            O => \N__62314\,
            I => \N__62295\
        );

    \I__14436\ : InMux
    port map (
            O => \N__62311\,
            I => \N__62292\
        );

    \I__14435\ : Span4Mux_v
    port map (
            O => \N__62308\,
            I => \N__62289\
        );

    \I__14434\ : InMux
    port map (
            O => \N__62307\,
            I => \N__62286\
        );

    \I__14433\ : CascadeMux
    port map (
            O => \N__62306\,
            I => \N__62282\
        );

    \I__14432\ : InMux
    port map (
            O => \N__62303\,
            I => \N__62278\
        );

    \I__14431\ : CascadeMux
    port map (
            O => \N__62302\,
            I => \N__62275\
        );

    \I__14430\ : InMux
    port map (
            O => \N__62299\,
            I => \N__62266\
        );

    \I__14429\ : InMux
    port map (
            O => \N__62298\,
            I => \N__62262\
        );

    \I__14428\ : LocalMux
    port map (
            O => \N__62295\,
            I => \N__62256\
        );

    \I__14427\ : LocalMux
    port map (
            O => \N__62292\,
            I => \N__62256\
        );

    \I__14426\ : Span4Mux_h
    port map (
            O => \N__62289\,
            I => \N__62251\
        );

    \I__14425\ : LocalMux
    port map (
            O => \N__62286\,
            I => \N__62251\
        );

    \I__14424\ : InMux
    port map (
            O => \N__62285\,
            I => \N__62244\
        );

    \I__14423\ : InMux
    port map (
            O => \N__62282\,
            I => \N__62244\
        );

    \I__14422\ : InMux
    port map (
            O => \N__62281\,
            I => \N__62244\
        );

    \I__14421\ : LocalMux
    port map (
            O => \N__62278\,
            I => \N__62241\
        );

    \I__14420\ : InMux
    port map (
            O => \N__62275\,
            I => \N__62238\
        );

    \I__14419\ : InMux
    port map (
            O => \N__62274\,
            I => \N__62235\
        );

    \I__14418\ : InMux
    port map (
            O => \N__62273\,
            I => \N__62223\
        );

    \I__14417\ : InMux
    port map (
            O => \N__62272\,
            I => \N__62223\
        );

    \I__14416\ : InMux
    port map (
            O => \N__62271\,
            I => \N__62223\
        );

    \I__14415\ : InMux
    port map (
            O => \N__62270\,
            I => \N__62223\
        );

    \I__14414\ : InMux
    port map (
            O => \N__62269\,
            I => \N__62220\
        );

    \I__14413\ : LocalMux
    port map (
            O => \N__62266\,
            I => \N__62216\
        );

    \I__14412\ : InMux
    port map (
            O => \N__62265\,
            I => \N__62213\
        );

    \I__14411\ : LocalMux
    port map (
            O => \N__62262\,
            I => \N__62210\
        );

    \I__14410\ : InMux
    port map (
            O => \N__62261\,
            I => \N__62206\
        );

    \I__14409\ : Span4Mux_v
    port map (
            O => \N__62256\,
            I => \N__62199\
        );

    \I__14408\ : Span4Mux_h
    port map (
            O => \N__62251\,
            I => \N__62199\
        );

    \I__14407\ : LocalMux
    port map (
            O => \N__62244\,
            I => \N__62199\
        );

    \I__14406\ : Span4Mux_v
    port map (
            O => \N__62241\,
            I => \N__62192\
        );

    \I__14405\ : LocalMux
    port map (
            O => \N__62238\,
            I => \N__62192\
        );

    \I__14404\ : LocalMux
    port map (
            O => \N__62235\,
            I => \N__62192\
        );

    \I__14403\ : CascadeMux
    port map (
            O => \N__62234\,
            I => \N__62187\
        );

    \I__14402\ : InMux
    port map (
            O => \N__62233\,
            I => \N__62182\
        );

    \I__14401\ : InMux
    port map (
            O => \N__62232\,
            I => \N__62179\
        );

    \I__14400\ : LocalMux
    port map (
            O => \N__62223\,
            I => \N__62176\
        );

    \I__14399\ : LocalMux
    port map (
            O => \N__62220\,
            I => \N__62173\
        );

    \I__14398\ : InMux
    port map (
            O => \N__62219\,
            I => \N__62170\
        );

    \I__14397\ : Span4Mux_v
    port map (
            O => \N__62216\,
            I => \N__62165\
        );

    \I__14396\ : LocalMux
    port map (
            O => \N__62213\,
            I => \N__62165\
        );

    \I__14395\ : Span4Mux_v
    port map (
            O => \N__62210\,
            I => \N__62162\
        );

    \I__14394\ : InMux
    port map (
            O => \N__62209\,
            I => \N__62159\
        );

    \I__14393\ : LocalMux
    port map (
            O => \N__62206\,
            I => \N__62151\
        );

    \I__14392\ : Span4Mux_v
    port map (
            O => \N__62199\,
            I => \N__62151\
        );

    \I__14391\ : Span4Mux_v
    port map (
            O => \N__62192\,
            I => \N__62148\
        );

    \I__14390\ : InMux
    port map (
            O => \N__62191\,
            I => \N__62143\
        );

    \I__14389\ : InMux
    port map (
            O => \N__62190\,
            I => \N__62143\
        );

    \I__14388\ : InMux
    port map (
            O => \N__62187\,
            I => \N__62138\
        );

    \I__14387\ : InMux
    port map (
            O => \N__62186\,
            I => \N__62138\
        );

    \I__14386\ : InMux
    port map (
            O => \N__62185\,
            I => \N__62135\
        );

    \I__14385\ : LocalMux
    port map (
            O => \N__62182\,
            I => \N__62132\
        );

    \I__14384\ : LocalMux
    port map (
            O => \N__62179\,
            I => \N__62125\
        );

    \I__14383\ : Span4Mux_h
    port map (
            O => \N__62176\,
            I => \N__62125\
        );

    \I__14382\ : Span4Mux_v
    port map (
            O => \N__62173\,
            I => \N__62125\
        );

    \I__14381\ : LocalMux
    port map (
            O => \N__62170\,
            I => \N__62122\
        );

    \I__14380\ : Span4Mux_v
    port map (
            O => \N__62165\,
            I => \N__62119\
        );

    \I__14379\ : Span4Mux_h
    port map (
            O => \N__62162\,
            I => \N__62114\
        );

    \I__14378\ : LocalMux
    port map (
            O => \N__62159\,
            I => \N__62114\
        );

    \I__14377\ : InMux
    port map (
            O => \N__62158\,
            I => \N__62107\
        );

    \I__14376\ : InMux
    port map (
            O => \N__62157\,
            I => \N__62107\
        );

    \I__14375\ : InMux
    port map (
            O => \N__62156\,
            I => \N__62107\
        );

    \I__14374\ : Span4Mux_v
    port map (
            O => \N__62151\,
            I => \N__62100\
        );

    \I__14373\ : Span4Mux_h
    port map (
            O => \N__62148\,
            I => \N__62100\
        );

    \I__14372\ : LocalMux
    port map (
            O => \N__62143\,
            I => \N__62100\
        );

    \I__14371\ : LocalMux
    port map (
            O => \N__62138\,
            I => \N__62095\
        );

    \I__14370\ : LocalMux
    port map (
            O => \N__62135\,
            I => \N__62095\
        );

    \I__14369\ : Span4Mux_v
    port map (
            O => \N__62132\,
            I => \N__62090\
        );

    \I__14368\ : Span4Mux_h
    port map (
            O => \N__62125\,
            I => \N__62090\
        );

    \I__14367\ : Span4Mux_h
    port map (
            O => \N__62122\,
            I => \N__62087\
        );

    \I__14366\ : Span4Mux_h
    port map (
            O => \N__62119\,
            I => \N__62084\
        );

    \I__14365\ : Span4Mux_v
    port map (
            O => \N__62114\,
            I => \N__62079\
        );

    \I__14364\ : LocalMux
    port map (
            O => \N__62107\,
            I => \N__62079\
        );

    \I__14363\ : Span4Mux_h
    port map (
            O => \N__62100\,
            I => \N__62076\
        );

    \I__14362\ : Span12Mux_h
    port map (
            O => \N__62095\,
            I => \N__62071\
        );

    \I__14361\ : Sp12to4
    port map (
            O => \N__62090\,
            I => \N__62071\
        );

    \I__14360\ : Odrv4
    port map (
            O => \N__62087\,
            I => \aluOut_7\
        );

    \I__14359\ : Odrv4
    port map (
            O => \N__62084\,
            I => \aluOut_7\
        );

    \I__14358\ : Odrv4
    port map (
            O => \N__62079\,
            I => \aluOut_7\
        );

    \I__14357\ : Odrv4
    port map (
            O => \N__62076\,
            I => \aluOut_7\
        );

    \I__14356\ : Odrv12
    port map (
            O => \N__62071\,
            I => \aluOut_7\
        );

    \I__14355\ : CascadeMux
    port map (
            O => \N__62060\,
            I => \N__62057\
        );

    \I__14354\ : InMux
    port map (
            O => \N__62057\,
            I => \N__62054\
        );

    \I__14353\ : LocalMux
    port map (
            O => \N__62054\,
            I => \N__62051\
        );

    \I__14352\ : Odrv12
    port map (
            O => \N__62051\,
            I => \ALU.d_RNI500DGZ0Z_7\
        );

    \I__14351\ : InMux
    port map (
            O => \N__62048\,
            I => \N__62044\
        );

    \I__14350\ : InMux
    port map (
            O => \N__62047\,
            I => \N__62041\
        );

    \I__14349\ : LocalMux
    port map (
            O => \N__62044\,
            I => \N__62038\
        );

    \I__14348\ : LocalMux
    port map (
            O => \N__62041\,
            I => \N__62035\
        );

    \I__14347\ : Odrv4
    port map (
            O => \N__62038\,
            I => \ALU.addsub_7\
        );

    \I__14346\ : Odrv4
    port map (
            O => \N__62035\,
            I => \ALU.addsub_7\
        );

    \I__14345\ : InMux
    port map (
            O => \N__62030\,
            I => \bfn_23_15_0_\
        );

    \I__14344\ : InMux
    port map (
            O => \N__62027\,
            I => \N__62018\
        );

    \I__14343\ : CascadeMux
    port map (
            O => \N__62026\,
            I => \N__62014\
        );

    \I__14342\ : CascadeMux
    port map (
            O => \N__62025\,
            I => \N__62011\
        );

    \I__14341\ : InMux
    port map (
            O => \N__62024\,
            I => \N__62007\
        );

    \I__14340\ : InMux
    port map (
            O => \N__62023\,
            I => \N__62004\
        );

    \I__14339\ : CascadeMux
    port map (
            O => \N__62022\,
            I => \N__62001\
        );

    \I__14338\ : CascadeMux
    port map (
            O => \N__62021\,
            I => \N__61997\
        );

    \I__14337\ : LocalMux
    port map (
            O => \N__62018\,
            I => \N__61994\
        );

    \I__14336\ : InMux
    port map (
            O => \N__62017\,
            I => \N__61991\
        );

    \I__14335\ : InMux
    port map (
            O => \N__62014\,
            I => \N__61984\
        );

    \I__14334\ : InMux
    port map (
            O => \N__62011\,
            I => \N__61984\
        );

    \I__14333\ : InMux
    port map (
            O => \N__62010\,
            I => \N__61984\
        );

    \I__14332\ : LocalMux
    port map (
            O => \N__62007\,
            I => \N__61979\
        );

    \I__14331\ : LocalMux
    port map (
            O => \N__62004\,
            I => \N__61972\
        );

    \I__14330\ : InMux
    port map (
            O => \N__62001\,
            I => \N__61969\
        );

    \I__14329\ : CascadeMux
    port map (
            O => \N__62000\,
            I => \N__61966\
        );

    \I__14328\ : InMux
    port map (
            O => \N__61997\,
            I => \N__61963\
        );

    \I__14327\ : Span4Mux_h
    port map (
            O => \N__61994\,
            I => \N__61960\
        );

    \I__14326\ : LocalMux
    port map (
            O => \N__61991\,
            I => \N__61955\
        );

    \I__14325\ : LocalMux
    port map (
            O => \N__61984\,
            I => \N__61955\
        );

    \I__14324\ : InMux
    port map (
            O => \N__61983\,
            I => \N__61952\
        );

    \I__14323\ : CascadeMux
    port map (
            O => \N__61982\,
            I => \N__61949\
        );

    \I__14322\ : Span4Mux_h
    port map (
            O => \N__61979\,
            I => \N__61944\
        );

    \I__14321\ : InMux
    port map (
            O => \N__61978\,
            I => \N__61939\
        );

    \I__14320\ : InMux
    port map (
            O => \N__61977\,
            I => \N__61939\
        );

    \I__14319\ : CascadeMux
    port map (
            O => \N__61976\,
            I => \N__61936\
        );

    \I__14318\ : CascadeMux
    port map (
            O => \N__61975\,
            I => \N__61932\
        );

    \I__14317\ : Span4Mux_h
    port map (
            O => \N__61972\,
            I => \N__61925\
        );

    \I__14316\ : LocalMux
    port map (
            O => \N__61969\,
            I => \N__61925\
        );

    \I__14315\ : InMux
    port map (
            O => \N__61966\,
            I => \N__61922\
        );

    \I__14314\ : LocalMux
    port map (
            O => \N__61963\,
            I => \N__61919\
        );

    \I__14313\ : Span4Mux_v
    port map (
            O => \N__61960\,
            I => \N__61914\
        );

    \I__14312\ : Span4Mux_v
    port map (
            O => \N__61955\,
            I => \N__61914\
        );

    \I__14311\ : LocalMux
    port map (
            O => \N__61952\,
            I => \N__61911\
        );

    \I__14310\ : InMux
    port map (
            O => \N__61949\,
            I => \N__61908\
        );

    \I__14309\ : CascadeMux
    port map (
            O => \N__61948\,
            I => \N__61905\
        );

    \I__14308\ : InMux
    port map (
            O => \N__61947\,
            I => \N__61902\
        );

    \I__14307\ : Span4Mux_h
    port map (
            O => \N__61944\,
            I => \N__61896\
        );

    \I__14306\ : LocalMux
    port map (
            O => \N__61939\,
            I => \N__61896\
        );

    \I__14305\ : InMux
    port map (
            O => \N__61936\,
            I => \N__61893\
        );

    \I__14304\ : InMux
    port map (
            O => \N__61935\,
            I => \N__61890\
        );

    \I__14303\ : InMux
    port map (
            O => \N__61932\,
            I => \N__61887\
        );

    \I__14302\ : InMux
    port map (
            O => \N__61931\,
            I => \N__61882\
        );

    \I__14301\ : InMux
    port map (
            O => \N__61930\,
            I => \N__61882\
        );

    \I__14300\ : Span4Mux_h
    port map (
            O => \N__61925\,
            I => \N__61878\
        );

    \I__14299\ : LocalMux
    port map (
            O => \N__61922\,
            I => \N__61869\
        );

    \I__14298\ : Span4Mux_h
    port map (
            O => \N__61919\,
            I => \N__61869\
        );

    \I__14297\ : Span4Mux_h
    port map (
            O => \N__61914\,
            I => \N__61869\
        );

    \I__14296\ : Span4Mux_v
    port map (
            O => \N__61911\,
            I => \N__61869\
        );

    \I__14295\ : LocalMux
    port map (
            O => \N__61908\,
            I => \N__61866\
        );

    \I__14294\ : InMux
    port map (
            O => \N__61905\,
            I => \N__61863\
        );

    \I__14293\ : LocalMux
    port map (
            O => \N__61902\,
            I => \N__61860\
        );

    \I__14292\ : InMux
    port map (
            O => \N__61901\,
            I => \N__61857\
        );

    \I__14291\ : Span4Mux_h
    port map (
            O => \N__61896\,
            I => \N__61852\
        );

    \I__14290\ : LocalMux
    port map (
            O => \N__61893\,
            I => \N__61852\
        );

    \I__14289\ : LocalMux
    port map (
            O => \N__61890\,
            I => \N__61849\
        );

    \I__14288\ : LocalMux
    port map (
            O => \N__61887\,
            I => \N__61846\
        );

    \I__14287\ : LocalMux
    port map (
            O => \N__61882\,
            I => \N__61843\
        );

    \I__14286\ : InMux
    port map (
            O => \N__61881\,
            I => \N__61840\
        );

    \I__14285\ : Span4Mux_v
    port map (
            O => \N__61878\,
            I => \N__61837\
        );

    \I__14284\ : Span4Mux_h
    port map (
            O => \N__61869\,
            I => \N__61833\
        );

    \I__14283\ : Span4Mux_h
    port map (
            O => \N__61866\,
            I => \N__61830\
        );

    \I__14282\ : LocalMux
    port map (
            O => \N__61863\,
            I => \N__61827\
        );

    \I__14281\ : Span4Mux_h
    port map (
            O => \N__61860\,
            I => \N__61820\
        );

    \I__14280\ : LocalMux
    port map (
            O => \N__61857\,
            I => \N__61820\
        );

    \I__14279\ : Span4Mux_v
    port map (
            O => \N__61852\,
            I => \N__61820\
        );

    \I__14278\ : Span12Mux_v
    port map (
            O => \N__61849\,
            I => \N__61817\
        );

    \I__14277\ : Span4Mux_v
    port map (
            O => \N__61846\,
            I => \N__61812\
        );

    \I__14276\ : Span4Mux_h
    port map (
            O => \N__61843\,
            I => \N__61812\
        );

    \I__14275\ : LocalMux
    port map (
            O => \N__61840\,
            I => \N__61807\
        );

    \I__14274\ : Span4Mux_v
    port map (
            O => \N__61837\,
            I => \N__61807\
        );

    \I__14273\ : InMux
    port map (
            O => \N__61836\,
            I => \N__61804\
        );

    \I__14272\ : Span4Mux_v
    port map (
            O => \N__61833\,
            I => \N__61799\
        );

    \I__14271\ : Span4Mux_h
    port map (
            O => \N__61830\,
            I => \N__61799\
        );

    \I__14270\ : Span4Mux_h
    port map (
            O => \N__61827\,
            I => \N__61794\
        );

    \I__14269\ : Span4Mux_v
    port map (
            O => \N__61820\,
            I => \N__61794\
        );

    \I__14268\ : Odrv12
    port map (
            O => \N__61817\,
            I => \aluOut_8\
        );

    \I__14267\ : Odrv4
    port map (
            O => \N__61812\,
            I => \aluOut_8\
        );

    \I__14266\ : Odrv4
    port map (
            O => \N__61807\,
            I => \aluOut_8\
        );

    \I__14265\ : LocalMux
    port map (
            O => \N__61804\,
            I => \aluOut_8\
        );

    \I__14264\ : Odrv4
    port map (
            O => \N__61799\,
            I => \aluOut_8\
        );

    \I__14263\ : Odrv4
    port map (
            O => \N__61794\,
            I => \aluOut_8\
        );

    \I__14262\ : CascadeMux
    port map (
            O => \N__61781\,
            I => \N__61778\
        );

    \I__14261\ : InMux
    port map (
            O => \N__61778\,
            I => \N__61775\
        );

    \I__14260\ : LocalMux
    port map (
            O => \N__61775\,
            I => \N__61772\
        );

    \I__14259\ : Span4Mux_h
    port map (
            O => \N__61772\,
            I => \N__61769\
        );

    \I__14258\ : Span4Mux_v
    port map (
            O => \N__61769\,
            I => \N__61766\
        );

    \I__14257\ : Span4Mux_h
    port map (
            O => \N__61766\,
            I => \N__61763\
        );

    \I__14256\ : Odrv4
    port map (
            O => \N__61763\,
            I => \ALU.d_RNIAJ1KHZ0Z_8\
        );

    \I__14255\ : InMux
    port map (
            O => \N__61760\,
            I => \N__61757\
        );

    \I__14254\ : LocalMux
    port map (
            O => \N__61757\,
            I => \N__61754\
        );

    \I__14253\ : Span4Mux_v
    port map (
            O => \N__61754\,
            I => \N__61750\
        );

    \I__14252\ : InMux
    port map (
            O => \N__61753\,
            I => \N__61747\
        );

    \I__14251\ : Odrv4
    port map (
            O => \N__61750\,
            I => \ALU.addsub_8\
        );

    \I__14250\ : LocalMux
    port map (
            O => \N__61747\,
            I => \ALU.addsub_8\
        );

    \I__14249\ : InMux
    port map (
            O => \N__61742\,
            I => \ALU.addsub_cry_7\
        );

    \I__14248\ : InMux
    port map (
            O => \N__61739\,
            I => \ALU.addsub_cry_8\
        );

    \I__14247\ : InMux
    port map (
            O => \N__61736\,
            I => \N__61733\
        );

    \I__14246\ : LocalMux
    port map (
            O => \N__61733\,
            I => \N__61730\
        );

    \I__14245\ : Span4Mux_v
    port map (
            O => \N__61730\,
            I => \N__61727\
        );

    \I__14244\ : Sp12to4
    port map (
            O => \N__61727\,
            I => \N__61724\
        );

    \I__14243\ : Span12Mux_h
    port map (
            O => \N__61724\,
            I => \N__61721\
        );

    \I__14242\ : Odrv12
    port map (
            O => \N__61721\,
            I => \ALU.c_RNI1QK5KZ0Z_10\
        );

    \I__14241\ : CascadeMux
    port map (
            O => \N__61718\,
            I => \N__61711\
        );

    \I__14240\ : CascadeMux
    port map (
            O => \N__61717\,
            I => \N__61707\
        );

    \I__14239\ : CascadeMux
    port map (
            O => \N__61716\,
            I => \N__61704\
        );

    \I__14238\ : CascadeMux
    port map (
            O => \N__61715\,
            I => \N__61698\
        );

    \I__14237\ : InMux
    port map (
            O => \N__61714\,
            I => \N__61692\
        );

    \I__14236\ : InMux
    port map (
            O => \N__61711\,
            I => \N__61692\
        );

    \I__14235\ : CascadeMux
    port map (
            O => \N__61710\,
            I => \N__61689\
        );

    \I__14234\ : InMux
    port map (
            O => \N__61707\,
            I => \N__61686\
        );

    \I__14233\ : InMux
    port map (
            O => \N__61704\,
            I => \N__61683\
        );

    \I__14232\ : InMux
    port map (
            O => \N__61703\,
            I => \N__61676\
        );

    \I__14231\ : InMux
    port map (
            O => \N__61702\,
            I => \N__61676\
        );

    \I__14230\ : InMux
    port map (
            O => \N__61701\,
            I => \N__61672\
        );

    \I__14229\ : InMux
    port map (
            O => \N__61698\,
            I => \N__61669\
        );

    \I__14228\ : InMux
    port map (
            O => \N__61697\,
            I => \N__61663\
        );

    \I__14227\ : LocalMux
    port map (
            O => \N__61692\,
            I => \N__61658\
        );

    \I__14226\ : InMux
    port map (
            O => \N__61689\,
            I => \N__61655\
        );

    \I__14225\ : LocalMux
    port map (
            O => \N__61686\,
            I => \N__61650\
        );

    \I__14224\ : LocalMux
    port map (
            O => \N__61683\,
            I => \N__61650\
        );

    \I__14223\ : InMux
    port map (
            O => \N__61682\,
            I => \N__61647\
        );

    \I__14222\ : InMux
    port map (
            O => \N__61681\,
            I => \N__61644\
        );

    \I__14221\ : LocalMux
    port map (
            O => \N__61676\,
            I => \N__61641\
        );

    \I__14220\ : CascadeMux
    port map (
            O => \N__61675\,
            I => \N__61637\
        );

    \I__14219\ : LocalMux
    port map (
            O => \N__61672\,
            I => \N__61633\
        );

    \I__14218\ : LocalMux
    port map (
            O => \N__61669\,
            I => \N__61630\
        );

    \I__14217\ : CascadeMux
    port map (
            O => \N__61668\,
            I => \N__61627\
        );

    \I__14216\ : InMux
    port map (
            O => \N__61667\,
            I => \N__61624\
        );

    \I__14215\ : InMux
    port map (
            O => \N__61666\,
            I => \N__61621\
        );

    \I__14214\ : LocalMux
    port map (
            O => \N__61663\,
            I => \N__61618\
        );

    \I__14213\ : InMux
    port map (
            O => \N__61662\,
            I => \N__61613\
        );

    \I__14212\ : InMux
    port map (
            O => \N__61661\,
            I => \N__61613\
        );

    \I__14211\ : Span4Mux_v
    port map (
            O => \N__61658\,
            I => \N__61610\
        );

    \I__14210\ : LocalMux
    port map (
            O => \N__61655\,
            I => \N__61607\
        );

    \I__14209\ : Span4Mux_v
    port map (
            O => \N__61650\,
            I => \N__61604\
        );

    \I__14208\ : LocalMux
    port map (
            O => \N__61647\,
            I => \N__61599\
        );

    \I__14207\ : LocalMux
    port map (
            O => \N__61644\,
            I => \N__61599\
        );

    \I__14206\ : Span4Mux_h
    port map (
            O => \N__61641\,
            I => \N__61596\
        );

    \I__14205\ : InMux
    port map (
            O => \N__61640\,
            I => \N__61593\
        );

    \I__14204\ : InMux
    port map (
            O => \N__61637\,
            I => \N__61588\
        );

    \I__14203\ : InMux
    port map (
            O => \N__61636\,
            I => \N__61588\
        );

    \I__14202\ : Span4Mux_v
    port map (
            O => \N__61633\,
            I => \N__61583\
        );

    \I__14201\ : Span4Mux_v
    port map (
            O => \N__61630\,
            I => \N__61583\
        );

    \I__14200\ : InMux
    port map (
            O => \N__61627\,
            I => \N__61580\
        );

    \I__14199\ : LocalMux
    port map (
            O => \N__61624\,
            I => \N__61577\
        );

    \I__14198\ : LocalMux
    port map (
            O => \N__61621\,
            I => \N__61574\
        );

    \I__14197\ : Span4Mux_h
    port map (
            O => \N__61618\,
            I => \N__61571\
        );

    \I__14196\ : LocalMux
    port map (
            O => \N__61613\,
            I => \N__61568\
        );

    \I__14195\ : Sp12to4
    port map (
            O => \N__61610\,
            I => \N__61565\
        );

    \I__14194\ : Span4Mux_v
    port map (
            O => \N__61607\,
            I => \N__61562\
        );

    \I__14193\ : Span4Mux_v
    port map (
            O => \N__61604\,
            I => \N__61559\
        );

    \I__14192\ : Span4Mux_v
    port map (
            O => \N__61599\,
            I => \N__61556\
        );

    \I__14191\ : Span4Mux_h
    port map (
            O => \N__61596\,
            I => \N__61553\
        );

    \I__14190\ : LocalMux
    port map (
            O => \N__61593\,
            I => \N__61546\
        );

    \I__14189\ : LocalMux
    port map (
            O => \N__61588\,
            I => \N__61546\
        );

    \I__14188\ : Sp12to4
    port map (
            O => \N__61583\,
            I => \N__61546\
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__61580\,
            I => \N__61541\
        );

    \I__14186\ : Span4Mux_h
    port map (
            O => \N__61577\,
            I => \N__61541\
        );

    \I__14185\ : Span4Mux_v
    port map (
            O => \N__61574\,
            I => \N__61536\
        );

    \I__14184\ : Span4Mux_h
    port map (
            O => \N__61571\,
            I => \N__61536\
        );

    \I__14183\ : Span4Mux_h
    port map (
            O => \N__61568\,
            I => \N__61533\
        );

    \I__14182\ : Span12Mux_s11_h
    port map (
            O => \N__61565\,
            I => \N__61526\
        );

    \I__14181\ : Sp12to4
    port map (
            O => \N__61562\,
            I => \N__61526\
        );

    \I__14180\ : Sp12to4
    port map (
            O => \N__61559\,
            I => \N__61526\
        );

    \I__14179\ : Span4Mux_h
    port map (
            O => \N__61556\,
            I => \N__61521\
        );

    \I__14178\ : Span4Mux_v
    port map (
            O => \N__61553\,
            I => \N__61521\
        );

    \I__14177\ : Span12Mux_h
    port map (
            O => \N__61546\,
            I => \N__61516\
        );

    \I__14176\ : Sp12to4
    port map (
            O => \N__61541\,
            I => \N__61516\
        );

    \I__14175\ : Odrv4
    port map (
            O => \N__61536\,
            I => \aluOut_10\
        );

    \I__14174\ : Odrv4
    port map (
            O => \N__61533\,
            I => \aluOut_10\
        );

    \I__14173\ : Odrv12
    port map (
            O => \N__61526\,
            I => \aluOut_10\
        );

    \I__14172\ : Odrv4
    port map (
            O => \N__61521\,
            I => \aluOut_10\
        );

    \I__14171\ : Odrv12
    port map (
            O => \N__61516\,
            I => \aluOut_10\
        );

    \I__14170\ : InMux
    port map (
            O => \N__61505\,
            I => \N__61502\
        );

    \I__14169\ : LocalMux
    port map (
            O => \N__61502\,
            I => \N__61499\
        );

    \I__14168\ : Span4Mux_h
    port map (
            O => \N__61499\,
            I => \N__61496\
        );

    \I__14167\ : Span4Mux_h
    port map (
            O => \N__61496\,
            I => \N__61493\
        );

    \I__14166\ : Span4Mux_h
    port map (
            O => \N__61493\,
            I => \N__61489\
        );

    \I__14165\ : InMux
    port map (
            O => \N__61492\,
            I => \N__61486\
        );

    \I__14164\ : Span4Mux_v
    port map (
            O => \N__61489\,
            I => \N__61483\
        );

    \I__14163\ : LocalMux
    port map (
            O => \N__61486\,
            I => \ALU.addsub_10\
        );

    \I__14162\ : Odrv4
    port map (
            O => \N__61483\,
            I => \ALU.addsub_10\
        );

    \I__14161\ : InMux
    port map (
            O => \N__61478\,
            I => \ALU.addsub_cry_9\
        );

    \I__14160\ : InMux
    port map (
            O => \N__61475\,
            I => \N__61467\
        );

    \I__14159\ : InMux
    port map (
            O => \N__61474\,
            I => \N__61457\
        );

    \I__14158\ : InMux
    port map (
            O => \N__61473\,
            I => \N__61454\
        );

    \I__14157\ : InMux
    port map (
            O => \N__61472\,
            I => \N__61447\
        );

    \I__14156\ : InMux
    port map (
            O => \N__61471\,
            I => \N__61447\
        );

    \I__14155\ : InMux
    port map (
            O => \N__61470\,
            I => \N__61447\
        );

    \I__14154\ : LocalMux
    port map (
            O => \N__61467\,
            I => \N__61443\
        );

    \I__14153\ : InMux
    port map (
            O => \N__61466\,
            I => \N__61440\
        );

    \I__14152\ : InMux
    port map (
            O => \N__61465\,
            I => \N__61436\
        );

    \I__14151\ : InMux
    port map (
            O => \N__61464\,
            I => \N__61428\
        );

    \I__14150\ : InMux
    port map (
            O => \N__61463\,
            I => \N__61428\
        );

    \I__14149\ : InMux
    port map (
            O => \N__61462\,
            I => \N__61422\
        );

    \I__14148\ : InMux
    port map (
            O => \N__61461\,
            I => \N__61417\
        );

    \I__14147\ : InMux
    port map (
            O => \N__61460\,
            I => \N__61417\
        );

    \I__14146\ : LocalMux
    port map (
            O => \N__61457\,
            I => \N__61410\
        );

    \I__14145\ : LocalMux
    port map (
            O => \N__61454\,
            I => \N__61410\
        );

    \I__14144\ : LocalMux
    port map (
            O => \N__61447\,
            I => \N__61410\
        );

    \I__14143\ : InMux
    port map (
            O => \N__61446\,
            I => \N__61407\
        );

    \I__14142\ : Span4Mux_v
    port map (
            O => \N__61443\,
            I => \N__61404\
        );

    \I__14141\ : LocalMux
    port map (
            O => \N__61440\,
            I => \N__61401\
        );

    \I__14140\ : InMux
    port map (
            O => \N__61439\,
            I => \N__61398\
        );

    \I__14139\ : LocalMux
    port map (
            O => \N__61436\,
            I => \N__61395\
        );

    \I__14138\ : InMux
    port map (
            O => \N__61435\,
            I => \N__61390\
        );

    \I__14137\ : InMux
    port map (
            O => \N__61434\,
            I => \N__61390\
        );

    \I__14136\ : InMux
    port map (
            O => \N__61433\,
            I => \N__61387\
        );

    \I__14135\ : LocalMux
    port map (
            O => \N__61428\,
            I => \N__61384\
        );

    \I__14134\ : InMux
    port map (
            O => \N__61427\,
            I => \N__61381\
        );

    \I__14133\ : InMux
    port map (
            O => \N__61426\,
            I => \N__61378\
        );

    \I__14132\ : InMux
    port map (
            O => \N__61425\,
            I => \N__61375\
        );

    \I__14131\ : LocalMux
    port map (
            O => \N__61422\,
            I => \N__61372\
        );

    \I__14130\ : LocalMux
    port map (
            O => \N__61417\,
            I => \N__61365\
        );

    \I__14129\ : Span4Mux_v
    port map (
            O => \N__61410\,
            I => \N__61365\
        );

    \I__14128\ : LocalMux
    port map (
            O => \N__61407\,
            I => \N__61365\
        );

    \I__14127\ : Span4Mux_h
    port map (
            O => \N__61404\,
            I => \N__61353\
        );

    \I__14126\ : Span4Mux_v
    port map (
            O => \N__61401\,
            I => \N__61353\
        );

    \I__14125\ : LocalMux
    port map (
            O => \N__61398\,
            I => \N__61353\
        );

    \I__14124\ : Span4Mux_v
    port map (
            O => \N__61395\,
            I => \N__61353\
        );

    \I__14123\ : LocalMux
    port map (
            O => \N__61390\,
            I => \N__61353\
        );

    \I__14122\ : LocalMux
    port map (
            O => \N__61387\,
            I => \N__61350\
        );

    \I__14121\ : Span4Mux_h
    port map (
            O => \N__61384\,
            I => \N__61347\
        );

    \I__14120\ : LocalMux
    port map (
            O => \N__61381\,
            I => \N__61344\
        );

    \I__14119\ : LocalMux
    port map (
            O => \N__61378\,
            I => \N__61341\
        );

    \I__14118\ : LocalMux
    port map (
            O => \N__61375\,
            I => \N__61334\
        );

    \I__14117\ : Span4Mux_v
    port map (
            O => \N__61372\,
            I => \N__61334\
        );

    \I__14116\ : Span4Mux_h
    port map (
            O => \N__61365\,
            I => \N__61334\
        );

    \I__14115\ : InMux
    port map (
            O => \N__61364\,
            I => \N__61331\
        );

    \I__14114\ : Span4Mux_v
    port map (
            O => \N__61353\,
            I => \N__61328\
        );

    \I__14113\ : Span4Mux_v
    port map (
            O => \N__61350\,
            I => \N__61325\
        );

    \I__14112\ : Span4Mux_h
    port map (
            O => \N__61347\,
            I => \N__61322\
        );

    \I__14111\ : Span4Mux_h
    port map (
            O => \N__61344\,
            I => \N__61317\
        );

    \I__14110\ : Span4Mux_v
    port map (
            O => \N__61341\,
            I => \N__61317\
        );

    \I__14109\ : Span4Mux_h
    port map (
            O => \N__61334\,
            I => \N__61314\
        );

    \I__14108\ : LocalMux
    port map (
            O => \N__61331\,
            I => \N__61309\
        );

    \I__14107\ : Sp12to4
    port map (
            O => \N__61328\,
            I => \N__61309\
        );

    \I__14106\ : Odrv4
    port map (
            O => \N__61325\,
            I => \aluOut_11\
        );

    \I__14105\ : Odrv4
    port map (
            O => \N__61322\,
            I => \aluOut_11\
        );

    \I__14104\ : Odrv4
    port map (
            O => \N__61317\,
            I => \aluOut_11\
        );

    \I__14103\ : Odrv4
    port map (
            O => \N__61314\,
            I => \aluOut_11\
        );

    \I__14102\ : Odrv12
    port map (
            O => \N__61309\,
            I => \aluOut_11\
        );

    \I__14101\ : CascadeMux
    port map (
            O => \N__61298\,
            I => \N__61295\
        );

    \I__14100\ : InMux
    port map (
            O => \N__61295\,
            I => \N__61292\
        );

    \I__14099\ : LocalMux
    port map (
            O => \N__61292\,
            I => \N__61289\
        );

    \I__14098\ : Span4Mux_v
    port map (
            O => \N__61289\,
            I => \N__61286\
        );

    \I__14097\ : Sp12to4
    port map (
            O => \N__61286\,
            I => \N__61283\
        );

    \I__14096\ : Span12Mux_h
    port map (
            O => \N__61283\,
            I => \N__61280\
        );

    \I__14095\ : Odrv12
    port map (
            O => \N__61280\,
            I => \ALU.c_RNIRRB4IZ0Z_11\
        );

    \I__14094\ : InMux
    port map (
            O => \N__61277\,
            I => \N__61273\
        );

    \I__14093\ : InMux
    port map (
            O => \N__61276\,
            I => \N__61270\
        );

    \I__14092\ : LocalMux
    port map (
            O => \N__61273\,
            I => \N__61267\
        );

    \I__14091\ : LocalMux
    port map (
            O => \N__61270\,
            I => \N__61264\
        );

    \I__14090\ : Span4Mux_v
    port map (
            O => \N__61267\,
            I => \N__61261\
        );

    \I__14089\ : Span4Mux_h
    port map (
            O => \N__61264\,
            I => \N__61258\
        );

    \I__14088\ : Span4Mux_h
    port map (
            O => \N__61261\,
            I => \N__61255\
        );

    \I__14087\ : Span4Mux_h
    port map (
            O => \N__61258\,
            I => \N__61252\
        );

    \I__14086\ : Odrv4
    port map (
            O => \N__61255\,
            I => \ALU.addsub_11\
        );

    \I__14085\ : Odrv4
    port map (
            O => \N__61252\,
            I => \ALU.addsub_11\
        );

    \I__14084\ : InMux
    port map (
            O => \N__61247\,
            I => \ALU.addsub_cry_10\
        );

    \I__14083\ : InMux
    port map (
            O => \N__61244\,
            I => \N__61241\
        );

    \I__14082\ : LocalMux
    port map (
            O => \N__61241\,
            I => \N__61238\
        );

    \I__14081\ : Span4Mux_h
    port map (
            O => \N__61238\,
            I => \N__61235\
        );

    \I__14080\ : Span4Mux_v
    port map (
            O => \N__61235\,
            I => \N__61232\
        );

    \I__14079\ : Span4Mux_h
    port map (
            O => \N__61232\,
            I => \N__61229\
        );

    \I__14078\ : Odrv4
    port map (
            O => \N__61229\,
            I => \ALU.c_RNITVOEKZ0Z_12\
        );

    \I__14077\ : InMux
    port map (
            O => \N__61226\,
            I => \N__61221\
        );

    \I__14076\ : CascadeMux
    port map (
            O => \N__61225\,
            I => \N__61218\
        );

    \I__14075\ : CascadeMux
    port map (
            O => \N__61224\,
            I => \N__61213\
        );

    \I__14074\ : LocalMux
    port map (
            O => \N__61221\,
            I => \N__61207\
        );

    \I__14073\ : InMux
    port map (
            O => \N__61218\,
            I => \N__61204\
        );

    \I__14072\ : CascadeMux
    port map (
            O => \N__61217\,
            I => \N__61200\
        );

    \I__14071\ : CascadeMux
    port map (
            O => \N__61216\,
            I => \N__61196\
        );

    \I__14070\ : InMux
    port map (
            O => \N__61213\,
            I => \N__61190\
        );

    \I__14069\ : InMux
    port map (
            O => \N__61212\,
            I => \N__61187\
        );

    \I__14068\ : InMux
    port map (
            O => \N__61211\,
            I => \N__61184\
        );

    \I__14067\ : CascadeMux
    port map (
            O => \N__61210\,
            I => \N__61181\
        );

    \I__14066\ : Span4Mux_v
    port map (
            O => \N__61207\,
            I => \N__61176\
        );

    \I__14065\ : LocalMux
    port map (
            O => \N__61204\,
            I => \N__61176\
        );

    \I__14064\ : InMux
    port map (
            O => \N__61203\,
            I => \N__61171\
        );

    \I__14063\ : InMux
    port map (
            O => \N__61200\,
            I => \N__61171\
        );

    \I__14062\ : InMux
    port map (
            O => \N__61199\,
            I => \N__61167\
        );

    \I__14061\ : InMux
    port map (
            O => \N__61196\,
            I => \N__61164\
        );

    \I__14060\ : InMux
    port map (
            O => \N__61195\,
            I => \N__61161\
        );

    \I__14059\ : CascadeMux
    port map (
            O => \N__61194\,
            I => \N__61158\
        );

    \I__14058\ : InMux
    port map (
            O => \N__61193\,
            I => \N__61153\
        );

    \I__14057\ : LocalMux
    port map (
            O => \N__61190\,
            I => \N__61148\
        );

    \I__14056\ : LocalMux
    port map (
            O => \N__61187\,
            I => \N__61143\
        );

    \I__14055\ : LocalMux
    port map (
            O => \N__61184\,
            I => \N__61143\
        );

    \I__14054\ : InMux
    port map (
            O => \N__61181\,
            I => \N__61140\
        );

    \I__14053\ : Span4Mux_h
    port map (
            O => \N__61176\,
            I => \N__61135\
        );

    \I__14052\ : LocalMux
    port map (
            O => \N__61171\,
            I => \N__61135\
        );

    \I__14051\ : InMux
    port map (
            O => \N__61170\,
            I => \N__61132\
        );

    \I__14050\ : LocalMux
    port map (
            O => \N__61167\,
            I => \N__61129\
        );

    \I__14049\ : LocalMux
    port map (
            O => \N__61164\,
            I => \N__61126\
        );

    \I__14048\ : LocalMux
    port map (
            O => \N__61161\,
            I => \N__61123\
        );

    \I__14047\ : InMux
    port map (
            O => \N__61158\,
            I => \N__61120\
        );

    \I__14046\ : InMux
    port map (
            O => \N__61157\,
            I => \N__61115\
        );

    \I__14045\ : InMux
    port map (
            O => \N__61156\,
            I => \N__61115\
        );

    \I__14044\ : LocalMux
    port map (
            O => \N__61153\,
            I => \N__61112\
        );

    \I__14043\ : InMux
    port map (
            O => \N__61152\,
            I => \N__61107\
        );

    \I__14042\ : InMux
    port map (
            O => \N__61151\,
            I => \N__61107\
        );

    \I__14041\ : Span4Mux_v
    port map (
            O => \N__61148\,
            I => \N__61104\
        );

    \I__14040\ : Span4Mux_v
    port map (
            O => \N__61143\,
            I => \N__61101\
        );

    \I__14039\ : LocalMux
    port map (
            O => \N__61140\,
            I => \N__61094\
        );

    \I__14038\ : Span4Mux_h
    port map (
            O => \N__61135\,
            I => \N__61094\
        );

    \I__14037\ : LocalMux
    port map (
            O => \N__61132\,
            I => \N__61094\
        );

    \I__14036\ : Span4Mux_h
    port map (
            O => \N__61129\,
            I => \N__61091\
        );

    \I__14035\ : Span4Mux_v
    port map (
            O => \N__61126\,
            I => \N__61082\
        );

    \I__14034\ : Span4Mux_v
    port map (
            O => \N__61123\,
            I => \N__61082\
        );

    \I__14033\ : LocalMux
    port map (
            O => \N__61120\,
            I => \N__61082\
        );

    \I__14032\ : LocalMux
    port map (
            O => \N__61115\,
            I => \N__61082\
        );

    \I__14031\ : Span4Mux_v
    port map (
            O => \N__61112\,
            I => \N__61079\
        );

    \I__14030\ : LocalMux
    port map (
            O => \N__61107\,
            I => \N__61076\
        );

    \I__14029\ : Span4Mux_h
    port map (
            O => \N__61104\,
            I => \N__61071\
        );

    \I__14028\ : Span4Mux_v
    port map (
            O => \N__61101\,
            I => \N__61071\
        );

    \I__14027\ : Span4Mux_v
    port map (
            O => \N__61094\,
            I => \N__61068\
        );

    \I__14026\ : Span4Mux_v
    port map (
            O => \N__61091\,
            I => \N__61063\
        );

    \I__14025\ : Span4Mux_h
    port map (
            O => \N__61082\,
            I => \N__61063\
        );

    \I__14024\ : Span4Mux_h
    port map (
            O => \N__61079\,
            I => \N__61058\
        );

    \I__14023\ : Span4Mux_h
    port map (
            O => \N__61076\,
            I => \N__61058\
        );

    \I__14022\ : Span4Mux_h
    port map (
            O => \N__61071\,
            I => \N__61053\
        );

    \I__14021\ : Span4Mux_v
    port map (
            O => \N__61068\,
            I => \N__61053\
        );

    \I__14020\ : Span4Mux_v
    port map (
            O => \N__61063\,
            I => \N__61050\
        );

    \I__14019\ : Odrv4
    port map (
            O => \N__61058\,
            I => \aluOut_12\
        );

    \I__14018\ : Odrv4
    port map (
            O => \N__61053\,
            I => \aluOut_12\
        );

    \I__14017\ : Odrv4
    port map (
            O => \N__61050\,
            I => \aluOut_12\
        );

    \I__14016\ : InMux
    port map (
            O => \N__61043\,
            I => \N__61037\
        );

    \I__14015\ : InMux
    port map (
            O => \N__61042\,
            I => \N__61037\
        );

    \I__14014\ : LocalMux
    port map (
            O => \N__61037\,
            I => \N__61034\
        );

    \I__14013\ : Span4Mux_v
    port map (
            O => \N__61034\,
            I => \N__61031\
        );

    \I__14012\ : Odrv4
    port map (
            O => \N__61031\,
            I => \ALU.addsub_12\
        );

    \I__14011\ : InMux
    port map (
            O => \N__61028\,
            I => \ALU.addsub_cry_11\
        );

    \I__14010\ : InMux
    port map (
            O => \N__61025\,
            I => \N__61022\
        );

    \I__14009\ : LocalMux
    port map (
            O => \N__61022\,
            I => \ALU.c_RNIVHVMKZ0Z_13\
        );

    \I__14008\ : CascadeMux
    port map (
            O => \N__61019\,
            I => \N__61015\
        );

    \I__14007\ : InMux
    port map (
            O => \N__61018\,
            I => \N__61005\
        );

    \I__14006\ : InMux
    port map (
            O => \N__61015\,
            I => \N__61002\
        );

    \I__14005\ : InMux
    port map (
            O => \N__61014\,
            I => \N__60999\
        );

    \I__14004\ : CascadeMux
    port map (
            O => \N__61013\,
            I => \N__60996\
        );

    \I__14003\ : InMux
    port map (
            O => \N__61012\,
            I => \N__60991\
        );

    \I__14002\ : InMux
    port map (
            O => \N__61011\,
            I => \N__60987\
        );

    \I__14001\ : InMux
    port map (
            O => \N__61010\,
            I => \N__60984\
        );

    \I__14000\ : InMux
    port map (
            O => \N__61009\,
            I => \N__60979\
        );

    \I__13999\ : InMux
    port map (
            O => \N__61008\,
            I => \N__60979\
        );

    \I__13998\ : LocalMux
    port map (
            O => \N__61005\,
            I => \N__60972\
        );

    \I__13997\ : LocalMux
    port map (
            O => \N__61002\,
            I => \N__60972\
        );

    \I__13996\ : LocalMux
    port map (
            O => \N__60999\,
            I => \N__60972\
        );

    \I__13995\ : InMux
    port map (
            O => \N__60996\,
            I => \N__60969\
        );

    \I__13994\ : InMux
    port map (
            O => \N__60995\,
            I => \N__60966\
        );

    \I__13993\ : InMux
    port map (
            O => \N__60994\,
            I => \N__60961\
        );

    \I__13992\ : LocalMux
    port map (
            O => \N__60991\,
            I => \N__60958\
        );

    \I__13991\ : InMux
    port map (
            O => \N__60990\,
            I => \N__60955\
        );

    \I__13990\ : LocalMux
    port map (
            O => \N__60987\,
            I => \N__60950\
        );

    \I__13989\ : LocalMux
    port map (
            O => \N__60984\,
            I => \N__60947\
        );

    \I__13988\ : LocalMux
    port map (
            O => \N__60979\,
            I => \N__60944\
        );

    \I__13987\ : Span4Mux_h
    port map (
            O => \N__60972\,
            I => \N__60941\
        );

    \I__13986\ : LocalMux
    port map (
            O => \N__60969\,
            I => \N__60933\
        );

    \I__13985\ : LocalMux
    port map (
            O => \N__60966\,
            I => \N__60933\
        );

    \I__13984\ : InMux
    port map (
            O => \N__60965\,
            I => \N__60928\
        );

    \I__13983\ : InMux
    port map (
            O => \N__60964\,
            I => \N__60928\
        );

    \I__13982\ : LocalMux
    port map (
            O => \N__60961\,
            I => \N__60925\
        );

    \I__13981\ : Span4Mux_v
    port map (
            O => \N__60958\,
            I => \N__60920\
        );

    \I__13980\ : LocalMux
    port map (
            O => \N__60955\,
            I => \N__60920\
        );

    \I__13979\ : InMux
    port map (
            O => \N__60954\,
            I => \N__60917\
        );

    \I__13978\ : InMux
    port map (
            O => \N__60953\,
            I => \N__60914\
        );

    \I__13977\ : Span4Mux_v
    port map (
            O => \N__60950\,
            I => \N__60911\
        );

    \I__13976\ : Span4Mux_v
    port map (
            O => \N__60947\,
            I => \N__60906\
        );

    \I__13975\ : Span4Mux_v
    port map (
            O => \N__60944\,
            I => \N__60906\
        );

    \I__13974\ : Span4Mux_v
    port map (
            O => \N__60941\,
            I => \N__60903\
        );

    \I__13973\ : InMux
    port map (
            O => \N__60940\,
            I => \N__60896\
        );

    \I__13972\ : InMux
    port map (
            O => \N__60939\,
            I => \N__60896\
        );

    \I__13971\ : InMux
    port map (
            O => \N__60938\,
            I => \N__60896\
        );

    \I__13970\ : Span4Mux_v
    port map (
            O => \N__60933\,
            I => \N__60893\
        );

    \I__13969\ : LocalMux
    port map (
            O => \N__60928\,
            I => \N__60890\
        );

    \I__13968\ : Span4Mux_v
    port map (
            O => \N__60925\,
            I => \N__60887\
        );

    \I__13967\ : Span4Mux_v
    port map (
            O => \N__60920\,
            I => \N__60884\
        );

    \I__13966\ : LocalMux
    port map (
            O => \N__60917\,
            I => \N__60879\
        );

    \I__13965\ : LocalMux
    port map (
            O => \N__60914\,
            I => \N__60879\
        );

    \I__13964\ : Sp12to4
    port map (
            O => \N__60911\,
            I => \N__60870\
        );

    \I__13963\ : Sp12to4
    port map (
            O => \N__60906\,
            I => \N__60870\
        );

    \I__13962\ : Sp12to4
    port map (
            O => \N__60903\,
            I => \N__60870\
        );

    \I__13961\ : LocalMux
    port map (
            O => \N__60896\,
            I => \N__60870\
        );

    \I__13960\ : Span4Mux_v
    port map (
            O => \N__60893\,
            I => \N__60867\
        );

    \I__13959\ : Span4Mux_v
    port map (
            O => \N__60890\,
            I => \N__60864\
        );

    \I__13958\ : Span4Mux_v
    port map (
            O => \N__60887\,
            I => \N__60861\
        );

    \I__13957\ : Span4Mux_v
    port map (
            O => \N__60884\,
            I => \N__60858\
        );

    \I__13956\ : Sp12to4
    port map (
            O => \N__60879\,
            I => \N__60853\
        );

    \I__13955\ : Span12Mux_h
    port map (
            O => \N__60870\,
            I => \N__60853\
        );

    \I__13954\ : Span4Mux_h
    port map (
            O => \N__60867\,
            I => \N__60848\
        );

    \I__13953\ : Span4Mux_v
    port map (
            O => \N__60864\,
            I => \N__60848\
        );

    \I__13952\ : Odrv4
    port map (
            O => \N__60861\,
            I => \aluOut_13\
        );

    \I__13951\ : Odrv4
    port map (
            O => \N__60858\,
            I => \aluOut_13\
        );

    \I__13950\ : Odrv12
    port map (
            O => \N__60853\,
            I => \aluOut_13\
        );

    \I__13949\ : Odrv4
    port map (
            O => \N__60848\,
            I => \aluOut_13\
        );

    \I__13948\ : InMux
    port map (
            O => \N__60839\,
            I => \N__60836\
        );

    \I__13947\ : LocalMux
    port map (
            O => \N__60836\,
            I => \N__60832\
        );

    \I__13946\ : InMux
    port map (
            O => \N__60835\,
            I => \N__60829\
        );

    \I__13945\ : Span4Mux_h
    port map (
            O => \N__60832\,
            I => \N__60826\
        );

    \I__13944\ : LocalMux
    port map (
            O => \N__60829\,
            I => \N__60823\
        );

    \I__13943\ : Odrv4
    port map (
            O => \N__60826\,
            I => \ALU.addsub_13\
        );

    \I__13942\ : Odrv12
    port map (
            O => \N__60823\,
            I => \ALU.addsub_13\
        );

    \I__13941\ : CascadeMux
    port map (
            O => \N__60818\,
            I => \N__60815\
        );

    \I__13940\ : InMux
    port map (
            O => \N__60815\,
            I => \N__60809\
        );

    \I__13939\ : CascadeMux
    port map (
            O => \N__60814\,
            I => \N__60806\
        );

    \I__13938\ : InMux
    port map (
            O => \N__60813\,
            I => \N__60802\
        );

    \I__13937\ : CascadeMux
    port map (
            O => \N__60812\,
            I => \N__60799\
        );

    \I__13936\ : LocalMux
    port map (
            O => \N__60809\,
            I => \N__60796\
        );

    \I__13935\ : InMux
    port map (
            O => \N__60806\,
            I => \N__60793\
        );

    \I__13934\ : CascadeMux
    port map (
            O => \N__60805\,
            I => \N__60790\
        );

    \I__13933\ : LocalMux
    port map (
            O => \N__60802\,
            I => \N__60787\
        );

    \I__13932\ : InMux
    port map (
            O => \N__60799\,
            I => \N__60784\
        );

    \I__13931\ : Sp12to4
    port map (
            O => \N__60796\,
            I => \N__60781\
        );

    \I__13930\ : LocalMux
    port map (
            O => \N__60793\,
            I => \N__60777\
        );

    \I__13929\ : InMux
    port map (
            O => \N__60790\,
            I => \N__60774\
        );

    \I__13928\ : Span4Mux_v
    port map (
            O => \N__60787\,
            I => \N__60769\
        );

    \I__13927\ : LocalMux
    port map (
            O => \N__60784\,
            I => \N__60769\
        );

    \I__13926\ : Span12Mux_v
    port map (
            O => \N__60781\,
            I => \N__60766\
        );

    \I__13925\ : InMux
    port map (
            O => \N__60780\,
            I => \N__60763\
        );

    \I__13924\ : Span4Mux_v
    port map (
            O => \N__60777\,
            I => \N__60760\
        );

    \I__13923\ : LocalMux
    port map (
            O => \N__60774\,
            I => \N__60755\
        );

    \I__13922\ : Span4Mux_h
    port map (
            O => \N__60769\,
            I => \N__60755\
        );

    \I__13921\ : Span12Mux_h
    port map (
            O => \N__60766\,
            I => \N__60752\
        );

    \I__13920\ : LocalMux
    port map (
            O => \N__60763\,
            I => \CONTROL.addrstackptrZ0Z_4\
        );

    \I__13919\ : Odrv4
    port map (
            O => \N__60760\,
            I => \CONTROL.addrstackptrZ0Z_4\
        );

    \I__13918\ : Odrv4
    port map (
            O => \N__60755\,
            I => \CONTROL.addrstackptrZ0Z_4\
        );

    \I__13917\ : Odrv12
    port map (
            O => \N__60752\,
            I => \CONTROL.addrstackptrZ0Z_4\
        );

    \I__13916\ : CascadeMux
    port map (
            O => \N__60743\,
            I => \N__60740\
        );

    \I__13915\ : InMux
    port map (
            O => \N__60740\,
            I => \N__60737\
        );

    \I__13914\ : LocalMux
    port map (
            O => \N__60737\,
            I => \N__60731\
        );

    \I__13913\ : InMux
    port map (
            O => \N__60736\,
            I => \N__60727\
        );

    \I__13912\ : CascadeMux
    port map (
            O => \N__60735\,
            I => \N__60724\
        );

    \I__13911\ : CascadeMux
    port map (
            O => \N__60734\,
            I => \N__60720\
        );

    \I__13910\ : Span4Mux_v
    port map (
            O => \N__60731\,
            I => \N__60717\
        );

    \I__13909\ : InMux
    port map (
            O => \N__60730\,
            I => \N__60714\
        );

    \I__13908\ : LocalMux
    port map (
            O => \N__60727\,
            I => \N__60711\
        );

    \I__13907\ : InMux
    port map (
            O => \N__60724\,
            I => \N__60708\
        );

    \I__13906\ : InMux
    port map (
            O => \N__60723\,
            I => \N__60705\
        );

    \I__13905\ : InMux
    port map (
            O => \N__60720\,
            I => \N__60702\
        );

    \I__13904\ : Span4Mux_h
    port map (
            O => \N__60717\,
            I => \N__60696\
        );

    \I__13903\ : LocalMux
    port map (
            O => \N__60714\,
            I => \N__60696\
        );

    \I__13902\ : Span4Mux_h
    port map (
            O => \N__60711\,
            I => \N__60693\
        );

    \I__13901\ : LocalMux
    port map (
            O => \N__60708\,
            I => \N__60686\
        );

    \I__13900\ : LocalMux
    port map (
            O => \N__60705\,
            I => \N__60686\
        );

    \I__13899\ : LocalMux
    port map (
            O => \N__60702\,
            I => \N__60686\
        );

    \I__13898\ : CascadeMux
    port map (
            O => \N__60701\,
            I => \N__60683\
        );

    \I__13897\ : Sp12to4
    port map (
            O => \N__60696\,
            I => \N__60679\
        );

    \I__13896\ : Sp12to4
    port map (
            O => \N__60693\,
            I => \N__60676\
        );

    \I__13895\ : Span4Mux_v
    port map (
            O => \N__60686\,
            I => \N__60673\
        );

    \I__13894\ : InMux
    port map (
            O => \N__60683\,
            I => \N__60668\
        );

    \I__13893\ : InMux
    port map (
            O => \N__60682\,
            I => \N__60668\
        );

    \I__13892\ : Span12Mux_h
    port map (
            O => \N__60679\,
            I => \N__60663\
        );

    \I__13891\ : Span12Mux_v
    port map (
            O => \N__60676\,
            I => \N__60663\
        );

    \I__13890\ : Sp12to4
    port map (
            O => \N__60673\,
            I => \N__60660\
        );

    \I__13889\ : LocalMux
    port map (
            O => \N__60668\,
            I => \CONTROL.addrstackptrZ0Z_2\
        );

    \I__13888\ : Odrv12
    port map (
            O => \N__60663\,
            I => \CONTROL.addrstackptrZ0Z_2\
        );

    \I__13887\ : Odrv12
    port map (
            O => \N__60660\,
            I => \CONTROL.addrstackptrZ0Z_2\
        );

    \I__13886\ : InMux
    port map (
            O => \N__60653\,
            I => \N__60650\
        );

    \I__13885\ : LocalMux
    port map (
            O => \N__60650\,
            I => \N__60647\
        );

    \I__13884\ : Span4Mux_v
    port map (
            O => \N__60647\,
            I => \N__60644\
        );

    \I__13883\ : Span4Mux_h
    port map (
            O => \N__60644\,
            I => \N__60641\
        );

    \I__13882\ : Span4Mux_h
    port map (
            O => \N__60641\,
            I => \N__60638\
        );

    \I__13881\ : Span4Mux_v
    port map (
            O => \N__60638\,
            I => \N__60635\
        );

    \I__13880\ : Span4Mux_v
    port map (
            O => \N__60635\,
            I => \N__60632\
        );

    \I__13879\ : Odrv4
    port map (
            O => \N__60632\,
            I => \CONTROL.g1_1_3\
        );

    \I__13878\ : CascadeMux
    port map (
            O => \N__60629\,
            I => \N__60621\
        );

    \I__13877\ : CascadeMux
    port map (
            O => \N__60628\,
            I => \N__60618\
        );

    \I__13876\ : CascadeMux
    port map (
            O => \N__60627\,
            I => \N__60613\
        );

    \I__13875\ : CascadeMux
    port map (
            O => \N__60626\,
            I => \N__60610\
        );

    \I__13874\ : InMux
    port map (
            O => \N__60625\,
            I => \N__60606\
        );

    \I__13873\ : InMux
    port map (
            O => \N__60624\,
            I => \N__60603\
        );

    \I__13872\ : InMux
    port map (
            O => \N__60621\,
            I => \N__60599\
        );

    \I__13871\ : InMux
    port map (
            O => \N__60618\,
            I => \N__60595\
        );

    \I__13870\ : InMux
    port map (
            O => \N__60617\,
            I => \N__60590\
        );

    \I__13869\ : InMux
    port map (
            O => \N__60616\,
            I => \N__60586\
        );

    \I__13868\ : InMux
    port map (
            O => \N__60613\,
            I => \N__60580\
        );

    \I__13867\ : InMux
    port map (
            O => \N__60610\,
            I => \N__60580\
        );

    \I__13866\ : CascadeMux
    port map (
            O => \N__60609\,
            I => \N__60576\
        );

    \I__13865\ : LocalMux
    port map (
            O => \N__60606\,
            I => \N__60569\
        );

    \I__13864\ : LocalMux
    port map (
            O => \N__60603\,
            I => \N__60563\
        );

    \I__13863\ : InMux
    port map (
            O => \N__60602\,
            I => \N__60560\
        );

    \I__13862\ : LocalMux
    port map (
            O => \N__60599\,
            I => \N__60557\
        );

    \I__13861\ : InMux
    port map (
            O => \N__60598\,
            I => \N__60554\
        );

    \I__13860\ : LocalMux
    port map (
            O => \N__60595\,
            I => \N__60551\
        );

    \I__13859\ : InMux
    port map (
            O => \N__60594\,
            I => \N__60546\
        );

    \I__13858\ : InMux
    port map (
            O => \N__60593\,
            I => \N__60546\
        );

    \I__13857\ : LocalMux
    port map (
            O => \N__60590\,
            I => \N__60536\
        );

    \I__13856\ : InMux
    port map (
            O => \N__60589\,
            I => \N__60533\
        );

    \I__13855\ : LocalMux
    port map (
            O => \N__60586\,
            I => \N__60530\
        );

    \I__13854\ : InMux
    port map (
            O => \N__60585\,
            I => \N__60527\
        );

    \I__13853\ : LocalMux
    port map (
            O => \N__60580\,
            I => \N__60524\
        );

    \I__13852\ : InMux
    port map (
            O => \N__60579\,
            I => \N__60521\
        );

    \I__13851\ : InMux
    port map (
            O => \N__60576\,
            I => \N__60518\
        );

    \I__13850\ : InMux
    port map (
            O => \N__60575\,
            I => \N__60513\
        );

    \I__13849\ : InMux
    port map (
            O => \N__60574\,
            I => \N__60513\
        );

    \I__13848\ : InMux
    port map (
            O => \N__60573\,
            I => \N__60508\
        );

    \I__13847\ : InMux
    port map (
            O => \N__60572\,
            I => \N__60508\
        );

    \I__13846\ : Span4Mux_v
    port map (
            O => \N__60569\,
            I => \N__60505\
        );

    \I__13845\ : InMux
    port map (
            O => \N__60568\,
            I => \N__60500\
        );

    \I__13844\ : InMux
    port map (
            O => \N__60567\,
            I => \N__60500\
        );

    \I__13843\ : InMux
    port map (
            O => \N__60566\,
            I => \N__60497\
        );

    \I__13842\ : Span4Mux_v
    port map (
            O => \N__60563\,
            I => \N__60492\
        );

    \I__13841\ : LocalMux
    port map (
            O => \N__60560\,
            I => \N__60492\
        );

    \I__13840\ : Span4Mux_v
    port map (
            O => \N__60557\,
            I => \N__60485\
        );

    \I__13839\ : LocalMux
    port map (
            O => \N__60554\,
            I => \N__60485\
        );

    \I__13838\ : Span4Mux_h
    port map (
            O => \N__60551\,
            I => \N__60485\
        );

    \I__13837\ : LocalMux
    port map (
            O => \N__60546\,
            I => \N__60482\
        );

    \I__13836\ : InMux
    port map (
            O => \N__60545\,
            I => \N__60471\
        );

    \I__13835\ : InMux
    port map (
            O => \N__60544\,
            I => \N__60471\
        );

    \I__13834\ : InMux
    port map (
            O => \N__60543\,
            I => \N__60471\
        );

    \I__13833\ : InMux
    port map (
            O => \N__60542\,
            I => \N__60471\
        );

    \I__13832\ : InMux
    port map (
            O => \N__60541\,
            I => \N__60471\
        );

    \I__13831\ : InMux
    port map (
            O => \N__60540\,
            I => \N__60466\
        );

    \I__13830\ : InMux
    port map (
            O => \N__60539\,
            I => \N__60466\
        );

    \I__13829\ : Span4Mux_h
    port map (
            O => \N__60536\,
            I => \N__60461\
        );

    \I__13828\ : LocalMux
    port map (
            O => \N__60533\,
            I => \N__60461\
        );

    \I__13827\ : Span4Mux_v
    port map (
            O => \N__60530\,
            I => \N__60454\
        );

    \I__13826\ : LocalMux
    port map (
            O => \N__60527\,
            I => \N__60454\
        );

    \I__13825\ : Span4Mux_v
    port map (
            O => \N__60524\,
            I => \N__60454\
        );

    \I__13824\ : LocalMux
    port map (
            O => \N__60521\,
            I => \N__60451\
        );

    \I__13823\ : LocalMux
    port map (
            O => \N__60518\,
            I => \N__60448\
        );

    \I__13822\ : LocalMux
    port map (
            O => \N__60513\,
            I => \N__60445\
        );

    \I__13821\ : LocalMux
    port map (
            O => \N__60508\,
            I => \N__60438\
        );

    \I__13820\ : Span4Mux_h
    port map (
            O => \N__60505\,
            I => \N__60438\
        );

    \I__13819\ : LocalMux
    port map (
            O => \N__60500\,
            I => \N__60438\
        );

    \I__13818\ : LocalMux
    port map (
            O => \N__60497\,
            I => \N__60433\
        );

    \I__13817\ : Span4Mux_v
    port map (
            O => \N__60492\,
            I => \N__60433\
        );

    \I__13816\ : Span4Mux_v
    port map (
            O => \N__60485\,
            I => \N__60430\
        );

    \I__13815\ : Span4Mux_v
    port map (
            O => \N__60482\,
            I => \N__60427\
        );

    \I__13814\ : LocalMux
    port map (
            O => \N__60471\,
            I => \N__60418\
        );

    \I__13813\ : LocalMux
    port map (
            O => \N__60466\,
            I => \N__60418\
        );

    \I__13812\ : Span4Mux_h
    port map (
            O => \N__60461\,
            I => \N__60418\
        );

    \I__13811\ : Span4Mux_h
    port map (
            O => \N__60454\,
            I => \N__60418\
        );

    \I__13810\ : Span12Mux_v
    port map (
            O => \N__60451\,
            I => \N__60415\
        );

    \I__13809\ : Span4Mux_v
    port map (
            O => \N__60448\,
            I => \N__60412\
        );

    \I__13808\ : Span4Mux_v
    port map (
            O => \N__60445\,
            I => \N__60407\
        );

    \I__13807\ : Span4Mux_h
    port map (
            O => \N__60438\,
            I => \N__60407\
        );

    \I__13806\ : Span4Mux_v
    port map (
            O => \N__60433\,
            I => \N__60402\
        );

    \I__13805\ : Span4Mux_v
    port map (
            O => \N__60430\,
            I => \N__60402\
        );

    \I__13804\ : Span4Mux_h
    port map (
            O => \N__60427\,
            I => \N__60397\
        );

    \I__13803\ : Span4Mux_v
    port map (
            O => \N__60418\,
            I => \N__60397\
        );

    \I__13802\ : Odrv12
    port map (
            O => \N__60415\,
            I => \aluOut_0\
        );

    \I__13801\ : Odrv4
    port map (
            O => \N__60412\,
            I => \aluOut_0\
        );

    \I__13800\ : Odrv4
    port map (
            O => \N__60407\,
            I => \aluOut_0\
        );

    \I__13799\ : Odrv4
    port map (
            O => \N__60402\,
            I => \aluOut_0\
        );

    \I__13798\ : Odrv4
    port map (
            O => \N__60397\,
            I => \aluOut_0\
        );

    \I__13797\ : CascadeMux
    port map (
            O => \N__60386\,
            I => \N__60383\
        );

    \I__13796\ : InMux
    port map (
            O => \N__60383\,
            I => \N__60380\
        );

    \I__13795\ : LocalMux
    port map (
            O => \N__60380\,
            I => \N__60377\
        );

    \I__13794\ : Span4Mux_h
    port map (
            O => \N__60377\,
            I => \N__60374\
        );

    \I__13793\ : Span4Mux_h
    port map (
            O => \N__60374\,
            I => \N__60371\
        );

    \I__13792\ : Span4Mux_v
    port map (
            O => \N__60371\,
            I => \N__60368\
        );

    \I__13791\ : Odrv4
    port map (
            O => \N__60368\,
            I => \ALU.d_RNI27KBDZ0Z_0\
        );

    \I__13790\ : InMux
    port map (
            O => \N__60365\,
            I => \N__60362\
        );

    \I__13789\ : LocalMux
    port map (
            O => \N__60362\,
            I => \N__60359\
        );

    \I__13788\ : Span12Mux_h
    port map (
            O => \N__60359\,
            I => \N__60355\
        );

    \I__13787\ : InMux
    port map (
            O => \N__60358\,
            I => \N__60352\
        );

    \I__13786\ : Odrv12
    port map (
            O => \N__60355\,
            I => \ALU.addsub_0\
        );

    \I__13785\ : LocalMux
    port map (
            O => \N__60352\,
            I => \ALU.addsub_0\
        );

    \I__13784\ : InMux
    port map (
            O => \N__60347\,
            I => \ALU.addsub_cry_0_c_THRU_CO\
        );

    \I__13783\ : CascadeMux
    port map (
            O => \N__60344\,
            I => \N__60341\
        );

    \I__13782\ : InMux
    port map (
            O => \N__60341\,
            I => \N__60338\
        );

    \I__13781\ : LocalMux
    port map (
            O => \N__60338\,
            I => \N__60335\
        );

    \I__13780\ : Span4Mux_v
    port map (
            O => \N__60335\,
            I => \N__60332\
        );

    \I__13779\ : Span4Mux_h
    port map (
            O => \N__60332\,
            I => \N__60329\
        );

    \I__13778\ : Odrv4
    port map (
            O => \N__60329\,
            I => \ALU.d_RNIIEOKOZ0Z_1\
        );

    \I__13777\ : InMux
    port map (
            O => \N__60326\,
            I => \N__60323\
        );

    \I__13776\ : LocalMux
    port map (
            O => \N__60323\,
            I => \N__60320\
        );

    \I__13775\ : Span12Mux_v
    port map (
            O => \N__60320\,
            I => \N__60316\
        );

    \I__13774\ : InMux
    port map (
            O => \N__60319\,
            I => \N__60313\
        );

    \I__13773\ : Odrv12
    port map (
            O => \N__60316\,
            I => \ALU.addsub_1\
        );

    \I__13772\ : LocalMux
    port map (
            O => \N__60313\,
            I => \ALU.addsub_1\
        );

    \I__13771\ : InMux
    port map (
            O => \N__60308\,
            I => \ALU.addsub_cry_0\
        );

    \I__13770\ : CascadeMux
    port map (
            O => \N__60305\,
            I => \N__60302\
        );

    \I__13769\ : InMux
    port map (
            O => \N__60302\,
            I => \N__60299\
        );

    \I__13768\ : LocalMux
    port map (
            O => \N__60299\,
            I => \N__60296\
        );

    \I__13767\ : Span12Mux_h
    port map (
            O => \N__60296\,
            I => \N__60293\
        );

    \I__13766\ : Odrv12
    port map (
            O => \N__60293\,
            I => \ALU.d_RNIN178LZ0Z_2\
        );

    \I__13765\ : InMux
    port map (
            O => \N__60290\,
            I => \N__60287\
        );

    \I__13764\ : LocalMux
    port map (
            O => \N__60287\,
            I => \N__60284\
        );

    \I__13763\ : Span4Mux_h
    port map (
            O => \N__60284\,
            I => \N__60281\
        );

    \I__13762\ : Span4Mux_h
    port map (
            O => \N__60281\,
            I => \N__60277\
        );

    \I__13761\ : InMux
    port map (
            O => \N__60280\,
            I => \N__60274\
        );

    \I__13760\ : Odrv4
    port map (
            O => \N__60277\,
            I => \ALU.addsub_2\
        );

    \I__13759\ : LocalMux
    port map (
            O => \N__60274\,
            I => \ALU.addsub_2\
        );

    \I__13758\ : InMux
    port map (
            O => \N__60269\,
            I => \ALU.addsub_cry_1\
        );

    \I__13757\ : InMux
    port map (
            O => \N__60266\,
            I => \N__60257\
        );

    \I__13756\ : InMux
    port map (
            O => \N__60265\,
            I => \N__60254\
        );

    \I__13755\ : CascadeMux
    port map (
            O => \N__60264\,
            I => \N__60251\
        );

    \I__13754\ : CascadeMux
    port map (
            O => \N__60263\,
            I => \N__60248\
        );

    \I__13753\ : CascadeMux
    port map (
            O => \N__60262\,
            I => \N__60242\
        );

    \I__13752\ : InMux
    port map (
            O => \N__60261\,
            I => \N__60238\
        );

    \I__13751\ : InMux
    port map (
            O => \N__60260\,
            I => \N__60233\
        );

    \I__13750\ : LocalMux
    port map (
            O => \N__60257\,
            I => \N__60228\
        );

    \I__13749\ : LocalMux
    port map (
            O => \N__60254\,
            I => \N__60228\
        );

    \I__13748\ : InMux
    port map (
            O => \N__60251\,
            I => \N__60224\
        );

    \I__13747\ : InMux
    port map (
            O => \N__60248\,
            I => \N__60221\
        );

    \I__13746\ : CascadeMux
    port map (
            O => \N__60247\,
            I => \N__60215\
        );

    \I__13745\ : InMux
    port map (
            O => \N__60246\,
            I => \N__60210\
        );

    \I__13744\ : InMux
    port map (
            O => \N__60245\,
            I => \N__60202\
        );

    \I__13743\ : InMux
    port map (
            O => \N__60242\,
            I => \N__60199\
        );

    \I__13742\ : CascadeMux
    port map (
            O => \N__60241\,
            I => \N__60193\
        );

    \I__13741\ : LocalMux
    port map (
            O => \N__60238\,
            I => \N__60184\
        );

    \I__13740\ : InMux
    port map (
            O => \N__60237\,
            I => \N__60181\
        );

    \I__13739\ : InMux
    port map (
            O => \N__60236\,
            I => \N__60178\
        );

    \I__13738\ : LocalMux
    port map (
            O => \N__60233\,
            I => \N__60173\
        );

    \I__13737\ : Span4Mux_v
    port map (
            O => \N__60228\,
            I => \N__60173\
        );

    \I__13736\ : InMux
    port map (
            O => \N__60227\,
            I => \N__60170\
        );

    \I__13735\ : LocalMux
    port map (
            O => \N__60224\,
            I => \N__60165\
        );

    \I__13734\ : LocalMux
    port map (
            O => \N__60221\,
            I => \N__60165\
        );

    \I__13733\ : InMux
    port map (
            O => \N__60220\,
            I => \N__60162\
        );

    \I__13732\ : InMux
    port map (
            O => \N__60219\,
            I => \N__60159\
        );

    \I__13731\ : InMux
    port map (
            O => \N__60218\,
            I => \N__60152\
        );

    \I__13730\ : InMux
    port map (
            O => \N__60215\,
            I => \N__60152\
        );

    \I__13729\ : InMux
    port map (
            O => \N__60214\,
            I => \N__60147\
        );

    \I__13728\ : InMux
    port map (
            O => \N__60213\,
            I => \N__60147\
        );

    \I__13727\ : LocalMux
    port map (
            O => \N__60210\,
            I => \N__60144\
        );

    \I__13726\ : InMux
    port map (
            O => \N__60209\,
            I => \N__60139\
        );

    \I__13725\ : InMux
    port map (
            O => \N__60208\,
            I => \N__60139\
        );

    \I__13724\ : InMux
    port map (
            O => \N__60207\,
            I => \N__60134\
        );

    \I__13723\ : InMux
    port map (
            O => \N__60206\,
            I => \N__60134\
        );

    \I__13722\ : CascadeMux
    port map (
            O => \N__60205\,
            I => \N__60130\
        );

    \I__13721\ : LocalMux
    port map (
            O => \N__60202\,
            I => \N__60127\
        );

    \I__13720\ : LocalMux
    port map (
            O => \N__60199\,
            I => \N__60124\
        );

    \I__13719\ : InMux
    port map (
            O => \N__60198\,
            I => \N__60119\
        );

    \I__13718\ : InMux
    port map (
            O => \N__60197\,
            I => \N__60119\
        );

    \I__13717\ : InMux
    port map (
            O => \N__60196\,
            I => \N__60109\
        );

    \I__13716\ : InMux
    port map (
            O => \N__60193\,
            I => \N__60109\
        );

    \I__13715\ : InMux
    port map (
            O => \N__60192\,
            I => \N__60109\
        );

    \I__13714\ : InMux
    port map (
            O => \N__60191\,
            I => \N__60109\
        );

    \I__13713\ : InMux
    port map (
            O => \N__60190\,
            I => \N__60102\
        );

    \I__13712\ : InMux
    port map (
            O => \N__60189\,
            I => \N__60102\
        );

    \I__13711\ : InMux
    port map (
            O => \N__60188\,
            I => \N__60102\
        );

    \I__13710\ : InMux
    port map (
            O => \N__60187\,
            I => \N__60096\
        );

    \I__13709\ : Span4Mux_v
    port map (
            O => \N__60184\,
            I => \N__60093\
        );

    \I__13708\ : LocalMux
    port map (
            O => \N__60181\,
            I => \N__60090\
        );

    \I__13707\ : LocalMux
    port map (
            O => \N__60178\,
            I => \N__60087\
        );

    \I__13706\ : Span4Mux_h
    port map (
            O => \N__60173\,
            I => \N__60084\
        );

    \I__13705\ : LocalMux
    port map (
            O => \N__60170\,
            I => \N__60079\
        );

    \I__13704\ : Span4Mux_v
    port map (
            O => \N__60165\,
            I => \N__60079\
        );

    \I__13703\ : LocalMux
    port map (
            O => \N__60162\,
            I => \N__60074\
        );

    \I__13702\ : LocalMux
    port map (
            O => \N__60159\,
            I => \N__60074\
        );

    \I__13701\ : InMux
    port map (
            O => \N__60158\,
            I => \N__60069\
        );

    \I__13700\ : InMux
    port map (
            O => \N__60157\,
            I => \N__60069\
        );

    \I__13699\ : LocalMux
    port map (
            O => \N__60152\,
            I => \N__60066\
        );

    \I__13698\ : LocalMux
    port map (
            O => \N__60147\,
            I => \N__60057\
        );

    \I__13697\ : Span4Mux_h
    port map (
            O => \N__60144\,
            I => \N__60057\
        );

    \I__13696\ : LocalMux
    port map (
            O => \N__60139\,
            I => \N__60057\
        );

    \I__13695\ : LocalMux
    port map (
            O => \N__60134\,
            I => \N__60057\
        );

    \I__13694\ : InMux
    port map (
            O => \N__60133\,
            I => \N__60052\
        );

    \I__13693\ : InMux
    port map (
            O => \N__60130\,
            I => \N__60052\
        );

    \I__13692\ : Span4Mux_v
    port map (
            O => \N__60127\,
            I => \N__60045\
        );

    \I__13691\ : Span4Mux_v
    port map (
            O => \N__60124\,
            I => \N__60045\
        );

    \I__13690\ : LocalMux
    port map (
            O => \N__60119\,
            I => \N__60045\
        );

    \I__13689\ : InMux
    port map (
            O => \N__60118\,
            I => \N__60042\
        );

    \I__13688\ : LocalMux
    port map (
            O => \N__60109\,
            I => \N__60037\
        );

    \I__13687\ : LocalMux
    port map (
            O => \N__60102\,
            I => \N__60037\
        );

    \I__13686\ : InMux
    port map (
            O => \N__60101\,
            I => \N__60030\
        );

    \I__13685\ : InMux
    port map (
            O => \N__60100\,
            I => \N__60030\
        );

    \I__13684\ : InMux
    port map (
            O => \N__60099\,
            I => \N__60030\
        );

    \I__13683\ : LocalMux
    port map (
            O => \N__60096\,
            I => \N__60027\
        );

    \I__13682\ : Span4Mux_v
    port map (
            O => \N__60093\,
            I => \N__60024\
        );

    \I__13681\ : Span4Mux_v
    port map (
            O => \N__60090\,
            I => \N__60017\
        );

    \I__13680\ : Span4Mux_h
    port map (
            O => \N__60087\,
            I => \N__60017\
        );

    \I__13679\ : Span4Mux_v
    port map (
            O => \N__60084\,
            I => \N__60017\
        );

    \I__13678\ : Span4Mux_v
    port map (
            O => \N__60079\,
            I => \N__60010\
        );

    \I__13677\ : Span4Mux_h
    port map (
            O => \N__60074\,
            I => \N__60010\
        );

    \I__13676\ : LocalMux
    port map (
            O => \N__60069\,
            I => \N__60010\
        );

    \I__13675\ : Span4Mux_h
    port map (
            O => \N__60066\,
            I => \N__60007\
        );

    \I__13674\ : Span4Mux_h
    port map (
            O => \N__60057\,
            I => \N__60004\
        );

    \I__13673\ : LocalMux
    port map (
            O => \N__60052\,
            I => \N__59999\
        );

    \I__13672\ : Span4Mux_h
    port map (
            O => \N__60045\,
            I => \N__59999\
        );

    \I__13671\ : LocalMux
    port map (
            O => \N__60042\,
            I => \N__59992\
        );

    \I__13670\ : Span4Mux_v
    port map (
            O => \N__60037\,
            I => \N__59992\
        );

    \I__13669\ : LocalMux
    port map (
            O => \N__60030\,
            I => \N__59992\
        );

    \I__13668\ : Span12Mux_v
    port map (
            O => \N__60027\,
            I => \N__59989\
        );

    \I__13667\ : Span4Mux_h
    port map (
            O => \N__60024\,
            I => \N__59986\
        );

    \I__13666\ : Span4Mux_h
    port map (
            O => \N__60017\,
            I => \N__59983\
        );

    \I__13665\ : Span4Mux_v
    port map (
            O => \N__60010\,
            I => \N__59980\
        );

    \I__13664\ : Span4Mux_h
    port map (
            O => \N__60007\,
            I => \N__59975\
        );

    \I__13663\ : Span4Mux_v
    port map (
            O => \N__60004\,
            I => \N__59975\
        );

    \I__13662\ : Span4Mux_v
    port map (
            O => \N__59999\,
            I => \N__59970\
        );

    \I__13661\ : Span4Mux_h
    port map (
            O => \N__59992\,
            I => \N__59970\
        );

    \I__13660\ : Odrv12
    port map (
            O => \N__59989\,
            I => \aluOut_3\
        );

    \I__13659\ : Odrv4
    port map (
            O => \N__59986\,
            I => \aluOut_3\
        );

    \I__13658\ : Odrv4
    port map (
            O => \N__59983\,
            I => \aluOut_3\
        );

    \I__13657\ : Odrv4
    port map (
            O => \N__59980\,
            I => \aluOut_3\
        );

    \I__13656\ : Odrv4
    port map (
            O => \N__59975\,
            I => \aluOut_3\
        );

    \I__13655\ : Odrv4
    port map (
            O => \N__59970\,
            I => \aluOut_3\
        );

    \I__13654\ : CascadeMux
    port map (
            O => \N__59957\,
            I => \N__59954\
        );

    \I__13653\ : InMux
    port map (
            O => \N__59954\,
            I => \N__59951\
        );

    \I__13652\ : LocalMux
    port map (
            O => \N__59951\,
            I => \N__59948\
        );

    \I__13651\ : Span4Mux_h
    port map (
            O => \N__59948\,
            I => \N__59945\
        );

    \I__13650\ : Span4Mux_v
    port map (
            O => \N__59945\,
            I => \N__59942\
        );

    \I__13649\ : Sp12to4
    port map (
            O => \N__59942\,
            I => \N__59939\
        );

    \I__13648\ : Odrv12
    port map (
            O => \N__59939\,
            I => \ALU.d_RNI04H8GZ0Z_3\
        );

    \I__13647\ : InMux
    port map (
            O => \N__59936\,
            I => \N__59933\
        );

    \I__13646\ : LocalMux
    port map (
            O => \N__59933\,
            I => \N__59930\
        );

    \I__13645\ : Span4Mux_v
    port map (
            O => \N__59930\,
            I => \N__59926\
        );

    \I__13644\ : InMux
    port map (
            O => \N__59929\,
            I => \N__59923\
        );

    \I__13643\ : Span4Mux_h
    port map (
            O => \N__59926\,
            I => \N__59920\
        );

    \I__13642\ : LocalMux
    port map (
            O => \N__59923\,
            I => \ALU.addsub_3\
        );

    \I__13641\ : Odrv4
    port map (
            O => \N__59920\,
            I => \ALU.addsub_3\
        );

    \I__13640\ : InMux
    port map (
            O => \N__59915\,
            I => \ALU.addsub_cry_2\
        );

    \I__13639\ : CascadeMux
    port map (
            O => \N__59912\,
            I => \N__59907\
        );

    \I__13638\ : CascadeMux
    port map (
            O => \N__59911\,
            I => \N__59904\
        );

    \I__13637\ : InMux
    port map (
            O => \N__59910\,
            I => \N__59899\
        );

    \I__13636\ : InMux
    port map (
            O => \N__59907\,
            I => \N__59895\
        );

    \I__13635\ : InMux
    port map (
            O => \N__59904\,
            I => \N__59891\
        );

    \I__13634\ : InMux
    port map (
            O => \N__59903\,
            I => \N__59888\
        );

    \I__13633\ : CascadeMux
    port map (
            O => \N__59902\,
            I => \N__59885\
        );

    \I__13632\ : LocalMux
    port map (
            O => \N__59899\,
            I => \N__59878\
        );

    \I__13631\ : InMux
    port map (
            O => \N__59898\,
            I => \N__59875\
        );

    \I__13630\ : LocalMux
    port map (
            O => \N__59895\,
            I => \N__59870\
        );

    \I__13629\ : InMux
    port map (
            O => \N__59894\,
            I => \N__59867\
        );

    \I__13628\ : LocalMux
    port map (
            O => \N__59891\,
            I => \N__59861\
        );

    \I__13627\ : LocalMux
    port map (
            O => \N__59888\,
            I => \N__59858\
        );

    \I__13626\ : InMux
    port map (
            O => \N__59885\,
            I => \N__59853\
        );

    \I__13625\ : InMux
    port map (
            O => \N__59884\,
            I => \N__59853\
        );

    \I__13624\ : InMux
    port map (
            O => \N__59883\,
            I => \N__59850\
        );

    \I__13623\ : InMux
    port map (
            O => \N__59882\,
            I => \N__59846\
        );

    \I__13622\ : InMux
    port map (
            O => \N__59881\,
            I => \N__59843\
        );

    \I__13621\ : Span4Mux_v
    port map (
            O => \N__59878\,
            I => \N__59837\
        );

    \I__13620\ : LocalMux
    port map (
            O => \N__59875\,
            I => \N__59834\
        );

    \I__13619\ : InMux
    port map (
            O => \N__59874\,
            I => \N__59830\
        );

    \I__13618\ : InMux
    port map (
            O => \N__59873\,
            I => \N__59827\
        );

    \I__13617\ : Span4Mux_v
    port map (
            O => \N__59870\,
            I => \N__59824\
        );

    \I__13616\ : LocalMux
    port map (
            O => \N__59867\,
            I => \N__59821\
        );

    \I__13615\ : CascadeMux
    port map (
            O => \N__59866\,
            I => \N__59818\
        );

    \I__13614\ : InMux
    port map (
            O => \N__59865\,
            I => \N__59814\
        );

    \I__13613\ : InMux
    port map (
            O => \N__59864\,
            I => \N__59811\
        );

    \I__13612\ : Span4Mux_v
    port map (
            O => \N__59861\,
            I => \N__59806\
        );

    \I__13611\ : Span4Mux_v
    port map (
            O => \N__59858\,
            I => \N__59806\
        );

    \I__13610\ : LocalMux
    port map (
            O => \N__59853\,
            I => \N__59803\
        );

    \I__13609\ : LocalMux
    port map (
            O => \N__59850\,
            I => \N__59797\
        );

    \I__13608\ : InMux
    port map (
            O => \N__59849\,
            I => \N__59794\
        );

    \I__13607\ : LocalMux
    port map (
            O => \N__59846\,
            I => \N__59791\
        );

    \I__13606\ : LocalMux
    port map (
            O => \N__59843\,
            I => \N__59788\
        );

    \I__13605\ : InMux
    port map (
            O => \N__59842\,
            I => \N__59785\
        );

    \I__13604\ : InMux
    port map (
            O => \N__59841\,
            I => \N__59780\
        );

    \I__13603\ : InMux
    port map (
            O => \N__59840\,
            I => \N__59780\
        );

    \I__13602\ : Span4Mux_h
    port map (
            O => \N__59837\,
            I => \N__59775\
        );

    \I__13601\ : Span4Mux_v
    port map (
            O => \N__59834\,
            I => \N__59775\
        );

    \I__13600\ : InMux
    port map (
            O => \N__59833\,
            I => \N__59772\
        );

    \I__13599\ : LocalMux
    port map (
            O => \N__59830\,
            I => \N__59769\
        );

    \I__13598\ : LocalMux
    port map (
            O => \N__59827\,
            I => \N__59766\
        );

    \I__13597\ : Span4Mux_h
    port map (
            O => \N__59824\,
            I => \N__59761\
        );

    \I__13596\ : Span4Mux_v
    port map (
            O => \N__59821\,
            I => \N__59761\
        );

    \I__13595\ : InMux
    port map (
            O => \N__59818\,
            I => \N__59756\
        );

    \I__13594\ : InMux
    port map (
            O => \N__59817\,
            I => \N__59756\
        );

    \I__13593\ : LocalMux
    port map (
            O => \N__59814\,
            I => \N__59747\
        );

    \I__13592\ : LocalMux
    port map (
            O => \N__59811\,
            I => \N__59747\
        );

    \I__13591\ : Span4Mux_h
    port map (
            O => \N__59806\,
            I => \N__59747\
        );

    \I__13590\ : Span4Mux_v
    port map (
            O => \N__59803\,
            I => \N__59747\
        );

    \I__13589\ : InMux
    port map (
            O => \N__59802\,
            I => \N__59742\
        );

    \I__13588\ : InMux
    port map (
            O => \N__59801\,
            I => \N__59742\
        );

    \I__13587\ : InMux
    port map (
            O => \N__59800\,
            I => \N__59739\
        );

    \I__13586\ : Span12Mux_v
    port map (
            O => \N__59797\,
            I => \N__59732\
        );

    \I__13585\ : LocalMux
    port map (
            O => \N__59794\,
            I => \N__59732\
        );

    \I__13584\ : Span12Mux_s9_h
    port map (
            O => \N__59791\,
            I => \N__59732\
        );

    \I__13583\ : Sp12to4
    port map (
            O => \N__59788\,
            I => \N__59725\
        );

    \I__13582\ : LocalMux
    port map (
            O => \N__59785\,
            I => \N__59725\
        );

    \I__13581\ : LocalMux
    port map (
            O => \N__59780\,
            I => \N__59725\
        );

    \I__13580\ : Span4Mux_h
    port map (
            O => \N__59775\,
            I => \N__59718\
        );

    \I__13579\ : LocalMux
    port map (
            O => \N__59772\,
            I => \N__59718\
        );

    \I__13578\ : Span4Mux_v
    port map (
            O => \N__59769\,
            I => \N__59718\
        );

    \I__13577\ : Span4Mux_v
    port map (
            O => \N__59766\,
            I => \N__59713\
        );

    \I__13576\ : Span4Mux_v
    port map (
            O => \N__59761\,
            I => \N__59713\
        );

    \I__13575\ : LocalMux
    port map (
            O => \N__59756\,
            I => \N__59708\
        );

    \I__13574\ : Span4Mux_h
    port map (
            O => \N__59747\,
            I => \N__59708\
        );

    \I__13573\ : LocalMux
    port map (
            O => \N__59742\,
            I => \aluOut_4\
        );

    \I__13572\ : LocalMux
    port map (
            O => \N__59739\,
            I => \aluOut_4\
        );

    \I__13571\ : Odrv12
    port map (
            O => \N__59732\,
            I => \aluOut_4\
        );

    \I__13570\ : Odrv12
    port map (
            O => \N__59725\,
            I => \aluOut_4\
        );

    \I__13569\ : Odrv4
    port map (
            O => \N__59718\,
            I => \aluOut_4\
        );

    \I__13568\ : Odrv4
    port map (
            O => \N__59713\,
            I => \aluOut_4\
        );

    \I__13567\ : Odrv4
    port map (
            O => \N__59708\,
            I => \aluOut_4\
        );

    \I__13566\ : CascadeMux
    port map (
            O => \N__59693\,
            I => \N__59690\
        );

    \I__13565\ : InMux
    port map (
            O => \N__59690\,
            I => \N__59687\
        );

    \I__13564\ : LocalMux
    port map (
            O => \N__59687\,
            I => \N__59684\
        );

    \I__13563\ : Span4Mux_v
    port map (
            O => \N__59684\,
            I => \N__59681\
        );

    \I__13562\ : Sp12to4
    port map (
            O => \N__59681\,
            I => \N__59678\
        );

    \I__13561\ : Span12Mux_h
    port map (
            O => \N__59678\,
            I => \N__59675\
        );

    \I__13560\ : Odrv12
    port map (
            O => \N__59675\,
            I => \ALU.d_RNI7BF7IZ0Z_4\
        );

    \I__13559\ : InMux
    port map (
            O => \N__59672\,
            I => \N__59669\
        );

    \I__13558\ : LocalMux
    port map (
            O => \N__59669\,
            I => \N__59666\
        );

    \I__13557\ : Span12Mux_v
    port map (
            O => \N__59666\,
            I => \N__59662\
        );

    \I__13556\ : InMux
    port map (
            O => \N__59665\,
            I => \N__59659\
        );

    \I__13555\ : Span12Mux_h
    port map (
            O => \N__59662\,
            I => \N__59656\
        );

    \I__13554\ : LocalMux
    port map (
            O => \N__59659\,
            I => \N__59653\
        );

    \I__13553\ : Odrv12
    port map (
            O => \N__59656\,
            I => \ALU.addsub_4\
        );

    \I__13552\ : Odrv4
    port map (
            O => \N__59653\,
            I => \ALU.addsub_4\
        );

    \I__13551\ : InMux
    port map (
            O => \N__59648\,
            I => \ALU.addsub_cry_3\
        );

    \I__13550\ : CascadeMux
    port map (
            O => \N__59645\,
            I => \N__59641\
        );

    \I__13549\ : InMux
    port map (
            O => \N__59644\,
            I => \N__59634\
        );

    \I__13548\ : InMux
    port map (
            O => \N__59641\,
            I => \N__59629\
        );

    \I__13547\ : InMux
    port map (
            O => \N__59640\,
            I => \N__59629\
        );

    \I__13546\ : InMux
    port map (
            O => \N__59639\,
            I => \N__59626\
        );

    \I__13545\ : InMux
    port map (
            O => \N__59638\,
            I => \N__59621\
        );

    \I__13544\ : InMux
    port map (
            O => \N__59637\,
            I => \N__59615\
        );

    \I__13543\ : LocalMux
    port map (
            O => \N__59634\,
            I => \N__59612\
        );

    \I__13542\ : LocalMux
    port map (
            O => \N__59629\,
            I => \N__59609\
        );

    \I__13541\ : LocalMux
    port map (
            O => \N__59626\,
            I => \N__59606\
        );

    \I__13540\ : InMux
    port map (
            O => \N__59625\,
            I => \N__59603\
        );

    \I__13539\ : CascadeMux
    port map (
            O => \N__59624\,
            I => \N__59596\
        );

    \I__13538\ : LocalMux
    port map (
            O => \N__59621\,
            I => \N__59592\
        );

    \I__13537\ : InMux
    port map (
            O => \N__59620\,
            I => \N__59589\
        );

    \I__13536\ : InMux
    port map (
            O => \N__59619\,
            I => \N__59577\
        );

    \I__13535\ : InMux
    port map (
            O => \N__59618\,
            I => \N__59577\
        );

    \I__13534\ : LocalMux
    port map (
            O => \N__59615\,
            I => \N__59574\
        );

    \I__13533\ : Span4Mux_v
    port map (
            O => \N__59612\,
            I => \N__59567\
        );

    \I__13532\ : Span4Mux_v
    port map (
            O => \N__59609\,
            I => \N__59567\
        );

    \I__13531\ : Span4Mux_v
    port map (
            O => \N__59606\,
            I => \N__59567\
        );

    \I__13530\ : LocalMux
    port map (
            O => \N__59603\,
            I => \N__59564\
        );

    \I__13529\ : InMux
    port map (
            O => \N__59602\,
            I => \N__59557\
        );

    \I__13528\ : InMux
    port map (
            O => \N__59601\,
            I => \N__59557\
        );

    \I__13527\ : InMux
    port map (
            O => \N__59600\,
            I => \N__59557\
        );

    \I__13526\ : CascadeMux
    port map (
            O => \N__59599\,
            I => \N__59554\
        );

    \I__13525\ : InMux
    port map (
            O => \N__59596\,
            I => \N__59551\
        );

    \I__13524\ : InMux
    port map (
            O => \N__59595\,
            I => \N__59546\
        );

    \I__13523\ : Span4Mux_h
    port map (
            O => \N__59592\,
            I => \N__59541\
        );

    \I__13522\ : LocalMux
    port map (
            O => \N__59589\,
            I => \N__59541\
        );

    \I__13521\ : InMux
    port map (
            O => \N__59588\,
            I => \N__59537\
        );

    \I__13520\ : InMux
    port map (
            O => \N__59587\,
            I => \N__59534\
        );

    \I__13519\ : InMux
    port map (
            O => \N__59586\,
            I => \N__59531\
        );

    \I__13518\ : InMux
    port map (
            O => \N__59585\,
            I => \N__59528\
        );

    \I__13517\ : InMux
    port map (
            O => \N__59584\,
            I => \N__59521\
        );

    \I__13516\ : InMux
    port map (
            O => \N__59583\,
            I => \N__59521\
        );

    \I__13515\ : InMux
    port map (
            O => \N__59582\,
            I => \N__59521\
        );

    \I__13514\ : LocalMux
    port map (
            O => \N__59577\,
            I => \N__59518\
        );

    \I__13513\ : Span4Mux_v
    port map (
            O => \N__59574\,
            I => \N__59515\
        );

    \I__13512\ : Span4Mux_h
    port map (
            O => \N__59567\,
            I => \N__59512\
        );

    \I__13511\ : Span4Mux_h
    port map (
            O => \N__59564\,
            I => \N__59507\
        );

    \I__13510\ : LocalMux
    port map (
            O => \N__59557\,
            I => \N__59507\
        );

    \I__13509\ : InMux
    port map (
            O => \N__59554\,
            I => \N__59504\
        );

    \I__13508\ : LocalMux
    port map (
            O => \N__59551\,
            I => \N__59500\
        );

    \I__13507\ : InMux
    port map (
            O => \N__59550\,
            I => \N__59497\
        );

    \I__13506\ : InMux
    port map (
            O => \N__59549\,
            I => \N__59494\
        );

    \I__13505\ : LocalMux
    port map (
            O => \N__59546\,
            I => \N__59491\
        );

    \I__13504\ : Span4Mux_h
    port map (
            O => \N__59541\,
            I => \N__59488\
        );

    \I__13503\ : CascadeMux
    port map (
            O => \N__59540\,
            I => \N__59480\
        );

    \I__13502\ : LocalMux
    port map (
            O => \N__59537\,
            I => \N__59473\
        );

    \I__13501\ : LocalMux
    port map (
            O => \N__59534\,
            I => \N__59470\
        );

    \I__13500\ : LocalMux
    port map (
            O => \N__59531\,
            I => \N__59463\
        );

    \I__13499\ : LocalMux
    port map (
            O => \N__59528\,
            I => \N__59463\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__59521\,
            I => \N__59463\
        );

    \I__13497\ : Span4Mux_v
    port map (
            O => \N__59518\,
            I => \N__59454\
        );

    \I__13496\ : Span4Mux_h
    port map (
            O => \N__59515\,
            I => \N__59454\
        );

    \I__13495\ : Span4Mux_h
    port map (
            O => \N__59512\,
            I => \N__59454\
        );

    \I__13494\ : Span4Mux_v
    port map (
            O => \N__59507\,
            I => \N__59454\
        );

    \I__13493\ : LocalMux
    port map (
            O => \N__59504\,
            I => \N__59451\
        );

    \I__13492\ : InMux
    port map (
            O => \N__59503\,
            I => \N__59448\
        );

    \I__13491\ : Span4Mux_h
    port map (
            O => \N__59500\,
            I => \N__59439\
        );

    \I__13490\ : LocalMux
    port map (
            O => \N__59497\,
            I => \N__59439\
        );

    \I__13489\ : LocalMux
    port map (
            O => \N__59494\,
            I => \N__59439\
        );

    \I__13488\ : Span4Mux_v
    port map (
            O => \N__59491\,
            I => \N__59439\
        );

    \I__13487\ : Span4Mux_h
    port map (
            O => \N__59488\,
            I => \N__59436\
        );

    \I__13486\ : InMux
    port map (
            O => \N__59487\,
            I => \N__59431\
        );

    \I__13485\ : InMux
    port map (
            O => \N__59486\,
            I => \N__59431\
        );

    \I__13484\ : InMux
    port map (
            O => \N__59485\,
            I => \N__59424\
        );

    \I__13483\ : InMux
    port map (
            O => \N__59484\,
            I => \N__59424\
        );

    \I__13482\ : InMux
    port map (
            O => \N__59483\,
            I => \N__59424\
        );

    \I__13481\ : InMux
    port map (
            O => \N__59480\,
            I => \N__59413\
        );

    \I__13480\ : InMux
    port map (
            O => \N__59479\,
            I => \N__59413\
        );

    \I__13479\ : InMux
    port map (
            O => \N__59478\,
            I => \N__59413\
        );

    \I__13478\ : InMux
    port map (
            O => \N__59477\,
            I => \N__59413\
        );

    \I__13477\ : InMux
    port map (
            O => \N__59476\,
            I => \N__59413\
        );

    \I__13476\ : Span4Mux_h
    port map (
            O => \N__59473\,
            I => \N__59406\
        );

    \I__13475\ : Span4Mux_v
    port map (
            O => \N__59470\,
            I => \N__59406\
        );

    \I__13474\ : Span4Mux_h
    port map (
            O => \N__59463\,
            I => \N__59406\
        );

    \I__13473\ : Span4Mux_h
    port map (
            O => \N__59454\,
            I => \N__59403\
        );

    \I__13472\ : Odrv12
    port map (
            O => \N__59451\,
            I => \aluOut_5\
        );

    \I__13471\ : LocalMux
    port map (
            O => \N__59448\,
            I => \aluOut_5\
        );

    \I__13470\ : Odrv4
    port map (
            O => \N__59439\,
            I => \aluOut_5\
        );

    \I__13469\ : Odrv4
    port map (
            O => \N__59436\,
            I => \aluOut_5\
        );

    \I__13468\ : LocalMux
    port map (
            O => \N__59431\,
            I => \aluOut_5\
        );

    \I__13467\ : LocalMux
    port map (
            O => \N__59424\,
            I => \aluOut_5\
        );

    \I__13466\ : LocalMux
    port map (
            O => \N__59413\,
            I => \aluOut_5\
        );

    \I__13465\ : Odrv4
    port map (
            O => \N__59406\,
            I => \aluOut_5\
        );

    \I__13464\ : Odrv4
    port map (
            O => \N__59403\,
            I => \aluOut_5\
        );

    \I__13463\ : CascadeMux
    port map (
            O => \N__59384\,
            I => \N__59381\
        );

    \I__13462\ : InMux
    port map (
            O => \N__59381\,
            I => \N__59378\
        );

    \I__13461\ : LocalMux
    port map (
            O => \N__59378\,
            I => \N__59375\
        );

    \I__13460\ : Span12Mux_s10_h
    port map (
            O => \N__59375\,
            I => \N__59372\
        );

    \I__13459\ : Odrv12
    port map (
            O => \N__59372\,
            I => \ALU.d_RNI58QFIZ0Z_5\
        );

    \I__13458\ : InMux
    port map (
            O => \N__59369\,
            I => \N__59366\
        );

    \I__13457\ : LocalMux
    port map (
            O => \N__59366\,
            I => \N__59363\
        );

    \I__13456\ : Span4Mux_h
    port map (
            O => \N__59363\,
            I => \N__59360\
        );

    \I__13455\ : Span4Mux_h
    port map (
            O => \N__59360\,
            I => \N__59357\
        );

    \I__13454\ : Span4Mux_h
    port map (
            O => \N__59357\,
            I => \N__59354\
        );

    \I__13453\ : Span4Mux_v
    port map (
            O => \N__59354\,
            I => \N__59350\
        );

    \I__13452\ : InMux
    port map (
            O => \N__59353\,
            I => \N__59347\
        );

    \I__13451\ : Odrv4
    port map (
            O => \N__59350\,
            I => \ALU.addsub_5\
        );

    \I__13450\ : LocalMux
    port map (
            O => \N__59347\,
            I => \ALU.addsub_5\
        );

    \I__13449\ : InMux
    port map (
            O => \N__59342\,
            I => \ALU.addsub_cry_4\
        );

    \I__13448\ : InMux
    port map (
            O => \N__59339\,
            I => \N__59335\
        );

    \I__13447\ : InMux
    port map (
            O => \N__59338\,
            I => \N__59332\
        );

    \I__13446\ : LocalMux
    port map (
            O => \N__59335\,
            I => \N__59329\
        );

    \I__13445\ : LocalMux
    port map (
            O => \N__59332\,
            I => \N__59325\
        );

    \I__13444\ : Span4Mux_v
    port map (
            O => \N__59329\,
            I => \N__59322\
        );

    \I__13443\ : InMux
    port map (
            O => \N__59328\,
            I => \N__59319\
        );

    \I__13442\ : Span4Mux_h
    port map (
            O => \N__59325\,
            I => \N__59316\
        );

    \I__13441\ : Span4Mux_h
    port map (
            O => \N__59322\,
            I => \N__59313\
        );

    \I__13440\ : LocalMux
    port map (
            O => \N__59319\,
            I => \ALU.a_15_m2_sZ0Z_15\
        );

    \I__13439\ : Odrv4
    port map (
            O => \N__59316\,
            I => \ALU.a_15_m2_sZ0Z_15\
        );

    \I__13438\ : Odrv4
    port map (
            O => \N__59313\,
            I => \ALU.a_15_m2_sZ0Z_15\
        );

    \I__13437\ : InMux
    port map (
            O => \N__59306\,
            I => \N__59302\
        );

    \I__13436\ : InMux
    port map (
            O => \N__59305\,
            I => \N__59299\
        );

    \I__13435\ : LocalMux
    port map (
            O => \N__59302\,
            I => \N__59292\
        );

    \I__13434\ : LocalMux
    port map (
            O => \N__59299\,
            I => \N__59283\
        );

    \I__13433\ : InMux
    port map (
            O => \N__59298\,
            I => \N__59276\
        );

    \I__13432\ : InMux
    port map (
            O => \N__59297\,
            I => \N__59276\
        );

    \I__13431\ : InMux
    port map (
            O => \N__59296\,
            I => \N__59271\
        );

    \I__13430\ : InMux
    port map (
            O => \N__59295\,
            I => \N__59271\
        );

    \I__13429\ : Span4Mux_v
    port map (
            O => \N__59292\,
            I => \N__59268\
        );

    \I__13428\ : InMux
    port map (
            O => \N__59291\,
            I => \N__59263\
        );

    \I__13427\ : InMux
    port map (
            O => \N__59290\,
            I => \N__59259\
        );

    \I__13426\ : InMux
    port map (
            O => \N__59289\,
            I => \N__59250\
        );

    \I__13425\ : InMux
    port map (
            O => \N__59288\,
            I => \N__59250\
        );

    \I__13424\ : InMux
    port map (
            O => \N__59287\,
            I => \N__59250\
        );

    \I__13423\ : InMux
    port map (
            O => \N__59286\,
            I => \N__59250\
        );

    \I__13422\ : Span4Mux_v
    port map (
            O => \N__59283\,
            I => \N__59245\
        );

    \I__13421\ : InMux
    port map (
            O => \N__59282\,
            I => \N__59240\
        );

    \I__13420\ : InMux
    port map (
            O => \N__59281\,
            I => \N__59240\
        );

    \I__13419\ : LocalMux
    port map (
            O => \N__59276\,
            I => \N__59235\
        );

    \I__13418\ : LocalMux
    port map (
            O => \N__59271\,
            I => \N__59235\
        );

    \I__13417\ : Span4Mux_h
    port map (
            O => \N__59268\,
            I => \N__59232\
        );

    \I__13416\ : InMux
    port map (
            O => \N__59267\,
            I => \N__59229\
        );

    \I__13415\ : InMux
    port map (
            O => \N__59266\,
            I => \N__59226\
        );

    \I__13414\ : LocalMux
    port map (
            O => \N__59263\,
            I => \N__59223\
        );

    \I__13413\ : InMux
    port map (
            O => \N__59262\,
            I => \N__59220\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__59259\,
            I => \N__59215\
        );

    \I__13411\ : LocalMux
    port map (
            O => \N__59250\,
            I => \N__59215\
        );

    \I__13410\ : InMux
    port map (
            O => \N__59249\,
            I => \N__59212\
        );

    \I__13409\ : InMux
    port map (
            O => \N__59248\,
            I => \N__59209\
        );

    \I__13408\ : Sp12to4
    port map (
            O => \N__59245\,
            I => \N__59202\
        );

    \I__13407\ : LocalMux
    port map (
            O => \N__59240\,
            I => \N__59202\
        );

    \I__13406\ : Span12Mux_v
    port map (
            O => \N__59235\,
            I => \N__59202\
        );

    \I__13405\ : Span4Mux_v
    port map (
            O => \N__59232\,
            I => \N__59195\
        );

    \I__13404\ : LocalMux
    port map (
            O => \N__59229\,
            I => \N__59195\
        );

    \I__13403\ : LocalMux
    port map (
            O => \N__59226\,
            I => \N__59195\
        );

    \I__13402\ : Span4Mux_h
    port map (
            O => \N__59223\,
            I => \N__59188\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__59220\,
            I => \N__59188\
        );

    \I__13400\ : Span4Mux_h
    port map (
            O => \N__59215\,
            I => \N__59188\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__59212\,
            I => \ALU.a_15_sm0\
        );

    \I__13398\ : LocalMux
    port map (
            O => \N__59209\,
            I => \ALU.a_15_sm0\
        );

    \I__13397\ : Odrv12
    port map (
            O => \N__59202\,
            I => \ALU.a_15_sm0\
        );

    \I__13396\ : Odrv4
    port map (
            O => \N__59195\,
            I => \ALU.a_15_sm0\
        );

    \I__13395\ : Odrv4
    port map (
            O => \N__59188\,
            I => \ALU.a_15_sm0\
        );

    \I__13394\ : CascadeMux
    port map (
            O => \N__59177\,
            I => \N__59173\
        );

    \I__13393\ : CascadeMux
    port map (
            O => \N__59176\,
            I => \N__59170\
        );

    \I__13392\ : InMux
    port map (
            O => \N__59173\,
            I => \N__59166\
        );

    \I__13391\ : InMux
    port map (
            O => \N__59170\,
            I => \N__59163\
        );

    \I__13390\ : InMux
    port map (
            O => \N__59169\,
            I => \N__59160\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__59166\,
            I => \N__59151\
        );

    \I__13388\ : LocalMux
    port map (
            O => \N__59163\,
            I => \N__59151\
        );

    \I__13387\ : LocalMux
    port map (
            O => \N__59160\,
            I => \N__59151\
        );

    \I__13386\ : InMux
    port map (
            O => \N__59159\,
            I => \N__59146\
        );

    \I__13385\ : InMux
    port map (
            O => \N__59158\,
            I => \N__59146\
        );

    \I__13384\ : Span4Mux_v
    port map (
            O => \N__59151\,
            I => \N__59133\
        );

    \I__13383\ : LocalMux
    port map (
            O => \N__59146\,
            I => \N__59130\
        );

    \I__13382\ : InMux
    port map (
            O => \N__59145\,
            I => \N__59125\
        );

    \I__13381\ : InMux
    port map (
            O => \N__59144\,
            I => \N__59125\
        );

    \I__13380\ : CascadeMux
    port map (
            O => \N__59143\,
            I => \N__59121\
        );

    \I__13379\ : CascadeMux
    port map (
            O => \N__59142\,
            I => \N__59117\
        );

    \I__13378\ : CascadeMux
    port map (
            O => \N__59141\,
            I => \N__59114\
        );

    \I__13377\ : CascadeMux
    port map (
            O => \N__59140\,
            I => \N__59111\
        );

    \I__13376\ : CascadeMux
    port map (
            O => \N__59139\,
            I => \N__59108\
        );

    \I__13375\ : CascadeMux
    port map (
            O => \N__59138\,
            I => \N__59103\
        );

    \I__13374\ : InMux
    port map (
            O => \N__59137\,
            I => \N__59095\
        );

    \I__13373\ : InMux
    port map (
            O => \N__59136\,
            I => \N__59095\
        );

    \I__13372\ : Span4Mux_v
    port map (
            O => \N__59133\,
            I => \N__59088\
        );

    \I__13371\ : Span4Mux_h
    port map (
            O => \N__59130\,
            I => \N__59088\
        );

    \I__13370\ : LocalMux
    port map (
            O => \N__59125\,
            I => \N__59088\
        );

    \I__13369\ : InMux
    port map (
            O => \N__59124\,
            I => \N__59085\
        );

    \I__13368\ : InMux
    port map (
            O => \N__59121\,
            I => \N__59082\
        );

    \I__13367\ : CascadeMux
    port map (
            O => \N__59120\,
            I => \N__59079\
        );

    \I__13366\ : InMux
    port map (
            O => \N__59117\,
            I => \N__59076\
        );

    \I__13365\ : InMux
    port map (
            O => \N__59114\,
            I => \N__59073\
        );

    \I__13364\ : InMux
    port map (
            O => \N__59111\,
            I => \N__59070\
        );

    \I__13363\ : InMux
    port map (
            O => \N__59108\,
            I => \N__59067\
        );

    \I__13362\ : InMux
    port map (
            O => \N__59107\,
            I => \N__59059\
        );

    \I__13361\ : InMux
    port map (
            O => \N__59106\,
            I => \N__59059\
        );

    \I__13360\ : InMux
    port map (
            O => \N__59103\,
            I => \N__59059\
        );

    \I__13359\ : InMux
    port map (
            O => \N__59102\,
            I => \N__59056\
        );

    \I__13358\ : InMux
    port map (
            O => \N__59101\,
            I => \N__59051\
        );

    \I__13357\ : InMux
    port map (
            O => \N__59100\,
            I => \N__59051\
        );

    \I__13356\ : LocalMux
    port map (
            O => \N__59095\,
            I => \N__59045\
        );

    \I__13355\ : Span4Mux_h
    port map (
            O => \N__59088\,
            I => \N__59037\
        );

    \I__13354\ : LocalMux
    port map (
            O => \N__59085\,
            I => \N__59037\
        );

    \I__13353\ : LocalMux
    port map (
            O => \N__59082\,
            I => \N__59034\
        );

    \I__13352\ : InMux
    port map (
            O => \N__59079\,
            I => \N__59031\
        );

    \I__13351\ : LocalMux
    port map (
            O => \N__59076\,
            I => \N__59024\
        );

    \I__13350\ : LocalMux
    port map (
            O => \N__59073\,
            I => \N__59024\
        );

    \I__13349\ : LocalMux
    port map (
            O => \N__59070\,
            I => \N__59024\
        );

    \I__13348\ : LocalMux
    port map (
            O => \N__59067\,
            I => \N__59021\
        );

    \I__13347\ : InMux
    port map (
            O => \N__59066\,
            I => \N__59018\
        );

    \I__13346\ : LocalMux
    port map (
            O => \N__59059\,
            I => \N__59013\
        );

    \I__13345\ : LocalMux
    port map (
            O => \N__59056\,
            I => \N__59013\
        );

    \I__13344\ : LocalMux
    port map (
            O => \N__59051\,
            I => \N__59010\
        );

    \I__13343\ : CascadeMux
    port map (
            O => \N__59050\,
            I => \N__59006\
        );

    \I__13342\ : CascadeMux
    port map (
            O => \N__59049\,
            I => \N__59002\
        );

    \I__13341\ : CascadeMux
    port map (
            O => \N__59048\,
            I => \N__58998\
        );

    \I__13340\ : Span4Mux_v
    port map (
            O => \N__59045\,
            I => \N__58995\
        );

    \I__13339\ : InMux
    port map (
            O => \N__59044\,
            I => \N__58988\
        );

    \I__13338\ : InMux
    port map (
            O => \N__59043\,
            I => \N__58988\
        );

    \I__13337\ : InMux
    port map (
            O => \N__59042\,
            I => \N__58988\
        );

    \I__13336\ : Span4Mux_v
    port map (
            O => \N__59037\,
            I => \N__58984\
        );

    \I__13335\ : Span4Mux_v
    port map (
            O => \N__59034\,
            I => \N__58981\
        );

    \I__13334\ : LocalMux
    port map (
            O => \N__59031\,
            I => \N__58976\
        );

    \I__13333\ : Span4Mux_v
    port map (
            O => \N__59024\,
            I => \N__58976\
        );

    \I__13332\ : Span4Mux_v
    port map (
            O => \N__59021\,
            I => \N__58971\
        );

    \I__13331\ : LocalMux
    port map (
            O => \N__59018\,
            I => \N__58971\
        );

    \I__13330\ : Span4Mux_v
    port map (
            O => \N__59013\,
            I => \N__58968\
        );

    \I__13329\ : Span4Mux_h
    port map (
            O => \N__59010\,
            I => \N__58965\
        );

    \I__13328\ : InMux
    port map (
            O => \N__59009\,
            I => \N__58958\
        );

    \I__13327\ : InMux
    port map (
            O => \N__59006\,
            I => \N__58958\
        );

    \I__13326\ : InMux
    port map (
            O => \N__59005\,
            I => \N__58958\
        );

    \I__13325\ : InMux
    port map (
            O => \N__59002\,
            I => \N__58951\
        );

    \I__13324\ : InMux
    port map (
            O => \N__59001\,
            I => \N__58951\
        );

    \I__13323\ : InMux
    port map (
            O => \N__58998\,
            I => \N__58951\
        );

    \I__13322\ : Span4Mux_h
    port map (
            O => \N__58995\,
            I => \N__58946\
        );

    \I__13321\ : LocalMux
    port map (
            O => \N__58988\,
            I => \N__58946\
        );

    \I__13320\ : InMux
    port map (
            O => \N__58987\,
            I => \N__58943\
        );

    \I__13319\ : Sp12to4
    port map (
            O => \N__58984\,
            I => \N__58940\
        );

    \I__13318\ : Span4Mux_h
    port map (
            O => \N__58981\,
            I => \N__58933\
        );

    \I__13317\ : Span4Mux_v
    port map (
            O => \N__58976\,
            I => \N__58933\
        );

    \I__13316\ : Span4Mux_v
    port map (
            O => \N__58971\,
            I => \N__58933\
        );

    \I__13315\ : Span4Mux_v
    port map (
            O => \N__58968\,
            I => \N__58930\
        );

    \I__13314\ : Span4Mux_v
    port map (
            O => \N__58965\,
            I => \N__58927\
        );

    \I__13313\ : LocalMux
    port map (
            O => \N__58958\,
            I => \N__58920\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__58951\,
            I => \N__58920\
        );

    \I__13311\ : Span4Mux_h
    port map (
            O => \N__58946\,
            I => \N__58920\
        );

    \I__13310\ : LocalMux
    port map (
            O => \N__58943\,
            I => \N__58915\
        );

    \I__13309\ : Span12Mux_h
    port map (
            O => \N__58940\,
            I => \N__58915\
        );

    \I__13308\ : Sp12to4
    port map (
            O => \N__58933\,
            I => \N__58910\
        );

    \I__13307\ : Sp12to4
    port map (
            O => \N__58930\,
            I => \N__58910\
        );

    \I__13306\ : Span4Mux_v
    port map (
            O => \N__58927\,
            I => \N__58907\
        );

    \I__13305\ : Span4Mux_v
    port map (
            O => \N__58920\,
            I => \N__58904\
        );

    \I__13304\ : Span12Mux_v
    port map (
            O => \N__58915\,
            I => \N__58899\
        );

    \I__13303\ : Span12Mux_h
    port map (
            O => \N__58910\,
            I => \N__58899\
        );

    \I__13302\ : Span4Mux_h
    port map (
            O => \N__58907\,
            I => \N__58894\
        );

    \I__13301\ : Span4Mux_v
    port map (
            O => \N__58904\,
            I => \N__58894\
        );

    \I__13300\ : Odrv12
    port map (
            O => \N__58899\,
            I => \aluOperation_1\
        );

    \I__13299\ : Odrv4
    port map (
            O => \N__58894\,
            I => \aluOperation_1\
        );

    \I__13298\ : InMux
    port map (
            O => \N__58889\,
            I => \N__58881\
        );

    \I__13297\ : InMux
    port map (
            O => \N__58888\,
            I => \N__58878\
        );

    \I__13296\ : InMux
    port map (
            O => \N__58887\,
            I => \N__58874\
        );

    \I__13295\ : InMux
    port map (
            O => \N__58886\,
            I => \N__58871\
        );

    \I__13294\ : InMux
    port map (
            O => \N__58885\,
            I => \N__58868\
        );

    \I__13293\ : InMux
    port map (
            O => \N__58884\,
            I => \N__58865\
        );

    \I__13292\ : LocalMux
    port map (
            O => \N__58881\,
            I => \N__58861\
        );

    \I__13291\ : LocalMux
    port map (
            O => \N__58878\,
            I => \N__58858\
        );

    \I__13290\ : InMux
    port map (
            O => \N__58877\,
            I => \N__58855\
        );

    \I__13289\ : LocalMux
    port map (
            O => \N__58874\,
            I => \N__58850\
        );

    \I__13288\ : LocalMux
    port map (
            O => \N__58871\,
            I => \N__58850\
        );

    \I__13287\ : LocalMux
    port map (
            O => \N__58868\,
            I => \N__58845\
        );

    \I__13286\ : LocalMux
    port map (
            O => \N__58865\,
            I => \N__58845\
        );

    \I__13285\ : InMux
    port map (
            O => \N__58864\,
            I => \N__58842\
        );

    \I__13284\ : Span4Mux_h
    port map (
            O => \N__58861\,
            I => \N__58839\
        );

    \I__13283\ : Span4Mux_h
    port map (
            O => \N__58858\,
            I => \N__58836\
        );

    \I__13282\ : LocalMux
    port map (
            O => \N__58855\,
            I => \N__58831\
        );

    \I__13281\ : Span4Mux_v
    port map (
            O => \N__58850\,
            I => \N__58831\
        );

    \I__13280\ : Span4Mux_v
    port map (
            O => \N__58845\,
            I => \N__58828\
        );

    \I__13279\ : LocalMux
    port map (
            O => \N__58842\,
            I => \ALU.a_15_ns_1_7\
        );

    \I__13278\ : Odrv4
    port map (
            O => \N__58839\,
            I => \ALU.a_15_ns_1_7\
        );

    \I__13277\ : Odrv4
    port map (
            O => \N__58836\,
            I => \ALU.a_15_ns_1_7\
        );

    \I__13276\ : Odrv4
    port map (
            O => \N__58831\,
            I => \ALU.a_15_ns_1_7\
        );

    \I__13275\ : Odrv4
    port map (
            O => \N__58828\,
            I => \ALU.a_15_ns_1_7\
        );

    \I__13274\ : InMux
    port map (
            O => \N__58817\,
            I => \N__58813\
        );

    \I__13273\ : InMux
    port map (
            O => \N__58816\,
            I => \N__58809\
        );

    \I__13272\ : LocalMux
    port map (
            O => \N__58813\,
            I => \N__58805\
        );

    \I__13271\ : InMux
    port map (
            O => \N__58812\,
            I => \N__58802\
        );

    \I__13270\ : LocalMux
    port map (
            O => \N__58809\,
            I => \N__58796\
        );

    \I__13269\ : InMux
    port map (
            O => \N__58808\,
            I => \N__58793\
        );

    \I__13268\ : Span4Mux_h
    port map (
            O => \N__58805\,
            I => \N__58790\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__58802\,
            I => \N__58787\
        );

    \I__13266\ : InMux
    port map (
            O => \N__58801\,
            I => \N__58784\
        );

    \I__13265\ : InMux
    port map (
            O => \N__58800\,
            I => \N__58781\
        );

    \I__13264\ : InMux
    port map (
            O => \N__58799\,
            I => \N__58778\
        );

    \I__13263\ : Span4Mux_v
    port map (
            O => \N__58796\,
            I => \N__58773\
        );

    \I__13262\ : LocalMux
    port map (
            O => \N__58793\,
            I => \N__58773\
        );

    \I__13261\ : Span4Mux_h
    port map (
            O => \N__58790\,
            I => \N__58768\
        );

    \I__13260\ : Span4Mux_v
    port map (
            O => \N__58787\,
            I => \N__58768\
        );

    \I__13259\ : LocalMux
    port map (
            O => \N__58784\,
            I => \ALU.mult_388_c_RNIPGN6QZ0Z7\
        );

    \I__13258\ : LocalMux
    port map (
            O => \N__58781\,
            I => \ALU.mult_388_c_RNIPGN6QZ0Z7\
        );

    \I__13257\ : LocalMux
    port map (
            O => \N__58778\,
            I => \ALU.mult_388_c_RNIPGN6QZ0Z7\
        );

    \I__13256\ : Odrv4
    port map (
            O => \N__58773\,
            I => \ALU.mult_388_c_RNIPGN6QZ0Z7\
        );

    \I__13255\ : Odrv4
    port map (
            O => \N__58768\,
            I => \ALU.mult_388_c_RNIPGN6QZ0Z7\
        );

    \I__13254\ : InMux
    port map (
            O => \N__58757\,
            I => \N__58753\
        );

    \I__13253\ : CascadeMux
    port map (
            O => \N__58756\,
            I => \N__58749\
        );

    \I__13252\ : LocalMux
    port map (
            O => \N__58753\,
            I => \N__58746\
        );

    \I__13251\ : InMux
    port map (
            O => \N__58752\,
            I => \N__58742\
        );

    \I__13250\ : InMux
    port map (
            O => \N__58749\,
            I => \N__58736\
        );

    \I__13249\ : Span4Mux_v
    port map (
            O => \N__58746\,
            I => \N__58733\
        );

    \I__13248\ : InMux
    port map (
            O => \N__58745\,
            I => \N__58730\
        );

    \I__13247\ : LocalMux
    port map (
            O => \N__58742\,
            I => \N__58727\
        );

    \I__13246\ : InMux
    port map (
            O => \N__58741\,
            I => \N__58724\
        );

    \I__13245\ : InMux
    port map (
            O => \N__58740\,
            I => \N__58721\
        );

    \I__13244\ : InMux
    port map (
            O => \N__58739\,
            I => \N__58718\
        );

    \I__13243\ : LocalMux
    port map (
            O => \N__58736\,
            I => \N__58714\
        );

    \I__13242\ : Span4Mux_h
    port map (
            O => \N__58733\,
            I => \N__58709\
        );

    \I__13241\ : LocalMux
    port map (
            O => \N__58730\,
            I => \N__58709\
        );

    \I__13240\ : Span4Mux_v
    port map (
            O => \N__58727\,
            I => \N__58706\
        );

    \I__13239\ : LocalMux
    port map (
            O => \N__58724\,
            I => \N__58699\
        );

    \I__13238\ : LocalMux
    port map (
            O => \N__58721\,
            I => \N__58699\
        );

    \I__13237\ : LocalMux
    port map (
            O => \N__58718\,
            I => \N__58699\
        );

    \I__13236\ : InMux
    port map (
            O => \N__58717\,
            I => \N__58696\
        );

    \I__13235\ : Span4Mux_v
    port map (
            O => \N__58714\,
            I => \N__58691\
        );

    \I__13234\ : Span4Mux_v
    port map (
            O => \N__58709\,
            I => \N__58691\
        );

    \I__13233\ : Span4Mux_h
    port map (
            O => \N__58706\,
            I => \N__58684\
        );

    \I__13232\ : Span4Mux_v
    port map (
            O => \N__58699\,
            I => \N__58684\
        );

    \I__13231\ : LocalMux
    port map (
            O => \N__58696\,
            I => \N__58684\
        );

    \I__13230\ : Odrv4
    port map (
            O => \N__58691\,
            I => \ALU.rshift_3\
        );

    \I__13229\ : Odrv4
    port map (
            O => \N__58684\,
            I => \ALU.rshift_3\
        );

    \I__13228\ : InMux
    port map (
            O => \N__58679\,
            I => \N__58673\
        );

    \I__13227\ : InMux
    port map (
            O => \N__58678\,
            I => \N__58670\
        );

    \I__13226\ : InMux
    port map (
            O => \N__58677\,
            I => \N__58667\
        );

    \I__13225\ : InMux
    port map (
            O => \N__58676\,
            I => \N__58660\
        );

    \I__13224\ : LocalMux
    port map (
            O => \N__58673\,
            I => \N__58657\
        );

    \I__13223\ : LocalMux
    port map (
            O => \N__58670\,
            I => \N__58654\
        );

    \I__13222\ : LocalMux
    port map (
            O => \N__58667\,
            I => \N__58651\
        );

    \I__13221\ : InMux
    port map (
            O => \N__58666\,
            I => \N__58648\
        );

    \I__13220\ : InMux
    port map (
            O => \N__58665\,
            I => \N__58645\
        );

    \I__13219\ : InMux
    port map (
            O => \N__58664\,
            I => \N__58642\
        );

    \I__13218\ : InMux
    port map (
            O => \N__58663\,
            I => \N__58639\
        );

    \I__13217\ : LocalMux
    port map (
            O => \N__58660\,
            I => \N__58636\
        );

    \I__13216\ : Span4Mux_v
    port map (
            O => \N__58657\,
            I => \N__58633\
        );

    \I__13215\ : Span4Mux_h
    port map (
            O => \N__58654\,
            I => \N__58630\
        );

    \I__13214\ : Span12Mux_h
    port map (
            O => \N__58651\,
            I => \N__58627\
        );

    \I__13213\ : LocalMux
    port map (
            O => \N__58648\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13212\ : LocalMux
    port map (
            O => \N__58645\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13211\ : LocalMux
    port map (
            O => \N__58642\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13210\ : LocalMux
    port map (
            O => \N__58639\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13209\ : Odrv4
    port map (
            O => \N__58636\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13208\ : Odrv4
    port map (
            O => \N__58633\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13207\ : Odrv4
    port map (
            O => \N__58630\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13206\ : Odrv12
    port map (
            O => \N__58627\,
            I => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\
        );

    \I__13205\ : InMux
    port map (
            O => \N__58610\,
            I => \N__58607\
        );

    \I__13204\ : LocalMux
    port map (
            O => \N__58607\,
            I => \N__58603\
        );

    \I__13203\ : InMux
    port map (
            O => \N__58606\,
            I => \N__58599\
        );

    \I__13202\ : Span4Mux_v
    port map (
            O => \N__58603\,
            I => \N__58596\
        );

    \I__13201\ : InMux
    port map (
            O => \N__58602\,
            I => \N__58593\
        );

    \I__13200\ : LocalMux
    port map (
            O => \N__58599\,
            I => \N__58590\
        );

    \I__13199\ : Span4Mux_h
    port map (
            O => \N__58596\,
            I => \N__58585\
        );

    \I__13198\ : LocalMux
    port map (
            O => \N__58593\,
            I => \N__58585\
        );

    \I__13197\ : Span4Mux_h
    port map (
            O => \N__58590\,
            I => \N__58582\
        );

    \I__13196\ : Span4Mux_h
    port map (
            O => \N__58585\,
            I => \N__58579\
        );

    \I__13195\ : Span4Mux_h
    port map (
            O => \N__58582\,
            I => \N__58576\
        );

    \I__13194\ : Span4Mux_v
    port map (
            O => \N__58579\,
            I => \N__58573\
        );

    \I__13193\ : Span4Mux_v
    port map (
            O => \N__58576\,
            I => \N__58570\
        );

    \I__13192\ : Odrv4
    port map (
            O => \N__58573\,
            I => h_3
        );

    \I__13191\ : Odrv4
    port map (
            O => \N__58570\,
            I => h_3
        );

    \I__13190\ : CascadeMux
    port map (
            O => \N__58565\,
            I => \N__58559\
        );

    \I__13189\ : CascadeMux
    port map (
            O => \N__58564\,
            I => \N__58556\
        );

    \I__13188\ : CascadeMux
    port map (
            O => \N__58563\,
            I => \N__58553\
        );

    \I__13187\ : InMux
    port map (
            O => \N__58562\,
            I => \N__58548\
        );

    \I__13186\ : InMux
    port map (
            O => \N__58559\,
            I => \N__58544\
        );

    \I__13185\ : InMux
    port map (
            O => \N__58556\,
            I => \N__58541\
        );

    \I__13184\ : InMux
    port map (
            O => \N__58553\,
            I => \N__58538\
        );

    \I__13183\ : InMux
    port map (
            O => \N__58552\,
            I => \N__58535\
        );

    \I__13182\ : CascadeMux
    port map (
            O => \N__58551\,
            I => \N__58530\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__58548\,
            I => \N__58527\
        );

    \I__13180\ : CascadeMux
    port map (
            O => \N__58547\,
            I => \N__58521\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__58544\,
            I => \N__58516\
        );

    \I__13178\ : LocalMux
    port map (
            O => \N__58541\,
            I => \N__58516\
        );

    \I__13177\ : LocalMux
    port map (
            O => \N__58538\,
            I => \N__58511\
        );

    \I__13176\ : LocalMux
    port map (
            O => \N__58535\,
            I => \N__58511\
        );

    \I__13175\ : InMux
    port map (
            O => \N__58534\,
            I => \N__58505\
        );

    \I__13174\ : InMux
    port map (
            O => \N__58533\,
            I => \N__58505\
        );

    \I__13173\ : InMux
    port map (
            O => \N__58530\,
            I => \N__58502\
        );

    \I__13172\ : Span4Mux_v
    port map (
            O => \N__58527\,
            I => \N__58499\
        );

    \I__13171\ : InMux
    port map (
            O => \N__58526\,
            I => \N__58491\
        );

    \I__13170\ : InMux
    port map (
            O => \N__58525\,
            I => \N__58488\
        );

    \I__13169\ : InMux
    port map (
            O => \N__58524\,
            I => \N__58485\
        );

    \I__13168\ : InMux
    port map (
            O => \N__58521\,
            I => \N__58482\
        );

    \I__13167\ : Span4Mux_v
    port map (
            O => \N__58516\,
            I => \N__58479\
        );

    \I__13166\ : Span4Mux_h
    port map (
            O => \N__58511\,
            I => \N__58476\
        );

    \I__13165\ : InMux
    port map (
            O => \N__58510\,
            I => \N__58473\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__58505\,
            I => \N__58470\
        );

    \I__13163\ : LocalMux
    port map (
            O => \N__58502\,
            I => \N__58465\
        );

    \I__13162\ : Sp12to4
    port map (
            O => \N__58499\,
            I => \N__58465\
        );

    \I__13161\ : InMux
    port map (
            O => \N__58498\,
            I => \N__58462\
        );

    \I__13160\ : InMux
    port map (
            O => \N__58497\,
            I => \N__58457\
        );

    \I__13159\ : InMux
    port map (
            O => \N__58496\,
            I => \N__58457\
        );

    \I__13158\ : InMux
    port map (
            O => \N__58495\,
            I => \N__58452\
        );

    \I__13157\ : InMux
    port map (
            O => \N__58494\,
            I => \N__58449\
        );

    \I__13156\ : LocalMux
    port map (
            O => \N__58491\,
            I => \N__58444\
        );

    \I__13155\ : LocalMux
    port map (
            O => \N__58488\,
            I => \N__58444\
        );

    \I__13154\ : LocalMux
    port map (
            O => \N__58485\,
            I => \N__58439\
        );

    \I__13153\ : LocalMux
    port map (
            O => \N__58482\,
            I => \N__58439\
        );

    \I__13152\ : Span4Mux_h
    port map (
            O => \N__58479\,
            I => \N__58434\
        );

    \I__13151\ : Span4Mux_v
    port map (
            O => \N__58476\,
            I => \N__58434\
        );

    \I__13150\ : LocalMux
    port map (
            O => \N__58473\,
            I => \N__58431\
        );

    \I__13149\ : Span4Mux_v
    port map (
            O => \N__58470\,
            I => \N__58428\
        );

    \I__13148\ : Span12Mux_h
    port map (
            O => \N__58465\,
            I => \N__58423\
        );

    \I__13147\ : LocalMux
    port map (
            O => \N__58462\,
            I => \N__58423\
        );

    \I__13146\ : LocalMux
    port map (
            O => \N__58457\,
            I => \N__58420\
        );

    \I__13145\ : InMux
    port map (
            O => \N__58456\,
            I => \N__58417\
        );

    \I__13144\ : InMux
    port map (
            O => \N__58455\,
            I => \N__58414\
        );

    \I__13143\ : LocalMux
    port map (
            O => \N__58452\,
            I => \N__58409\
        );

    \I__13142\ : LocalMux
    port map (
            O => \N__58449\,
            I => \N__58409\
        );

    \I__13141\ : Span12Mux_v
    port map (
            O => \N__58444\,
            I => \N__58406\
        );

    \I__13140\ : Span12Mux_v
    port map (
            O => \N__58439\,
            I => \N__58403\
        );

    \I__13139\ : Span4Mux_v
    port map (
            O => \N__58434\,
            I => \N__58396\
        );

    \I__13138\ : Span4Mux_v
    port map (
            O => \N__58431\,
            I => \N__58396\
        );

    \I__13137\ : Span4Mux_h
    port map (
            O => \N__58428\,
            I => \N__58396\
        );

    \I__13136\ : Span12Mux_v
    port map (
            O => \N__58423\,
            I => \N__58393\
        );

    \I__13135\ : Span4Mux_h
    port map (
            O => \N__58420\,
            I => \N__58390\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__58417\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13133\ : LocalMux
    port map (
            O => \N__58414\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13132\ : Odrv4
    port map (
            O => \N__58409\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13131\ : Odrv12
    port map (
            O => \N__58406\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13130\ : Odrv12
    port map (
            O => \N__58403\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13129\ : Odrv4
    port map (
            O => \N__58396\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13128\ : Odrv12
    port map (
            O => \N__58393\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13127\ : Odrv4
    port map (
            O => \N__58390\,
            I => \ALU.a_15_sZ0Z_13\
        );

    \I__13126\ : CascadeMux
    port map (
            O => \N__58373\,
            I => \N__58367\
        );

    \I__13125\ : InMux
    port map (
            O => \N__58372\,
            I => \N__58362\
        );

    \I__13124\ : InMux
    port map (
            O => \N__58371\,
            I => \N__58359\
        );

    \I__13123\ : InMux
    port map (
            O => \N__58370\,
            I => \N__58356\
        );

    \I__13122\ : InMux
    port map (
            O => \N__58367\,
            I => \N__58353\
        );

    \I__13121\ : InMux
    port map (
            O => \N__58366\,
            I => \N__58350\
        );

    \I__13120\ : InMux
    port map (
            O => \N__58365\,
            I => \N__58347\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__58362\,
            I => \N__58344\
        );

    \I__13118\ : LocalMux
    port map (
            O => \N__58359\,
            I => \N__58340\
        );

    \I__13117\ : LocalMux
    port map (
            O => \N__58356\,
            I => \N__58337\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__58353\,
            I => \N__58330\
        );

    \I__13115\ : LocalMux
    port map (
            O => \N__58350\,
            I => \N__58330\
        );

    \I__13114\ : LocalMux
    port map (
            O => \N__58347\,
            I => \N__58330\
        );

    \I__13113\ : Span4Mux_h
    port map (
            O => \N__58344\,
            I => \N__58327\
        );

    \I__13112\ : InMux
    port map (
            O => \N__58343\,
            I => \N__58324\
        );

    \I__13111\ : Span4Mux_h
    port map (
            O => \N__58340\,
            I => \N__58321\
        );

    \I__13110\ : Span4Mux_h
    port map (
            O => \N__58337\,
            I => \N__58318\
        );

    \I__13109\ : Span4Mux_v
    port map (
            O => \N__58330\,
            I => \N__58315\
        );

    \I__13108\ : Span4Mux_h
    port map (
            O => \N__58327\,
            I => \N__58312\
        );

    \I__13107\ : LocalMux
    port map (
            O => \N__58324\,
            I => \ALU.c_RNIO0KOKEZ0Z_10\
        );

    \I__13106\ : Odrv4
    port map (
            O => \N__58321\,
            I => \ALU.c_RNIO0KOKEZ0Z_10\
        );

    \I__13105\ : Odrv4
    port map (
            O => \N__58318\,
            I => \ALU.c_RNIO0KOKEZ0Z_10\
        );

    \I__13104\ : Odrv4
    port map (
            O => \N__58315\,
            I => \ALU.c_RNIO0KOKEZ0Z_10\
        );

    \I__13103\ : Odrv4
    port map (
            O => \N__58312\,
            I => \ALU.c_RNIO0KOKEZ0Z_10\
        );

    \I__13102\ : InMux
    port map (
            O => \N__58301\,
            I => \N__58296\
        );

    \I__13101\ : InMux
    port map (
            O => \N__58300\,
            I => \N__58291\
        );

    \I__13100\ : InMux
    port map (
            O => \N__58299\,
            I => \N__58288\
        );

    \I__13099\ : LocalMux
    port map (
            O => \N__58296\,
            I => \N__58285\
        );

    \I__13098\ : InMux
    port map (
            O => \N__58295\,
            I => \N__58280\
        );

    \I__13097\ : InMux
    port map (
            O => \N__58294\,
            I => \N__58277\
        );

    \I__13096\ : LocalMux
    port map (
            O => \N__58291\,
            I => \N__58274\
        );

    \I__13095\ : LocalMux
    port map (
            O => \N__58288\,
            I => \N__58271\
        );

    \I__13094\ : Span4Mux_v
    port map (
            O => \N__58285\,
            I => \N__58268\
        );

    \I__13093\ : InMux
    port map (
            O => \N__58284\,
            I => \N__58265\
        );

    \I__13092\ : InMux
    port map (
            O => \N__58283\,
            I => \N__58262\
        );

    \I__13091\ : LocalMux
    port map (
            O => \N__58280\,
            I => \N__58255\
        );

    \I__13090\ : LocalMux
    port map (
            O => \N__58277\,
            I => \N__58255\
        );

    \I__13089\ : Span4Mux_h
    port map (
            O => \N__58274\,
            I => \N__58255\
        );

    \I__13088\ : Span4Mux_v
    port map (
            O => \N__58271\,
            I => \N__58250\
        );

    \I__13087\ : Span4Mux_h
    port map (
            O => \N__58268\,
            I => \N__58250\
        );

    \I__13086\ : LocalMux
    port map (
            O => \N__58265\,
            I => \ALU.mult_549_c_RNIE7260OZ0\
        );

    \I__13085\ : LocalMux
    port map (
            O => \N__58262\,
            I => \ALU.mult_549_c_RNIE7260OZ0\
        );

    \I__13084\ : Odrv4
    port map (
            O => \N__58255\,
            I => \ALU.mult_549_c_RNIE7260OZ0\
        );

    \I__13083\ : Odrv4
    port map (
            O => \N__58250\,
            I => \ALU.mult_549_c_RNIE7260OZ0\
        );

    \I__13082\ : CascadeMux
    port map (
            O => \N__58241\,
            I => \N__58238\
        );

    \I__13081\ : InMux
    port map (
            O => \N__58238\,
            I => \N__58235\
        );

    \I__13080\ : LocalMux
    port map (
            O => \N__58235\,
            I => \N__58231\
        );

    \I__13079\ : InMux
    port map (
            O => \N__58234\,
            I => \N__58228\
        );

    \I__13078\ : Span4Mux_v
    port map (
            O => \N__58231\,
            I => \N__58222\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__58228\,
            I => \N__58222\
        );

    \I__13076\ : InMux
    port map (
            O => \N__58227\,
            I => \N__58219\
        );

    \I__13075\ : Span4Mux_v
    port map (
            O => \N__58222\,
            I => \N__58216\
        );

    \I__13074\ : LocalMux
    port map (
            O => \N__58219\,
            I => \N__58213\
        );

    \I__13073\ : Span4Mux_h
    port map (
            O => \N__58216\,
            I => \N__58210\
        );

    \I__13072\ : Span4Mux_v
    port map (
            O => \N__58213\,
            I => \N__58207\
        );

    \I__13071\ : Sp12to4
    port map (
            O => \N__58210\,
            I => \N__58202\
        );

    \I__13070\ : Sp12to4
    port map (
            O => \N__58207\,
            I => \N__58202\
        );

    \I__13069\ : Span12Mux_h
    port map (
            O => \N__58202\,
            I => \N__58199\
        );

    \I__13068\ : Odrv12
    port map (
            O => \N__58199\,
            I => h_10
        );

    \I__13067\ : InMux
    port map (
            O => \N__58196\,
            I => \N__58191\
        );

    \I__13066\ : InMux
    port map (
            O => \N__58195\,
            I => \N__58185\
        );

    \I__13065\ : InMux
    port map (
            O => \N__58194\,
            I => \N__58181\
        );

    \I__13064\ : LocalMux
    port map (
            O => \N__58191\,
            I => \N__58178\
        );

    \I__13063\ : InMux
    port map (
            O => \N__58190\,
            I => \N__58175\
        );

    \I__13062\ : InMux
    port map (
            O => \N__58189\,
            I => \N__58172\
        );

    \I__13061\ : InMux
    port map (
            O => \N__58188\,
            I => \N__58169\
        );

    \I__13060\ : LocalMux
    port map (
            O => \N__58185\,
            I => \N__58166\
        );

    \I__13059\ : InMux
    port map (
            O => \N__58184\,
            I => \N__58162\
        );

    \I__13058\ : LocalMux
    port map (
            O => \N__58181\,
            I => \N__58159\
        );

    \I__13057\ : Span4Mux_v
    port map (
            O => \N__58178\,
            I => \N__58150\
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__58175\,
            I => \N__58150\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__58172\,
            I => \N__58150\
        );

    \I__13054\ : LocalMux
    port map (
            O => \N__58169\,
            I => \N__58150\
        );

    \I__13053\ : Span4Mux_v
    port map (
            O => \N__58166\,
            I => \N__58147\
        );

    \I__13052\ : InMux
    port map (
            O => \N__58165\,
            I => \N__58144\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__58162\,
            I => \N__58139\
        );

    \I__13050\ : Span4Mux_h
    port map (
            O => \N__58159\,
            I => \N__58139\
        );

    \I__13049\ : Span4Mux_v
    port map (
            O => \N__58150\,
            I => \N__58134\
        );

    \I__13048\ : Span4Mux_h
    port map (
            O => \N__58147\,
            I => \N__58134\
        );

    \I__13047\ : LocalMux
    port map (
            O => \N__58144\,
            I => \ALU.c_RNIBN2FN8Z0Z_11\
        );

    \I__13046\ : Odrv4
    port map (
            O => \N__58139\,
            I => \ALU.c_RNIBN2FN8Z0Z_11\
        );

    \I__13045\ : Odrv4
    port map (
            O => \N__58134\,
            I => \ALU.c_RNIBN2FN8Z0Z_11\
        );

    \I__13044\ : CascadeMux
    port map (
            O => \N__58127\,
            I => \N__58123\
        );

    \I__13043\ : CascadeMux
    port map (
            O => \N__58126\,
            I => \N__58120\
        );

    \I__13042\ : InMux
    port map (
            O => \N__58123\,
            I => \N__58115\
        );

    \I__13041\ : InMux
    port map (
            O => \N__58120\,
            I => \N__58112\
        );

    \I__13040\ : InMux
    port map (
            O => \N__58119\,
            I => \N__58105\
        );

    \I__13039\ : InMux
    port map (
            O => \N__58118\,
            I => \N__58102\
        );

    \I__13038\ : LocalMux
    port map (
            O => \N__58115\,
            I => \N__58099\
        );

    \I__13037\ : LocalMux
    port map (
            O => \N__58112\,
            I => \N__58096\
        );

    \I__13036\ : InMux
    port map (
            O => \N__58111\,
            I => \N__58093\
        );

    \I__13035\ : InMux
    port map (
            O => \N__58110\,
            I => \N__58090\
        );

    \I__13034\ : InMux
    port map (
            O => \N__58109\,
            I => \N__58087\
        );

    \I__13033\ : InMux
    port map (
            O => \N__58108\,
            I => \N__58084\
        );

    \I__13032\ : LocalMux
    port map (
            O => \N__58105\,
            I => \N__58081\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__58102\,
            I => \N__58076\
        );

    \I__13030\ : Span4Mux_h
    port map (
            O => \N__58099\,
            I => \N__58076\
        );

    \I__13029\ : Span4Mux_h
    port map (
            O => \N__58096\,
            I => \N__58073\
        );

    \I__13028\ : LocalMux
    port map (
            O => \N__58093\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\
        );

    \I__13027\ : LocalMux
    port map (
            O => \N__58090\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\
        );

    \I__13026\ : LocalMux
    port map (
            O => \N__58087\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\
        );

    \I__13025\ : LocalMux
    port map (
            O => \N__58084\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\
        );

    \I__13024\ : Odrv4
    port map (
            O => \N__58081\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\
        );

    \I__13023\ : Odrv4
    port map (
            O => \N__58076\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\
        );

    \I__13022\ : Odrv4
    port map (
            O => \N__58073\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\
        );

    \I__13021\ : InMux
    port map (
            O => \N__58058\,
            I => \N__58053\
        );

    \I__13020\ : InMux
    port map (
            O => \N__58057\,
            I => \N__58046\
        );

    \I__13019\ : InMux
    port map (
            O => \N__58056\,
            I => \N__58043\
        );

    \I__13018\ : LocalMux
    port map (
            O => \N__58053\,
            I => \N__58040\
        );

    \I__13017\ : InMux
    port map (
            O => \N__58052\,
            I => \N__58037\
        );

    \I__13016\ : InMux
    port map (
            O => \N__58051\,
            I => \N__58034\
        );

    \I__13015\ : InMux
    port map (
            O => \N__58050\,
            I => \N__58031\
        );

    \I__13014\ : InMux
    port map (
            O => \N__58049\,
            I => \N__58028\
        );

    \I__13013\ : LocalMux
    port map (
            O => \N__58046\,
            I => \N__58025\
        );

    \I__13012\ : LocalMux
    port map (
            O => \N__58043\,
            I => \N__58022\
        );

    \I__13011\ : Span4Mux_v
    port map (
            O => \N__58040\,
            I => \N__58019\
        );

    \I__13010\ : LocalMux
    port map (
            O => \N__58037\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0\
        );

    \I__13009\ : LocalMux
    port map (
            O => \N__58034\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0\
        );

    \I__13008\ : LocalMux
    port map (
            O => \N__58031\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0\
        );

    \I__13007\ : LocalMux
    port map (
            O => \N__58028\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0\
        );

    \I__13006\ : Odrv4
    port map (
            O => \N__58025\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0\
        );

    \I__13005\ : Odrv12
    port map (
            O => \N__58022\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0\
        );

    \I__13004\ : Odrv4
    port map (
            O => \N__58019\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0\
        );

    \I__13003\ : CascadeMux
    port map (
            O => \N__58004\,
            I => \N__58001\
        );

    \I__13002\ : InMux
    port map (
            O => \N__58001\,
            I => \N__57998\
        );

    \I__13001\ : LocalMux
    port map (
            O => \N__57998\,
            I => \N__57994\
        );

    \I__13000\ : InMux
    port map (
            O => \N__57997\,
            I => \N__57991\
        );

    \I__12999\ : Span4Mux_v
    port map (
            O => \N__57994\,
            I => \N__57988\
        );

    \I__12998\ : LocalMux
    port map (
            O => \N__57991\,
            I => \N__57985\
        );

    \I__12997\ : Span4Mux_h
    port map (
            O => \N__57988\,
            I => \N__57982\
        );

    \I__12996\ : Span4Mux_v
    port map (
            O => \N__57985\,
            I => \N__57978\
        );

    \I__12995\ : Span4Mux_v
    port map (
            O => \N__57982\,
            I => \N__57975\
        );

    \I__12994\ : InMux
    port map (
            O => \N__57981\,
            I => \N__57972\
        );

    \I__12993\ : Span4Mux_h
    port map (
            O => \N__57978\,
            I => \N__57969\
        );

    \I__12992\ : Sp12to4
    port map (
            O => \N__57975\,
            I => \N__57964\
        );

    \I__12991\ : LocalMux
    port map (
            O => \N__57972\,
            I => \N__57964\
        );

    \I__12990\ : Span4Mux_h
    port map (
            O => \N__57969\,
            I => \N__57961\
        );

    \I__12989\ : Span12Mux_h
    port map (
            O => \N__57964\,
            I => \N__57958\
        );

    \I__12988\ : Span4Mux_v
    port map (
            O => \N__57961\,
            I => \N__57955\
        );

    \I__12987\ : Odrv12
    port map (
            O => \N__57958\,
            I => h_11
        );

    \I__12986\ : Odrv4
    port map (
            O => \N__57955\,
            I => h_11
        );

    \I__12985\ : InMux
    port map (
            O => \N__57950\,
            I => \N__57947\
        );

    \I__12984\ : LocalMux
    port map (
            O => \N__57947\,
            I => \N__57943\
        );

    \I__12983\ : InMux
    port map (
            O => \N__57946\,
            I => \N__57940\
        );

    \I__12982\ : Span4Mux_v
    port map (
            O => \N__57943\,
            I => \N__57935\
        );

    \I__12981\ : LocalMux
    port map (
            O => \N__57940\,
            I => \N__57935\
        );

    \I__12980\ : Span4Mux_v
    port map (
            O => \N__57935\,
            I => \N__57931\
        );

    \I__12979\ : InMux
    port map (
            O => \N__57934\,
            I => \N__57928\
        );

    \I__12978\ : Span4Mux_h
    port map (
            O => \N__57931\,
            I => \N__57925\
        );

    \I__12977\ : LocalMux
    port map (
            O => \N__57928\,
            I => \N__57922\
        );

    \I__12976\ : Span4Mux_h
    port map (
            O => \N__57925\,
            I => \N__57917\
        );

    \I__12975\ : Span4Mux_v
    port map (
            O => \N__57922\,
            I => \N__57917\
        );

    \I__12974\ : Sp12to4
    port map (
            O => \N__57917\,
            I => \N__57914\
        );

    \I__12973\ : Span12Mux_h
    port map (
            O => \N__57914\,
            I => \N__57911\
        );

    \I__12972\ : Odrv12
    port map (
            O => \N__57911\,
            I => h_12
        );

    \I__12971\ : InMux
    port map (
            O => \N__57908\,
            I => \N__57905\
        );

    \I__12970\ : LocalMux
    port map (
            O => \N__57905\,
            I => \N__57902\
        );

    \I__12969\ : Span4Mux_v
    port map (
            O => \N__57902\,
            I => \N__57899\
        );

    \I__12968\ : Span4Mux_h
    port map (
            O => \N__57899\,
            I => \N__57896\
        );

    \I__12967\ : Span4Mux_v
    port map (
            O => \N__57896\,
            I => \N__57893\
        );

    \I__12966\ : Sp12to4
    port map (
            O => \N__57893\,
            I => \N__57888\
        );

    \I__12965\ : InMux
    port map (
            O => \N__57892\,
            I => \N__57885\
        );

    \I__12964\ : InMux
    port map (
            O => \N__57891\,
            I => \N__57882\
        );

    \I__12963\ : Span12Mux_h
    port map (
            O => \N__57888\,
            I => \N__57877\
        );

    \I__12962\ : LocalMux
    port map (
            O => \N__57885\,
            I => \N__57877\
        );

    \I__12961\ : LocalMux
    port map (
            O => \N__57882\,
            I => \N__57872\
        );

    \I__12960\ : Span12Mux_v
    port map (
            O => \N__57877\,
            I => \N__57872\
        );

    \I__12959\ : Odrv12
    port map (
            O => \N__57872\,
            I => h_13
        );

    \I__12958\ : CascadeMux
    port map (
            O => \N__57869\,
            I => \N__57866\
        );

    \I__12957\ : InMux
    port map (
            O => \N__57866\,
            I => \N__57863\
        );

    \I__12956\ : LocalMux
    port map (
            O => \N__57863\,
            I => \N__57860\
        );

    \I__12955\ : Span4Mux_v
    port map (
            O => \N__57860\,
            I => \N__57856\
        );

    \I__12954\ : InMux
    port map (
            O => \N__57859\,
            I => \N__57853\
        );

    \I__12953\ : Span4Mux_h
    port map (
            O => \N__57856\,
            I => \N__57849\
        );

    \I__12952\ : LocalMux
    port map (
            O => \N__57853\,
            I => \N__57846\
        );

    \I__12951\ : InMux
    port map (
            O => \N__57852\,
            I => \N__57843\
        );

    \I__12950\ : Span4Mux_h
    port map (
            O => \N__57849\,
            I => \N__57840\
        );

    \I__12949\ : Span4Mux_v
    port map (
            O => \N__57846\,
            I => \N__57835\
        );

    \I__12948\ : LocalMux
    port map (
            O => \N__57843\,
            I => \N__57835\
        );

    \I__12947\ : Span4Mux_h
    port map (
            O => \N__57840\,
            I => \N__57830\
        );

    \I__12946\ : Span4Mux_h
    port map (
            O => \N__57835\,
            I => \N__57830\
        );

    \I__12945\ : Span4Mux_h
    port map (
            O => \N__57830\,
            I => \N__57827\
        );

    \I__12944\ : Span4Mux_h
    port map (
            O => \N__57827\,
            I => \N__57824\
        );

    \I__12943\ : Odrv4
    port map (
            O => \N__57824\,
            I => h_14
        );

    \I__12942\ : InMux
    port map (
            O => \N__57821\,
            I => \N__57816\
        );

    \I__12941\ : InMux
    port map (
            O => \N__57820\,
            I => \N__57813\
        );

    \I__12940\ : InMux
    port map (
            O => \N__57819\,
            I => \N__57810\
        );

    \I__12939\ : LocalMux
    port map (
            O => \N__57816\,
            I => \N__57805\
        );

    \I__12938\ : LocalMux
    port map (
            O => \N__57813\,
            I => \N__57802\
        );

    \I__12937\ : LocalMux
    port map (
            O => \N__57810\,
            I => \N__57798\
        );

    \I__12936\ : InMux
    port map (
            O => \N__57809\,
            I => \N__57793\
        );

    \I__12935\ : InMux
    port map (
            O => \N__57808\,
            I => \N__57793\
        );

    \I__12934\ : Span4Mux_v
    port map (
            O => \N__57805\,
            I => \N__57788\
        );

    \I__12933\ : Span4Mux_v
    port map (
            O => \N__57802\,
            I => \N__57785\
        );

    \I__12932\ : InMux
    port map (
            O => \N__57801\,
            I => \N__57782\
        );

    \I__12931\ : Span4Mux_h
    port map (
            O => \N__57798\,
            I => \N__57777\
        );

    \I__12930\ : LocalMux
    port map (
            O => \N__57793\,
            I => \N__57777\
        );

    \I__12929\ : InMux
    port map (
            O => \N__57792\,
            I => \N__57774\
        );

    \I__12928\ : InMux
    port map (
            O => \N__57791\,
            I => \N__57771\
        );

    \I__12927\ : Span4Mux_v
    port map (
            O => \N__57788\,
            I => \N__57768\
        );

    \I__12926\ : Sp12to4
    port map (
            O => \N__57785\,
            I => \N__57765\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__57782\,
            I => \N__57762\
        );

    \I__12924\ : Span4Mux_v
    port map (
            O => \N__57777\,
            I => \N__57758\
        );

    \I__12923\ : LocalMux
    port map (
            O => \N__57774\,
            I => \N__57755\
        );

    \I__12922\ : LocalMux
    port map (
            O => \N__57771\,
            I => \N__57752\
        );

    \I__12921\ : Span4Mux_v
    port map (
            O => \N__57768\,
            I => \N__57748\
        );

    \I__12920\ : Span12Mux_h
    port map (
            O => \N__57765\,
            I => \N__57743\
        );

    \I__12919\ : Sp12to4
    port map (
            O => \N__57762\,
            I => \N__57743\
        );

    \I__12918\ : InMux
    port map (
            O => \N__57761\,
            I => \N__57740\
        );

    \I__12917\ : Sp12to4
    port map (
            O => \N__57758\,
            I => \N__57737\
        );

    \I__12916\ : Span4Mux_h
    port map (
            O => \N__57755\,
            I => \N__57732\
        );

    \I__12915\ : Span4Mux_h
    port map (
            O => \N__57752\,
            I => \N__57732\
        );

    \I__12914\ : InMux
    port map (
            O => \N__57751\,
            I => \N__57729\
        );

    \I__12913\ : Span4Mux_h
    port map (
            O => \N__57748\,
            I => \N__57725\
        );

    \I__12912\ : Span12Mux_v
    port map (
            O => \N__57743\,
            I => \N__57722\
        );

    \I__12911\ : LocalMux
    port map (
            O => \N__57740\,
            I => \N__57715\
        );

    \I__12910\ : Span12Mux_h
    port map (
            O => \N__57737\,
            I => \N__57715\
        );

    \I__12909\ : Sp12to4
    port map (
            O => \N__57732\,
            I => \N__57715\
        );

    \I__12908\ : LocalMux
    port map (
            O => \N__57729\,
            I => \N__57712\
        );

    \I__12907\ : InMux
    port map (
            O => \N__57728\,
            I => \N__57709\
        );

    \I__12906\ : Span4Mux_v
    port map (
            O => \N__57725\,
            I => \N__57706\
        );

    \I__12905\ : Span12Mux_h
    port map (
            O => \N__57722\,
            I => \N__57703\
        );

    \I__12904\ : Span12Mux_v
    port map (
            O => \N__57715\,
            I => \N__57700\
        );

    \I__12903\ : Span4Mux_h
    port map (
            O => \N__57712\,
            I => \N__57697\
        );

    \I__12902\ : LocalMux
    port map (
            O => \N__57709\,
            I => \CONTROL.addrstack_1\
        );

    \I__12901\ : Odrv4
    port map (
            O => \N__57706\,
            I => \CONTROL.addrstack_1\
        );

    \I__12900\ : Odrv12
    port map (
            O => \N__57703\,
            I => \CONTROL.addrstack_1\
        );

    \I__12899\ : Odrv12
    port map (
            O => \N__57700\,
            I => \CONTROL.addrstack_1\
        );

    \I__12898\ : Odrv4
    port map (
            O => \N__57697\,
            I => \CONTROL.addrstack_1\
        );

    \I__12897\ : CascadeMux
    port map (
            O => \N__57686\,
            I => \N__57682\
        );

    \I__12896\ : InMux
    port map (
            O => \N__57685\,
            I => \N__57679\
        );

    \I__12895\ : InMux
    port map (
            O => \N__57682\,
            I => \N__57676\
        );

    \I__12894\ : LocalMux
    port map (
            O => \N__57679\,
            I => \N__57672\
        );

    \I__12893\ : LocalMux
    port map (
            O => \N__57676\,
            I => \N__57669\
        );

    \I__12892\ : InMux
    port map (
            O => \N__57675\,
            I => \N__57666\
        );

    \I__12891\ : Span4Mux_h
    port map (
            O => \N__57672\,
            I => \N__57661\
        );

    \I__12890\ : Span4Mux_v
    port map (
            O => \N__57669\,
            I => \N__57661\
        );

    \I__12889\ : LocalMux
    port map (
            O => \N__57666\,
            I => \N__57658\
        );

    \I__12888\ : Span4Mux_v
    port map (
            O => \N__57661\,
            I => \N__57655\
        );

    \I__12887\ : Span12Mux_v
    port map (
            O => \N__57658\,
            I => \N__57652\
        );

    \I__12886\ : Span4Mux_h
    port map (
            O => \N__57655\,
            I => \N__57649\
        );

    \I__12885\ : Span12Mux_h
    port map (
            O => \N__57652\,
            I => \N__57646\
        );

    \I__12884\ : Span4Mux_h
    port map (
            O => \N__57649\,
            I => \N__57643\
        );

    \I__12883\ : Odrv12
    port map (
            O => \N__57646\,
            I => f_12
        );

    \I__12882\ : Odrv4
    port map (
            O => \N__57643\,
            I => f_12
        );

    \I__12881\ : CascadeMux
    port map (
            O => \N__57638\,
            I => \N__57635\
        );

    \I__12880\ : InMux
    port map (
            O => \N__57635\,
            I => \N__57632\
        );

    \I__12879\ : LocalMux
    port map (
            O => \N__57632\,
            I => \N__57628\
        );

    \I__12878\ : InMux
    port map (
            O => \N__57631\,
            I => \N__57625\
        );

    \I__12877\ : Span4Mux_v
    port map (
            O => \N__57628\,
            I => \N__57622\
        );

    \I__12876\ : LocalMux
    port map (
            O => \N__57625\,
            I => \N__57616\
        );

    \I__12875\ : Span4Mux_v
    port map (
            O => \N__57622\,
            I => \N__57616\
        );

    \I__12874\ : InMux
    port map (
            O => \N__57621\,
            I => \N__57613\
        );

    \I__12873\ : Span4Mux_h
    port map (
            O => \N__57616\,
            I => \N__57610\
        );

    \I__12872\ : LocalMux
    port map (
            O => \N__57613\,
            I => \N__57607\
        );

    \I__12871\ : Span4Mux_h
    port map (
            O => \N__57610\,
            I => \N__57604\
        );

    \I__12870\ : Span12Mux_h
    port map (
            O => \N__57607\,
            I => \N__57601\
        );

    \I__12869\ : Span4Mux_h
    port map (
            O => \N__57604\,
            I => \N__57598\
        );

    \I__12868\ : Odrv12
    port map (
            O => \N__57601\,
            I => f_13
        );

    \I__12867\ : Odrv4
    port map (
            O => \N__57598\,
            I => f_13
        );

    \I__12866\ : CascadeMux
    port map (
            O => \N__57593\,
            I => \N__57590\
        );

    \I__12865\ : InMux
    port map (
            O => \N__57590\,
            I => \N__57587\
        );

    \I__12864\ : LocalMux
    port map (
            O => \N__57587\,
            I => \N__57583\
        );

    \I__12863\ : CascadeMux
    port map (
            O => \N__57586\,
            I => \N__57579\
        );

    \I__12862\ : Span4Mux_v
    port map (
            O => \N__57583\,
            I => \N__57576\
        );

    \I__12861\ : InMux
    port map (
            O => \N__57582\,
            I => \N__57573\
        );

    \I__12860\ : InMux
    port map (
            O => \N__57579\,
            I => \N__57570\
        );

    \I__12859\ : Span4Mux_h
    port map (
            O => \N__57576\,
            I => \N__57567\
        );

    \I__12858\ : LocalMux
    port map (
            O => \N__57573\,
            I => \N__57564\
        );

    \I__12857\ : LocalMux
    port map (
            O => \N__57570\,
            I => \N__57561\
        );

    \I__12856\ : Sp12to4
    port map (
            O => \N__57567\,
            I => \N__57558\
        );

    \I__12855\ : Span4Mux_h
    port map (
            O => \N__57564\,
            I => \N__57555\
        );

    \I__12854\ : Span4Mux_v
    port map (
            O => \N__57561\,
            I => \N__57552\
        );

    \I__12853\ : Span12Mux_s9_v
    port map (
            O => \N__57558\,
            I => \N__57549\
        );

    \I__12852\ : Span4Mux_h
    port map (
            O => \N__57555\,
            I => \N__57546\
        );

    \I__12851\ : Span4Mux_h
    port map (
            O => \N__57552\,
            I => \N__57543\
        );

    \I__12850\ : Span12Mux_v
    port map (
            O => \N__57549\,
            I => \N__57540\
        );

    \I__12849\ : Span4Mux_v
    port map (
            O => \N__57546\,
            I => \N__57537\
        );

    \I__12848\ : Span4Mux_v
    port map (
            O => \N__57543\,
            I => \N__57534\
        );

    \I__12847\ : Odrv12
    port map (
            O => \N__57540\,
            I => f_14
        );

    \I__12846\ : Odrv4
    port map (
            O => \N__57537\,
            I => f_14
        );

    \I__12845\ : Odrv4
    port map (
            O => \N__57534\,
            I => f_14
        );

    \I__12844\ : CascadeMux
    port map (
            O => \N__57527\,
            I => \N__57524\
        );

    \I__12843\ : InMux
    port map (
            O => \N__57524\,
            I => \N__57518\
        );

    \I__12842\ : InMux
    port map (
            O => \N__57523\,
            I => \N__57518\
        );

    \I__12841\ : LocalMux
    port map (
            O => \N__57518\,
            I => \N__57515\
        );

    \I__12840\ : Span4Mux_v
    port map (
            O => \N__57515\,
            I => \N__57511\
        );

    \I__12839\ : InMux
    port map (
            O => \N__57514\,
            I => \N__57508\
        );

    \I__12838\ : Odrv4
    port map (
            O => \N__57511\,
            I => \ALU.log_1_14\
        );

    \I__12837\ : LocalMux
    port map (
            O => \N__57508\,
            I => \ALU.log_1_14\
        );

    \I__12836\ : InMux
    port map (
            O => \N__57503\,
            I => \N__57500\
        );

    \I__12835\ : LocalMux
    port map (
            O => \N__57500\,
            I => \N__57497\
        );

    \I__12834\ : Span4Mux_h
    port map (
            O => \N__57497\,
            I => \N__57494\
        );

    \I__12833\ : Span4Mux_h
    port map (
            O => \N__57494\,
            I => \N__57491\
        );

    \I__12832\ : Odrv4
    port map (
            O => \N__57491\,
            I => \ALU.a_15_m0_14\
        );

    \I__12831\ : CascadeMux
    port map (
            O => \N__57488\,
            I => \ALU.addsub_cry_13_c_RNIBVHEA1Z0Z_0_cascade_\
        );

    \I__12830\ : InMux
    port map (
            O => \N__57485\,
            I => \N__57482\
        );

    \I__12829\ : LocalMux
    port map (
            O => \N__57482\,
            I => \ALU.addsub_cry_13_c_RNIBVHEAZ0Z1\
        );

    \I__12828\ : CascadeMux
    port map (
            O => \N__57479\,
            I => \ALU.addsub_cry_13_c_RNIJMTGAZ0Z5_cascade_\
        );

    \I__12827\ : InMux
    port map (
            O => \N__57476\,
            I => \N__57473\
        );

    \I__12826\ : LocalMux
    port map (
            O => \N__57473\,
            I => \N__57470\
        );

    \I__12825\ : Span4Mux_h
    port map (
            O => \N__57470\,
            I => \N__57467\
        );

    \I__12824\ : Span4Mux_h
    port map (
            O => \N__57467\,
            I => \N__57464\
        );

    \I__12823\ : Odrv4
    port map (
            O => \N__57464\,
            I => \ALU.mult_14\
        );

    \I__12822\ : CascadeMux
    port map (
            O => \N__57461\,
            I => \ALU.a_15_ns_rn_0_14_cascade_\
        );

    \I__12821\ : InMux
    port map (
            O => \N__57458\,
            I => \N__57455\
        );

    \I__12820\ : LocalMux
    port map (
            O => \N__57455\,
            I => \N__57451\
        );

    \I__12819\ : InMux
    port map (
            O => \N__57454\,
            I => \N__57448\
        );

    \I__12818\ : Span4Mux_v
    port map (
            O => \N__57451\,
            I => \N__57445\
        );

    \I__12817\ : LocalMux
    port map (
            O => \N__57448\,
            I => \N__57442\
        );

    \I__12816\ : Span4Mux_h
    port map (
            O => \N__57445\,
            I => \N__57439\
        );

    \I__12815\ : Span4Mux_h
    port map (
            O => \N__57442\,
            I => \N__57436\
        );

    \I__12814\ : Span4Mux_h
    port map (
            O => \N__57439\,
            I => \N__57433\
        );

    \I__12813\ : Span4Mux_v
    port map (
            O => \N__57436\,
            I => \N__57430\
        );

    \I__12812\ : Span4Mux_v
    port map (
            O => \N__57433\,
            I => \N__57427\
        );

    \I__12811\ : Odrv4
    port map (
            O => \N__57430\,
            I => \ALU.aZ0Z_14\
        );

    \I__12810\ : Odrv4
    port map (
            O => \N__57427\,
            I => \ALU.aZ0Z_14\
        );

    \I__12809\ : InMux
    port map (
            O => \N__57422\,
            I => \N__57416\
        );

    \I__12808\ : InMux
    port map (
            O => \N__57421\,
            I => \N__57413\
        );

    \I__12807\ : InMux
    port map (
            O => \N__57420\,
            I => \N__57407\
        );

    \I__12806\ : InMux
    port map (
            O => \N__57419\,
            I => \N__57407\
        );

    \I__12805\ : LocalMux
    port map (
            O => \N__57416\,
            I => \N__57400\
        );

    \I__12804\ : LocalMux
    port map (
            O => \N__57413\,
            I => \N__57400\
        );

    \I__12803\ : CascadeMux
    port map (
            O => \N__57412\,
            I => \N__57397\
        );

    \I__12802\ : LocalMux
    port map (
            O => \N__57407\,
            I => \N__57393\
        );

    \I__12801\ : InMux
    port map (
            O => \N__57406\,
            I => \N__57390\
        );

    \I__12800\ : CascadeMux
    port map (
            O => \N__57405\,
            I => \N__57385\
        );

    \I__12799\ : Span4Mux_h
    port map (
            O => \N__57400\,
            I => \N__57379\
        );

    \I__12798\ : InMux
    port map (
            O => \N__57397\,
            I => \N__57373\
        );

    \I__12797\ : InMux
    port map (
            O => \N__57396\,
            I => \N__57373\
        );

    \I__12796\ : Span4Mux_v
    port map (
            O => \N__57393\,
            I => \N__57368\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__57390\,
            I => \N__57365\
        );

    \I__12794\ : InMux
    port map (
            O => \N__57389\,
            I => \N__57360\
        );

    \I__12793\ : InMux
    port map (
            O => \N__57388\,
            I => \N__57360\
        );

    \I__12792\ : InMux
    port map (
            O => \N__57385\,
            I => \N__57355\
        );

    \I__12791\ : InMux
    port map (
            O => \N__57384\,
            I => \N__57355\
        );

    \I__12790\ : CascadeMux
    port map (
            O => \N__57383\,
            I => \N__57352\
        );

    \I__12789\ : InMux
    port map (
            O => \N__57382\,
            I => \N__57346\
        );

    \I__12788\ : Span4Mux_h
    port map (
            O => \N__57379\,
            I => \N__57343\
        );

    \I__12787\ : InMux
    port map (
            O => \N__57378\,
            I => \N__57340\
        );

    \I__12786\ : LocalMux
    port map (
            O => \N__57373\,
            I => \N__57337\
        );

    \I__12785\ : InMux
    port map (
            O => \N__57372\,
            I => \N__57332\
        );

    \I__12784\ : InMux
    port map (
            O => \N__57371\,
            I => \N__57332\
        );

    \I__12783\ : Span4Mux_h
    port map (
            O => \N__57368\,
            I => \N__57329\
        );

    \I__12782\ : Span4Mux_h
    port map (
            O => \N__57365\,
            I => \N__57322\
        );

    \I__12781\ : LocalMux
    port map (
            O => \N__57360\,
            I => \N__57322\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__57355\,
            I => \N__57322\
        );

    \I__12779\ : InMux
    port map (
            O => \N__57352\,
            I => \N__57316\
        );

    \I__12778\ : InMux
    port map (
            O => \N__57351\,
            I => \N__57316\
        );

    \I__12777\ : InMux
    port map (
            O => \N__57350\,
            I => \N__57311\
        );

    \I__12776\ : InMux
    port map (
            O => \N__57349\,
            I => \N__57311\
        );

    \I__12775\ : LocalMux
    port map (
            O => \N__57346\,
            I => \N__57300\
        );

    \I__12774\ : Span4Mux_v
    port map (
            O => \N__57343\,
            I => \N__57300\
        );

    \I__12773\ : LocalMux
    port map (
            O => \N__57340\,
            I => \N__57300\
        );

    \I__12772\ : Span4Mux_v
    port map (
            O => \N__57337\,
            I => \N__57300\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__57332\,
            I => \N__57300\
        );

    \I__12770\ : Span4Mux_v
    port map (
            O => \N__57329\,
            I => \N__57295\
        );

    \I__12769\ : Span4Mux_h
    port map (
            O => \N__57322\,
            I => \N__57295\
        );

    \I__12768\ : InMux
    port map (
            O => \N__57321\,
            I => \N__57292\
        );

    \I__12767\ : LocalMux
    port map (
            O => \N__57316\,
            I => \N__57285\
        );

    \I__12766\ : LocalMux
    port map (
            O => \N__57311\,
            I => \N__57285\
        );

    \I__12765\ : Span4Mux_v
    port map (
            O => \N__57300\,
            I => \N__57285\
        );

    \I__12764\ : Span4Mux_h
    port map (
            O => \N__57295\,
            I => \N__57282\
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__57292\,
            I => \N__57279\
        );

    \I__12762\ : Span4Mux_h
    port map (
            O => \N__57285\,
            I => \N__57276\
        );

    \I__12761\ : Span4Mux_h
    port map (
            O => \N__57282\,
            I => \N__57273\
        );

    \I__12760\ : Sp12to4
    port map (
            O => \N__57279\,
            I => \N__57270\
        );

    \I__12759\ : Span4Mux_h
    port map (
            O => \N__57276\,
            I => \N__57267\
        );

    \I__12758\ : Sp12to4
    port map (
            O => \N__57273\,
            I => \N__57264\
        );

    \I__12757\ : Span12Mux_s11_v
    port map (
            O => \N__57270\,
            I => \N__57261\
        );

    \I__12756\ : Span4Mux_h
    port map (
            O => \N__57267\,
            I => \N__57258\
        );

    \I__12755\ : Span12Mux_s11_v
    port map (
            O => \N__57264\,
            I => \N__57255\
        );

    \I__12754\ : Odrv12
    port map (
            O => \N__57261\,
            I => \ALU.a_15_sZ0Z_3\
        );

    \I__12753\ : Odrv4
    port map (
            O => \N__57258\,
            I => \ALU.a_15_sZ0Z_3\
        );

    \I__12752\ : Odrv12
    port map (
            O => \N__57255\,
            I => \ALU.a_15_sZ0Z_3\
        );

    \I__12751\ : InMux
    port map (
            O => \N__57248\,
            I => \N__57245\
        );

    \I__12750\ : LocalMux
    port map (
            O => \N__57245\,
            I => \ALU.log_1_3\
        );

    \I__12749\ : InMux
    port map (
            O => \N__57242\,
            I => \N__57239\
        );

    \I__12748\ : LocalMux
    port map (
            O => \N__57239\,
            I => \N__57235\
        );

    \I__12747\ : InMux
    port map (
            O => \N__57238\,
            I => \N__57232\
        );

    \I__12746\ : Span4Mux_h
    port map (
            O => \N__57235\,
            I => \N__57228\
        );

    \I__12745\ : LocalMux
    port map (
            O => \N__57232\,
            I => \N__57224\
        );

    \I__12744\ : InMux
    port map (
            O => \N__57231\,
            I => \N__57221\
        );

    \I__12743\ : Span4Mux_v
    port map (
            O => \N__57228\,
            I => \N__57218\
        );

    \I__12742\ : InMux
    port map (
            O => \N__57227\,
            I => \N__57215\
        );

    \I__12741\ : Span4Mux_v
    port map (
            O => \N__57224\,
            I => \N__57212\
        );

    \I__12740\ : LocalMux
    port map (
            O => \N__57221\,
            I => \N__57209\
        );

    \I__12739\ : Span4Mux_h
    port map (
            O => \N__57218\,
            I => \N__57204\
        );

    \I__12738\ : LocalMux
    port map (
            O => \N__57215\,
            I => \N__57204\
        );

    \I__12737\ : Span4Mux_v
    port map (
            O => \N__57212\,
            I => \N__57199\
        );

    \I__12736\ : Span4Mux_h
    port map (
            O => \N__57209\,
            I => \N__57199\
        );

    \I__12735\ : Span4Mux_h
    port map (
            O => \N__57204\,
            I => \N__57196\
        );

    \I__12734\ : Span4Mux_v
    port map (
            O => \N__57199\,
            I => \N__57193\
        );

    \I__12733\ : Span4Mux_h
    port map (
            O => \N__57196\,
            I => \N__57190\
        );

    \I__12732\ : Odrv4
    port map (
            O => \N__57193\,
            I => \ALU.lshift62_2\
        );

    \I__12731\ : Odrv4
    port map (
            O => \N__57190\,
            I => \ALU.lshift62_2\
        );

    \I__12730\ : InMux
    port map (
            O => \N__57185\,
            I => \N__57182\
        );

    \I__12729\ : LocalMux
    port map (
            O => \N__57182\,
            I => \N__57179\
        );

    \I__12728\ : Odrv12
    port map (
            O => \N__57179\,
            I => \ALU.mult_558_c_RNIB3E8DCZ0\
        );

    \I__12727\ : CascadeMux
    port map (
            O => \N__57176\,
            I => \ALU.a_15_d_ns_1_13_cascade_\
        );

    \I__12726\ : CascadeMux
    port map (
            O => \N__57173\,
            I => \ALU.mult_558_c_RNIB75F9GZ0_cascade_\
        );

    \I__12725\ : InMux
    port map (
            O => \N__57170\,
            I => \N__57167\
        );

    \I__12724\ : LocalMux
    port map (
            O => \N__57167\,
            I => \N__57163\
        );

    \I__12723\ : InMux
    port map (
            O => \N__57166\,
            I => \N__57160\
        );

    \I__12722\ : Span4Mux_v
    port map (
            O => \N__57163\,
            I => \N__57157\
        );

    \I__12721\ : LocalMux
    port map (
            O => \N__57160\,
            I => \N__57154\
        );

    \I__12720\ : Span4Mux_h
    port map (
            O => \N__57157\,
            I => \N__57151\
        );

    \I__12719\ : Span4Mux_v
    port map (
            O => \N__57154\,
            I => \N__57148\
        );

    \I__12718\ : Span4Mux_v
    port map (
            O => \N__57151\,
            I => \N__57145\
        );

    \I__12717\ : Sp12to4
    port map (
            O => \N__57148\,
            I => \N__57142\
        );

    \I__12716\ : Sp12to4
    port map (
            O => \N__57145\,
            I => \N__57137\
        );

    \I__12715\ : Span12Mux_h
    port map (
            O => \N__57142\,
            I => \N__57137\
        );

    \I__12714\ : Odrv12
    port map (
            O => \N__57137\,
            I => \ALU.aZ0Z_13\
        );

    \I__12713\ : InMux
    port map (
            O => \N__57134\,
            I => \N__57131\
        );

    \I__12712\ : LocalMux
    port map (
            O => \N__57131\,
            I => \N__57128\
        );

    \I__12711\ : Span4Mux_v
    port map (
            O => \N__57128\,
            I => \N__57125\
        );

    \I__12710\ : Odrv4
    port map (
            O => \N__57125\,
            I => \ALU.d_RNIJ7J1M5_0Z0Z_2\
        );

    \I__12709\ : CascadeMux
    port map (
            O => \N__57122\,
            I => \N__57118\
        );

    \I__12708\ : InMux
    port map (
            O => \N__57121\,
            I => \N__57113\
        );

    \I__12707\ : InMux
    port map (
            O => \N__57118\,
            I => \N__57113\
        );

    \I__12706\ : LocalMux
    port map (
            O => \N__57113\,
            I => \ALU.a_15_m3_d_sZ0Z_8\
        );

    \I__12705\ : InMux
    port map (
            O => \N__57110\,
            I => \N__57104\
        );

    \I__12704\ : InMux
    port map (
            O => \N__57109\,
            I => \N__57104\
        );

    \I__12703\ : LocalMux
    port map (
            O => \N__57104\,
            I => \N__57101\
        );

    \I__12702\ : Span4Mux_v
    port map (
            O => \N__57101\,
            I => \N__57098\
        );

    \I__12701\ : Span4Mux_v
    port map (
            O => \N__57098\,
            I => \N__57095\
        );

    \I__12700\ : Sp12to4
    port map (
            O => \N__57095\,
            I => \N__57091\
        );

    \I__12699\ : InMux
    port map (
            O => \N__57094\,
            I => \N__57088\
        );

    \I__12698\ : Span12Mux_h
    port map (
            O => \N__57091\,
            I => \N__57085\
        );

    \I__12697\ : LocalMux
    port map (
            O => \N__57088\,
            I => \N__57082\
        );

    \I__12696\ : Odrv12
    port map (
            O => \N__57085\,
            I => bus_0_8
        );

    \I__12695\ : Odrv4
    port map (
            O => \N__57082\,
            I => bus_0_8
        );

    \I__12694\ : CascadeMux
    port map (
            O => \N__57077\,
            I => \ALU.a_15_m3_d_sZ0Z_8_cascade_\
        );

    \I__12693\ : InMux
    port map (
            O => \N__57074\,
            I => \N__57068\
        );

    \I__12692\ : InMux
    port map (
            O => \N__57073\,
            I => \N__57068\
        );

    \I__12691\ : LocalMux
    port map (
            O => \N__57068\,
            I => \ALU.d_RNI12L8C5Z0Z_2\
        );

    \I__12690\ : InMux
    port map (
            O => \N__57065\,
            I => \N__57062\
        );

    \I__12689\ : LocalMux
    port map (
            O => \N__57062\,
            I => \N__57059\
        );

    \I__12688\ : Span4Mux_v
    port map (
            O => \N__57059\,
            I => \N__57056\
        );

    \I__12687\ : Odrv4
    port map (
            O => \N__57056\,
            I => \ALU.d_RNIJ7J1M5Z0Z_2\
        );

    \I__12686\ : InMux
    port map (
            O => \N__57053\,
            I => \N__57050\
        );

    \I__12685\ : LocalMux
    port map (
            O => \N__57050\,
            I => \N__57047\
        );

    \I__12684\ : Span4Mux_h
    port map (
            O => \N__57047\,
            I => \N__57043\
        );

    \I__12683\ : InMux
    port map (
            O => \N__57046\,
            I => \N__57040\
        );

    \I__12682\ : Span4Mux_h
    port map (
            O => \N__57043\,
            I => \N__57034\
        );

    \I__12681\ : LocalMux
    port map (
            O => \N__57040\,
            I => \N__57034\
        );

    \I__12680\ : InMux
    port map (
            O => \N__57039\,
            I => \N__57025\
        );

    \I__12679\ : Span4Mux_v
    port map (
            O => \N__57034\,
            I => \N__57021\
        );

    \I__12678\ : InMux
    port map (
            O => \N__57033\,
            I => \N__57016\
        );

    \I__12677\ : InMux
    port map (
            O => \N__57032\,
            I => \N__57016\
        );

    \I__12676\ : InMux
    port map (
            O => \N__57031\,
            I => \N__57012\
        );

    \I__12675\ : CascadeMux
    port map (
            O => \N__57030\,
            I => \N__57009\
        );

    \I__12674\ : CascadeMux
    port map (
            O => \N__57029\,
            I => \N__57006\
        );

    \I__12673\ : CascadeMux
    port map (
            O => \N__57028\,
            I => \N__57003\
        );

    \I__12672\ : LocalMux
    port map (
            O => \N__57025\,
            I => \N__57000\
        );

    \I__12671\ : CascadeMux
    port map (
            O => \N__57024\,
            I => \N__56997\
        );

    \I__12670\ : Span4Mux_v
    port map (
            O => \N__57021\,
            I => \N__56994\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__57016\,
            I => \N__56991\
        );

    \I__12668\ : InMux
    port map (
            O => \N__57015\,
            I => \N__56988\
        );

    \I__12667\ : LocalMux
    port map (
            O => \N__57012\,
            I => \N__56984\
        );

    \I__12666\ : InMux
    port map (
            O => \N__57009\,
            I => \N__56977\
        );

    \I__12665\ : InMux
    port map (
            O => \N__57006\,
            I => \N__56977\
        );

    \I__12664\ : InMux
    port map (
            O => \N__57003\,
            I => \N__56977\
        );

    \I__12663\ : Span4Mux_h
    port map (
            O => \N__57000\,
            I => \N__56974\
        );

    \I__12662\ : InMux
    port map (
            O => \N__56997\,
            I => \N__56971\
        );

    \I__12661\ : Span4Mux_h
    port map (
            O => \N__56994\,
            I => \N__56966\
        );

    \I__12660\ : Span4Mux_v
    port map (
            O => \N__56991\,
            I => \N__56966\
        );

    \I__12659\ : LocalMux
    port map (
            O => \N__56988\,
            I => \N__56963\
        );

    \I__12658\ : InMux
    port map (
            O => \N__56987\,
            I => \N__56960\
        );

    \I__12657\ : Span4Mux_h
    port map (
            O => \N__56984\,
            I => \N__56955\
        );

    \I__12656\ : LocalMux
    port map (
            O => \N__56977\,
            I => \N__56955\
        );

    \I__12655\ : Odrv4
    port map (
            O => \N__56974\,
            I => \ALU.status_19_10\
        );

    \I__12654\ : LocalMux
    port map (
            O => \N__56971\,
            I => \ALU.status_19_10\
        );

    \I__12653\ : Odrv4
    port map (
            O => \N__56966\,
            I => \ALU.status_19_10\
        );

    \I__12652\ : Odrv12
    port map (
            O => \N__56963\,
            I => \ALU.status_19_10\
        );

    \I__12651\ : LocalMux
    port map (
            O => \N__56960\,
            I => \ALU.status_19_10\
        );

    \I__12650\ : Odrv4
    port map (
            O => \N__56955\,
            I => \ALU.status_19_10\
        );

    \I__12649\ : CascadeMux
    port map (
            O => \N__56942\,
            I => \N__56939\
        );

    \I__12648\ : InMux
    port map (
            O => \N__56939\,
            I => \N__56936\
        );

    \I__12647\ : LocalMux
    port map (
            O => \N__56936\,
            I => \ALU.aluOut_i_11\
        );

    \I__12646\ : InMux
    port map (
            O => \N__56933\,
            I => \N__56930\
        );

    \I__12645\ : LocalMux
    port map (
            O => \N__56930\,
            I => \N__56925\
        );

    \I__12644\ : InMux
    port map (
            O => \N__56929\,
            I => \N__56920\
        );

    \I__12643\ : InMux
    port map (
            O => \N__56928\,
            I => \N__56920\
        );

    \I__12642\ : Span4Mux_h
    port map (
            O => \N__56925\,
            I => \N__56917\
        );

    \I__12641\ : LocalMux
    port map (
            O => \N__56920\,
            I => \N__56914\
        );

    \I__12640\ : Span4Mux_h
    port map (
            O => \N__56917\,
            I => \N__56911\
        );

    \I__12639\ : Span4Mux_v
    port map (
            O => \N__56914\,
            I => \N__56906\
        );

    \I__12638\ : Span4Mux_h
    port map (
            O => \N__56911\,
            I => \N__56901\
        );

    \I__12637\ : InMux
    port map (
            O => \N__56910\,
            I => \N__56895\
        );

    \I__12636\ : InMux
    port map (
            O => \N__56909\,
            I => \N__56895\
        );

    \I__12635\ : Span4Mux_h
    port map (
            O => \N__56906\,
            I => \N__56892\
        );

    \I__12634\ : InMux
    port map (
            O => \N__56905\,
            I => \N__56889\
        );

    \I__12633\ : InMux
    port map (
            O => \N__56904\,
            I => \N__56886\
        );

    \I__12632\ : Span4Mux_h
    port map (
            O => \N__56901\,
            I => \N__56883\
        );

    \I__12631\ : InMux
    port map (
            O => \N__56900\,
            I => \N__56880\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__56895\,
            I => \N__56877\
        );

    \I__12629\ : Span4Mux_h
    port map (
            O => \N__56892\,
            I => \N__56870\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__56889\,
            I => \N__56870\
        );

    \I__12627\ : LocalMux
    port map (
            O => \N__56886\,
            I => \N__56870\
        );

    \I__12626\ : Span4Mux_v
    port map (
            O => \N__56883\,
            I => \N__56865\
        );

    \I__12625\ : LocalMux
    port map (
            O => \N__56880\,
            I => \N__56865\
        );

    \I__12624\ : Span12Mux_v
    port map (
            O => \N__56877\,
            I => \N__56862\
        );

    \I__12623\ : Span4Mux_h
    port map (
            O => \N__56870\,
            I => \N__56859\
        );

    \I__12622\ : Odrv4
    port map (
            O => \N__56865\,
            I => \ALU.N_126\
        );

    \I__12621\ : Odrv12
    port map (
            O => \N__56862\,
            I => \ALU.N_126\
        );

    \I__12620\ : Odrv4
    port map (
            O => \N__56859\,
            I => \ALU.N_126\
        );

    \I__12619\ : CascadeMux
    port map (
            O => \N__56852\,
            I => \N__56849\
        );

    \I__12618\ : InMux
    port map (
            O => \N__56849\,
            I => \N__56846\
        );

    \I__12617\ : LocalMux
    port map (
            O => \N__56846\,
            I => \ALU.aluOut_i_12\
        );

    \I__12616\ : CascadeMux
    port map (
            O => \N__56843\,
            I => \N__56840\
        );

    \I__12615\ : InMux
    port map (
            O => \N__56840\,
            I => \N__56836\
        );

    \I__12614\ : CascadeMux
    port map (
            O => \N__56839\,
            I => \N__56833\
        );

    \I__12613\ : LocalMux
    port map (
            O => \N__56836\,
            I => \N__56830\
        );

    \I__12612\ : InMux
    port map (
            O => \N__56833\,
            I => \N__56825\
        );

    \I__12611\ : Span4Mux_v
    port map (
            O => \N__56830\,
            I => \N__56820\
        );

    \I__12610\ : InMux
    port map (
            O => \N__56829\,
            I => \N__56815\
        );

    \I__12609\ : InMux
    port map (
            O => \N__56828\,
            I => \N__56815\
        );

    \I__12608\ : LocalMux
    port map (
            O => \N__56825\,
            I => \N__56812\
        );

    \I__12607\ : CascadeMux
    port map (
            O => \N__56824\,
            I => \N__56809\
        );

    \I__12606\ : CascadeMux
    port map (
            O => \N__56823\,
            I => \N__56806\
        );

    \I__12605\ : Span4Mux_h
    port map (
            O => \N__56820\,
            I => \N__56799\
        );

    \I__12604\ : LocalMux
    port map (
            O => \N__56815\,
            I => \N__56799\
        );

    \I__12603\ : Span4Mux_v
    port map (
            O => \N__56812\,
            I => \N__56796\
        );

    \I__12602\ : InMux
    port map (
            O => \N__56809\,
            I => \N__56793\
        );

    \I__12601\ : InMux
    port map (
            O => \N__56806\,
            I => \N__56788\
        );

    \I__12600\ : InMux
    port map (
            O => \N__56805\,
            I => \N__56788\
        );

    \I__12599\ : CascadeMux
    port map (
            O => \N__56804\,
            I => \N__56784\
        );

    \I__12598\ : Span4Mux_h
    port map (
            O => \N__56799\,
            I => \N__56781\
        );

    \I__12597\ : Span4Mux_h
    port map (
            O => \N__56796\,
            I => \N__56778\
        );

    \I__12596\ : LocalMux
    port map (
            O => \N__56793\,
            I => \N__56773\
        );

    \I__12595\ : LocalMux
    port map (
            O => \N__56788\,
            I => \N__56773\
        );

    \I__12594\ : InMux
    port map (
            O => \N__56787\,
            I => \N__56768\
        );

    \I__12593\ : InMux
    port map (
            O => \N__56784\,
            I => \N__56768\
        );

    \I__12592\ : Odrv4
    port map (
            O => \N__56781\,
            I => \ALU.N_125\
        );

    \I__12591\ : Odrv4
    port map (
            O => \N__56778\,
            I => \ALU.N_125\
        );

    \I__12590\ : Odrv12
    port map (
            O => \N__56773\,
            I => \ALU.N_125\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__56768\,
            I => \ALU.N_125\
        );

    \I__12588\ : InMux
    port map (
            O => \N__56759\,
            I => \N__56756\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__56756\,
            I => \ALU.aluOut_i_13\
        );

    \I__12586\ : InMux
    port map (
            O => \N__56753\,
            I => \N__56750\
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__56750\,
            I => \N__56745\
        );

    \I__12584\ : InMux
    port map (
            O => \N__56749\,
            I => \N__56742\
        );

    \I__12583\ : CascadeMux
    port map (
            O => \N__56748\,
            I => \N__56738\
        );

    \I__12582\ : Span4Mux_v
    port map (
            O => \N__56745\,
            I => \N__56734\
        );

    \I__12581\ : LocalMux
    port map (
            O => \N__56742\,
            I => \N__56731\
        );

    \I__12580\ : InMux
    port map (
            O => \N__56741\,
            I => \N__56728\
        );

    \I__12579\ : InMux
    port map (
            O => \N__56738\,
            I => \N__56723\
        );

    \I__12578\ : InMux
    port map (
            O => \N__56737\,
            I => \N__56723\
        );

    \I__12577\ : Span4Mux_h
    port map (
            O => \N__56734\,
            I => \N__56720\
        );

    \I__12576\ : Span4Mux_h
    port map (
            O => \N__56731\,
            I => \N__56713\
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__56728\,
            I => \N__56713\
        );

    \I__12574\ : LocalMux
    port map (
            O => \N__56723\,
            I => \N__56710\
        );

    \I__12573\ : Sp12to4
    port map (
            O => \N__56720\,
            I => \N__56707\
        );

    \I__12572\ : InMux
    port map (
            O => \N__56719\,
            I => \N__56702\
        );

    \I__12571\ : InMux
    port map (
            O => \N__56718\,
            I => \N__56702\
        );

    \I__12570\ : Span4Mux_v
    port map (
            O => \N__56713\,
            I => \N__56699\
        );

    \I__12569\ : Span4Mux_h
    port map (
            O => \N__56710\,
            I => \N__56696\
        );

    \I__12568\ : Span12Mux_v
    port map (
            O => \N__56707\,
            I => \N__56693\
        );

    \I__12567\ : LocalMux
    port map (
            O => \N__56702\,
            I => \N__56688\
        );

    \I__12566\ : Span4Mux_v
    port map (
            O => \N__56699\,
            I => \N__56688\
        );

    \I__12565\ : Span4Mux_h
    port map (
            O => \N__56696\,
            I => \N__56685\
        );

    \I__12564\ : Odrv12
    port map (
            O => \N__56693\,
            I => \ALU.status_19_13\
        );

    \I__12563\ : Odrv4
    port map (
            O => \N__56688\,
            I => \ALU.status_19_13\
        );

    \I__12562\ : Odrv4
    port map (
            O => \N__56685\,
            I => \ALU.status_19_13\
        );

    \I__12561\ : CascadeMux
    port map (
            O => \N__56678\,
            I => \N__56675\
        );

    \I__12560\ : InMux
    port map (
            O => \N__56675\,
            I => \N__56672\
        );

    \I__12559\ : LocalMux
    port map (
            O => \N__56672\,
            I => \ALU.aluOut_i_14\
        );

    \I__12558\ : CascadeMux
    port map (
            O => \N__56669\,
            I => \N__56666\
        );

    \I__12557\ : InMux
    port map (
            O => \N__56666\,
            I => \N__56663\
        );

    \I__12556\ : LocalMux
    port map (
            O => \N__56663\,
            I => \ALU.aluOut_i_15\
        );

    \I__12555\ : InMux
    port map (
            O => \N__56660\,
            I => \bfn_23_9_0_\
        );

    \I__12554\ : InMux
    port map (
            O => \N__56657\,
            I => \N__56651\
        );

    \I__12553\ : InMux
    port map (
            O => \N__56656\,
            I => \N__56651\
        );

    \I__12552\ : LocalMux
    port map (
            O => \N__56651\,
            I => \N__56648\
        );

    \I__12551\ : Span4Mux_v
    port map (
            O => \N__56648\,
            I => \N__56644\
        );

    \I__12550\ : CascadeMux
    port map (
            O => \N__56647\,
            I => \N__56641\
        );

    \I__12549\ : Span4Mux_h
    port map (
            O => \N__56644\,
            I => \N__56638\
        );

    \I__12548\ : InMux
    port map (
            O => \N__56641\,
            I => \N__56635\
        );

    \I__12547\ : Sp12to4
    port map (
            O => \N__56638\,
            I => \N__56632\
        );

    \I__12546\ : LocalMux
    port map (
            O => \N__56635\,
            I => \aluStatus_5\
        );

    \I__12545\ : Odrv12
    port map (
            O => \N__56632\,
            I => \aluStatus_5\
        );

    \I__12544\ : CascadeMux
    port map (
            O => \N__56627\,
            I => \N__56624\
        );

    \I__12543\ : InMux
    port map (
            O => \N__56624\,
            I => \N__56618\
        );

    \I__12542\ : CascadeMux
    port map (
            O => \N__56623\,
            I => \N__56615\
        );

    \I__12541\ : InMux
    port map (
            O => \N__56622\,
            I => \N__56610\
        );

    \I__12540\ : InMux
    port map (
            O => \N__56621\,
            I => \N__56610\
        );

    \I__12539\ : LocalMux
    port map (
            O => \N__56618\,
            I => \N__56607\
        );

    \I__12538\ : InMux
    port map (
            O => \N__56615\,
            I => \N__56604\
        );

    \I__12537\ : LocalMux
    port map (
            O => \N__56610\,
            I => \N__56600\
        );

    \I__12536\ : Span4Mux_h
    port map (
            O => \N__56607\,
            I => \N__56595\
        );

    \I__12535\ : LocalMux
    port map (
            O => \N__56604\,
            I => \N__56595\
        );

    \I__12534\ : CEMux
    port map (
            O => \N__56603\,
            I => \N__56592\
        );

    \I__12533\ : Span4Mux_h
    port map (
            O => \N__56600\,
            I => \N__56589\
        );

    \I__12532\ : Span4Mux_v
    port map (
            O => \N__56595\,
            I => \N__56586\
        );

    \I__12531\ : LocalMux
    port map (
            O => \N__56592\,
            I => \N__56583\
        );

    \I__12530\ : Span4Mux_h
    port map (
            O => \N__56589\,
            I => \N__56580\
        );

    \I__12529\ : Span4Mux_v
    port map (
            O => \N__56586\,
            I => \N__56577\
        );

    \I__12528\ : Span4Mux_v
    port map (
            O => \N__56583\,
            I => \N__56574\
        );

    \I__12527\ : Sp12to4
    port map (
            O => \N__56580\,
            I => \N__56570\
        );

    \I__12526\ : Span4Mux_h
    port map (
            O => \N__56577\,
            I => \N__56567\
        );

    \I__12525\ : Span4Mux_v
    port map (
            O => \N__56574\,
            I => \N__56564\
        );

    \I__12524\ : InMux
    port map (
            O => \N__56573\,
            I => \N__56561\
        );

    \I__12523\ : Span12Mux_s8_v
    port map (
            O => \N__56570\,
            I => \N__56558\
        );

    \I__12522\ : Span4Mux_h
    port map (
            O => \N__56567\,
            I => \N__56555\
        );

    \I__12521\ : Span4Mux_h
    port map (
            O => \N__56564\,
            I => \N__56552\
        );

    \I__12520\ : LocalMux
    port map (
            O => \N__56561\,
            I => \ALU.un1_a41_0\
        );

    \I__12519\ : Odrv12
    port map (
            O => \N__56558\,
            I => \ALU.un1_a41_0\
        );

    \I__12518\ : Odrv4
    port map (
            O => \N__56555\,
            I => \ALU.un1_a41_0\
        );

    \I__12517\ : Odrv4
    port map (
            O => \N__56552\,
            I => \ALU.un1_a41_0\
        );

    \I__12516\ : InMux
    port map (
            O => \N__56543\,
            I => \N__56539\
        );

    \I__12515\ : CascadeMux
    port map (
            O => \N__56542\,
            I => \N__56536\
        );

    \I__12514\ : LocalMux
    port map (
            O => \N__56539\,
            I => \N__56533\
        );

    \I__12513\ : InMux
    port map (
            O => \N__56536\,
            I => \N__56529\
        );

    \I__12512\ : Span4Mux_h
    port map (
            O => \N__56533\,
            I => \N__56526\
        );

    \I__12511\ : InMux
    port map (
            O => \N__56532\,
            I => \N__56523\
        );

    \I__12510\ : LocalMux
    port map (
            O => \N__56529\,
            I => \N__56520\
        );

    \I__12509\ : Span4Mux_h
    port map (
            O => \N__56526\,
            I => \N__56517\
        );

    \I__12508\ : LocalMux
    port map (
            O => \N__56523\,
            I => \N__56514\
        );

    \I__12507\ : Span4Mux_v
    port map (
            O => \N__56520\,
            I => \N__56511\
        );

    \I__12506\ : Span4Mux_v
    port map (
            O => \N__56517\,
            I => \N__56506\
        );

    \I__12505\ : Span4Mux_v
    port map (
            O => \N__56514\,
            I => \N__56506\
        );

    \I__12504\ : Sp12to4
    port map (
            O => \N__56511\,
            I => \N__56503\
        );

    \I__12503\ : Sp12to4
    port map (
            O => \N__56506\,
            I => \N__56500\
        );

    \I__12502\ : Span12Mux_h
    port map (
            O => \N__56503\,
            I => \N__56495\
        );

    \I__12501\ : Span12Mux_h
    port map (
            O => \N__56500\,
            I => \N__56495\
        );

    \I__12500\ : Odrv12
    port map (
            O => \N__56495\,
            I => \ALU.aZ0Z32\
        );

    \I__12499\ : InMux
    port map (
            O => \N__56492\,
            I => \N__56487\
        );

    \I__12498\ : InMux
    port map (
            O => \N__56491\,
            I => \N__56482\
        );

    \I__12497\ : InMux
    port map (
            O => \N__56490\,
            I => \N__56482\
        );

    \I__12496\ : LocalMux
    port map (
            O => \N__56487\,
            I => \N__56479\
        );

    \I__12495\ : LocalMux
    port map (
            O => \N__56482\,
            I => \ALU.N_866\
        );

    \I__12494\ : Odrv12
    port map (
            O => \N__56479\,
            I => \ALU.N_866\
        );

    \I__12493\ : InMux
    port map (
            O => \N__56474\,
            I => \N__56469\
        );

    \I__12492\ : InMux
    port map (
            O => \N__56473\,
            I => \N__56466\
        );

    \I__12491\ : CascadeMux
    port map (
            O => \N__56472\,
            I => \N__56462\
        );

    \I__12490\ : LocalMux
    port map (
            O => \N__56469\,
            I => \N__56459\
        );

    \I__12489\ : LocalMux
    port map (
            O => \N__56466\,
            I => \N__56456\
        );

    \I__12488\ : InMux
    port map (
            O => \N__56465\,
            I => \N__56453\
        );

    \I__12487\ : InMux
    port map (
            O => \N__56462\,
            I => \N__56450\
        );

    \I__12486\ : Span4Mux_h
    port map (
            O => \N__56459\,
            I => \N__56445\
        );

    \I__12485\ : Span4Mux_h
    port map (
            O => \N__56456\,
            I => \N__56445\
        );

    \I__12484\ : LocalMux
    port map (
            O => \N__56453\,
            I => \N__56442\
        );

    \I__12483\ : LocalMux
    port map (
            O => \N__56450\,
            I => \N__56439\
        );

    \I__12482\ : Sp12to4
    port map (
            O => \N__56445\,
            I => \N__56434\
        );

    \I__12481\ : Span12Mux_h
    port map (
            O => \N__56442\,
            I => \N__56434\
        );

    \I__12480\ : Span4Mux_h
    port map (
            O => \N__56439\,
            I => \N__56431\
        );

    \I__12479\ : Odrv12
    port map (
            O => \N__56434\,
            I => \ALU.N_967\
        );

    \I__12478\ : Odrv4
    port map (
            O => \N__56431\,
            I => \ALU.N_967\
        );

    \I__12477\ : CascadeMux
    port map (
            O => \N__56426\,
            I => \N__56423\
        );

    \I__12476\ : InMux
    port map (
            O => \N__56423\,
            I => \N__56420\
        );

    \I__12475\ : LocalMux
    port map (
            O => \N__56420\,
            I => \ALU.aluOut_i_3\
        );

    \I__12474\ : InMux
    port map (
            O => \N__56417\,
            I => \N__56410\
        );

    \I__12473\ : InMux
    port map (
            O => \N__56416\,
            I => \N__56407\
        );

    \I__12472\ : InMux
    port map (
            O => \N__56415\,
            I => \N__56402\
        );

    \I__12471\ : InMux
    port map (
            O => \N__56414\,
            I => \N__56402\
        );

    \I__12470\ : InMux
    port map (
            O => \N__56413\,
            I => \N__56398\
        );

    \I__12469\ : LocalMux
    port map (
            O => \N__56410\,
            I => \N__56395\
        );

    \I__12468\ : LocalMux
    port map (
            O => \N__56407\,
            I => \N__56391\
        );

    \I__12467\ : LocalMux
    port map (
            O => \N__56402\,
            I => \N__56388\
        );

    \I__12466\ : InMux
    port map (
            O => \N__56401\,
            I => \N__56385\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__56398\,
            I => \N__56382\
        );

    \I__12464\ : Span4Mux_v
    port map (
            O => \N__56395\,
            I => \N__56379\
        );

    \I__12463\ : InMux
    port map (
            O => \N__56394\,
            I => \N__56374\
        );

    \I__12462\ : Span4Mux_h
    port map (
            O => \N__56391\,
            I => \N__56371\
        );

    \I__12461\ : Span4Mux_h
    port map (
            O => \N__56388\,
            I => \N__56366\
        );

    \I__12460\ : LocalMux
    port map (
            O => \N__56385\,
            I => \N__56366\
        );

    \I__12459\ : Span4Mux_v
    port map (
            O => \N__56382\,
            I => \N__56361\
        );

    \I__12458\ : Span4Mux_h
    port map (
            O => \N__56379\,
            I => \N__56361\
        );

    \I__12457\ : InMux
    port map (
            O => \N__56378\,
            I => \N__56352\
        );

    \I__12456\ : InMux
    port map (
            O => \N__56377\,
            I => \N__56352\
        );

    \I__12455\ : LocalMux
    port map (
            O => \N__56374\,
            I => \N__56347\
        );

    \I__12454\ : Span4Mux_h
    port map (
            O => \N__56371\,
            I => \N__56347\
        );

    \I__12453\ : Span4Mux_h
    port map (
            O => \N__56366\,
            I => \N__56342\
        );

    \I__12452\ : Span4Mux_h
    port map (
            O => \N__56361\,
            I => \N__56339\
        );

    \I__12451\ : InMux
    port map (
            O => \N__56360\,
            I => \N__56336\
        );

    \I__12450\ : InMux
    port map (
            O => \N__56359\,
            I => \N__56329\
        );

    \I__12449\ : InMux
    port map (
            O => \N__56358\,
            I => \N__56329\
        );

    \I__12448\ : InMux
    port map (
            O => \N__56357\,
            I => \N__56329\
        );

    \I__12447\ : LocalMux
    port map (
            O => \N__56352\,
            I => \N__56321\
        );

    \I__12446\ : Span4Mux_h
    port map (
            O => \N__56347\,
            I => \N__56321\
        );

    \I__12445\ : InMux
    port map (
            O => \N__56346\,
            I => \N__56316\
        );

    \I__12444\ : InMux
    port map (
            O => \N__56345\,
            I => \N__56316\
        );

    \I__12443\ : Span4Mux_v
    port map (
            O => \N__56342\,
            I => \N__56313\
        );

    \I__12442\ : Span4Mux_h
    port map (
            O => \N__56339\,
            I => \N__56306\
        );

    \I__12441\ : LocalMux
    port map (
            O => \N__56336\,
            I => \N__56306\
        );

    \I__12440\ : LocalMux
    port map (
            O => \N__56329\,
            I => \N__56306\
        );

    \I__12439\ : InMux
    port map (
            O => \N__56328\,
            I => \N__56303\
        );

    \I__12438\ : InMux
    port map (
            O => \N__56327\,
            I => \N__56298\
        );

    \I__12437\ : InMux
    port map (
            O => \N__56326\,
            I => \N__56298\
        );

    \I__12436\ : Odrv4
    port map (
            O => \N__56321\,
            I => \ALU.status_19_3\
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__56316\,
            I => \ALU.status_19_3\
        );

    \I__12434\ : Odrv4
    port map (
            O => \N__56313\,
            I => \ALU.status_19_3\
        );

    \I__12433\ : Odrv4
    port map (
            O => \N__56306\,
            I => \ALU.status_19_3\
        );

    \I__12432\ : LocalMux
    port map (
            O => \N__56303\,
            I => \ALU.status_19_3\
        );

    \I__12431\ : LocalMux
    port map (
            O => \N__56298\,
            I => \ALU.status_19_3\
        );

    \I__12430\ : CascadeMux
    port map (
            O => \N__56285\,
            I => \N__56282\
        );

    \I__12429\ : InMux
    port map (
            O => \N__56282\,
            I => \N__56279\
        );

    \I__12428\ : LocalMux
    port map (
            O => \N__56279\,
            I => \ALU.aluOut_i_4\
        );

    \I__12427\ : InMux
    port map (
            O => \N__56276\,
            I => \N__56273\
        );

    \I__12426\ : LocalMux
    port map (
            O => \N__56273\,
            I => \N__56269\
        );

    \I__12425\ : CascadeMux
    port map (
            O => \N__56272\,
            I => \N__56263\
        );

    \I__12424\ : Span4Mux_h
    port map (
            O => \N__56269\,
            I => \N__56260\
        );

    \I__12423\ : CascadeMux
    port map (
            O => \N__56268\,
            I => \N__56256\
        );

    \I__12422\ : InMux
    port map (
            O => \N__56267\,
            I => \N__56253\
        );

    \I__12421\ : InMux
    port map (
            O => \N__56266\,
            I => \N__56250\
        );

    \I__12420\ : InMux
    port map (
            O => \N__56263\,
            I => \N__56247\
        );

    \I__12419\ : Span4Mux_v
    port map (
            O => \N__56260\,
            I => \N__56244\
        );

    \I__12418\ : InMux
    port map (
            O => \N__56259\,
            I => \N__56241\
        );

    \I__12417\ : InMux
    port map (
            O => \N__56256\,
            I => \N__56236\
        );

    \I__12416\ : LocalMux
    port map (
            O => \N__56253\,
            I => \N__56233\
        );

    \I__12415\ : LocalMux
    port map (
            O => \N__56250\,
            I => \N__56230\
        );

    \I__12414\ : LocalMux
    port map (
            O => \N__56247\,
            I => \N__56225\
        );

    \I__12413\ : Sp12to4
    port map (
            O => \N__56244\,
            I => \N__56218\
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__56241\,
            I => \N__56218\
        );

    \I__12411\ : InMux
    port map (
            O => \N__56240\,
            I => \N__56213\
        );

    \I__12410\ : InMux
    port map (
            O => \N__56239\,
            I => \N__56213\
        );

    \I__12409\ : LocalMux
    port map (
            O => \N__56236\,
            I => \N__56206\
        );

    \I__12408\ : Span4Mux_v
    port map (
            O => \N__56233\,
            I => \N__56206\
        );

    \I__12407\ : Span4Mux_h
    port map (
            O => \N__56230\,
            I => \N__56206\
        );

    \I__12406\ : CascadeMux
    port map (
            O => \N__56229\,
            I => \N__56203\
        );

    \I__12405\ : CascadeMux
    port map (
            O => \N__56228\,
            I => \N__56197\
        );

    \I__12404\ : Span4Mux_v
    port map (
            O => \N__56225\,
            I => \N__56193\
        );

    \I__12403\ : InMux
    port map (
            O => \N__56224\,
            I => \N__56188\
        );

    \I__12402\ : InMux
    port map (
            O => \N__56223\,
            I => \N__56188\
        );

    \I__12401\ : Span12Mux_h
    port map (
            O => \N__56218\,
            I => \N__56185\
        );

    \I__12400\ : LocalMux
    port map (
            O => \N__56213\,
            I => \N__56182\
        );

    \I__12399\ : Span4Mux_h
    port map (
            O => \N__56206\,
            I => \N__56179\
        );

    \I__12398\ : InMux
    port map (
            O => \N__56203\,
            I => \N__56168\
        );

    \I__12397\ : InMux
    port map (
            O => \N__56202\,
            I => \N__56168\
        );

    \I__12396\ : InMux
    port map (
            O => \N__56201\,
            I => \N__56168\
        );

    \I__12395\ : InMux
    port map (
            O => \N__56200\,
            I => \N__56168\
        );

    \I__12394\ : InMux
    port map (
            O => \N__56197\,
            I => \N__56168\
        );

    \I__12393\ : InMux
    port map (
            O => \N__56196\,
            I => \N__56165\
        );

    \I__12392\ : Odrv4
    port map (
            O => \N__56193\,
            I => \ALU.status_19_4\
        );

    \I__12391\ : LocalMux
    port map (
            O => \N__56188\,
            I => \ALU.status_19_4\
        );

    \I__12390\ : Odrv12
    port map (
            O => \N__56185\,
            I => \ALU.status_19_4\
        );

    \I__12389\ : Odrv4
    port map (
            O => \N__56182\,
            I => \ALU.status_19_4\
        );

    \I__12388\ : Odrv4
    port map (
            O => \N__56179\,
            I => \ALU.status_19_4\
        );

    \I__12387\ : LocalMux
    port map (
            O => \N__56168\,
            I => \ALU.status_19_4\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__56165\,
            I => \ALU.status_19_4\
        );

    \I__12385\ : CascadeMux
    port map (
            O => \N__56150\,
            I => \N__56147\
        );

    \I__12384\ : InMux
    port map (
            O => \N__56147\,
            I => \N__56144\
        );

    \I__12383\ : LocalMux
    port map (
            O => \N__56144\,
            I => \ALU.aluOut_i_5\
        );

    \I__12382\ : CascadeMux
    port map (
            O => \N__56141\,
            I => \N__56138\
        );

    \I__12381\ : InMux
    port map (
            O => \N__56138\,
            I => \N__56135\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__56135\,
            I => \N__56132\
        );

    \I__12379\ : Span4Mux_v
    port map (
            O => \N__56132\,
            I => \N__56127\
        );

    \I__12378\ : InMux
    port map (
            O => \N__56131\,
            I => \N__56124\
        );

    \I__12377\ : CascadeMux
    port map (
            O => \N__56130\,
            I => \N__56121\
        );

    \I__12376\ : Span4Mux_v
    port map (
            O => \N__56127\,
            I => \N__56117\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__56124\,
            I => \N__56112\
        );

    \I__12374\ : InMux
    port map (
            O => \N__56121\,
            I => \N__56109\
        );

    \I__12373\ : InMux
    port map (
            O => \N__56120\,
            I => \N__56106\
        );

    \I__12372\ : Span4Mux_h
    port map (
            O => \N__56117\,
            I => \N__56103\
        );

    \I__12371\ : InMux
    port map (
            O => \N__56116\,
            I => \N__56100\
        );

    \I__12370\ : InMux
    port map (
            O => \N__56115\,
            I => \N__56097\
        );

    \I__12369\ : Span4Mux_v
    port map (
            O => \N__56112\,
            I => \N__56093\
        );

    \I__12368\ : LocalMux
    port map (
            O => \N__56109\,
            I => \N__56090\
        );

    \I__12367\ : LocalMux
    port map (
            O => \N__56106\,
            I => \N__56087\
        );

    \I__12366\ : Span4Mux_h
    port map (
            O => \N__56103\,
            I => \N__56083\
        );

    \I__12365\ : LocalMux
    port map (
            O => \N__56100\,
            I => \N__56079\
        );

    \I__12364\ : LocalMux
    port map (
            O => \N__56097\,
            I => \N__56073\
        );

    \I__12363\ : CascadeMux
    port map (
            O => \N__56096\,
            I => \N__56070\
        );

    \I__12362\ : Span4Mux_v
    port map (
            O => \N__56093\,
            I => \N__56065\
        );

    \I__12361\ : Span4Mux_v
    port map (
            O => \N__56090\,
            I => \N__56060\
        );

    \I__12360\ : Span4Mux_v
    port map (
            O => \N__56087\,
            I => \N__56060\
        );

    \I__12359\ : InMux
    port map (
            O => \N__56086\,
            I => \N__56057\
        );

    \I__12358\ : Span4Mux_v
    port map (
            O => \N__56083\,
            I => \N__56054\
        );

    \I__12357\ : InMux
    port map (
            O => \N__56082\,
            I => \N__56051\
        );

    \I__12356\ : Span4Mux_v
    port map (
            O => \N__56079\,
            I => \N__56048\
        );

    \I__12355\ : InMux
    port map (
            O => \N__56078\,
            I => \N__56043\
        );

    \I__12354\ : InMux
    port map (
            O => \N__56077\,
            I => \N__56043\
        );

    \I__12353\ : InMux
    port map (
            O => \N__56076\,
            I => \N__56040\
        );

    \I__12352\ : Span4Mux_h
    port map (
            O => \N__56073\,
            I => \N__56037\
        );

    \I__12351\ : InMux
    port map (
            O => \N__56070\,
            I => \N__56032\
        );

    \I__12350\ : InMux
    port map (
            O => \N__56069\,
            I => \N__56032\
        );

    \I__12349\ : InMux
    port map (
            O => \N__56068\,
            I => \N__56029\
        );

    \I__12348\ : Sp12to4
    port map (
            O => \N__56065\,
            I => \N__56022\
        );

    \I__12347\ : Sp12to4
    port map (
            O => \N__56060\,
            I => \N__56022\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__56057\,
            I => \N__56022\
        );

    \I__12345\ : Odrv4
    port map (
            O => \N__56054\,
            I => \ALU.status_19_5\
        );

    \I__12344\ : LocalMux
    port map (
            O => \N__56051\,
            I => \ALU.status_19_5\
        );

    \I__12343\ : Odrv4
    port map (
            O => \N__56048\,
            I => \ALU.status_19_5\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__56043\,
            I => \ALU.status_19_5\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__56040\,
            I => \ALU.status_19_5\
        );

    \I__12340\ : Odrv4
    port map (
            O => \N__56037\,
            I => \ALU.status_19_5\
        );

    \I__12339\ : LocalMux
    port map (
            O => \N__56032\,
            I => \ALU.status_19_5\
        );

    \I__12338\ : LocalMux
    port map (
            O => \N__56029\,
            I => \ALU.status_19_5\
        );

    \I__12337\ : Odrv12
    port map (
            O => \N__56022\,
            I => \ALU.status_19_5\
        );

    \I__12336\ : CascadeMux
    port map (
            O => \N__56003\,
            I => \N__56000\
        );

    \I__12335\ : InMux
    port map (
            O => \N__56000\,
            I => \N__55997\
        );

    \I__12334\ : LocalMux
    port map (
            O => \N__55997\,
            I => \ALU.aluOut_i_6\
        );

    \I__12333\ : InMux
    port map (
            O => \N__55994\,
            I => \N__55986\
        );

    \I__12332\ : InMux
    port map (
            O => \N__55993\,
            I => \N__55979\
        );

    \I__12331\ : InMux
    port map (
            O => \N__55992\,
            I => \N__55979\
        );

    \I__12330\ : InMux
    port map (
            O => \N__55991\,
            I => \N__55976\
        );

    \I__12329\ : CascadeMux
    port map (
            O => \N__55990\,
            I => \N__55973\
        );

    \I__12328\ : InMux
    port map (
            O => \N__55989\,
            I => \N__55970\
        );

    \I__12327\ : LocalMux
    port map (
            O => \N__55986\,
            I => \N__55967\
        );

    \I__12326\ : InMux
    port map (
            O => \N__55985\,
            I => \N__55964\
        );

    \I__12325\ : CascadeMux
    port map (
            O => \N__55984\,
            I => \N__55961\
        );

    \I__12324\ : LocalMux
    port map (
            O => \N__55979\,
            I => \N__55954\
        );

    \I__12323\ : LocalMux
    port map (
            O => \N__55976\,
            I => \N__55950\
        );

    \I__12322\ : InMux
    port map (
            O => \N__55973\,
            I => \N__55946\
        );

    \I__12321\ : LocalMux
    port map (
            O => \N__55970\,
            I => \N__55941\
        );

    \I__12320\ : Span4Mux_v
    port map (
            O => \N__55967\,
            I => \N__55941\
        );

    \I__12319\ : LocalMux
    port map (
            O => \N__55964\,
            I => \N__55938\
        );

    \I__12318\ : InMux
    port map (
            O => \N__55961\,
            I => \N__55931\
        );

    \I__12317\ : InMux
    port map (
            O => \N__55960\,
            I => \N__55931\
        );

    \I__12316\ : InMux
    port map (
            O => \N__55959\,
            I => \N__55931\
        );

    \I__12315\ : InMux
    port map (
            O => \N__55958\,
            I => \N__55928\
        );

    \I__12314\ : InMux
    port map (
            O => \N__55957\,
            I => \N__55925\
        );

    \I__12313\ : Span4Mux_h
    port map (
            O => \N__55954\,
            I => \N__55922\
        );

    \I__12312\ : InMux
    port map (
            O => \N__55953\,
            I => \N__55919\
        );

    \I__12311\ : Span4Mux_v
    port map (
            O => \N__55950\,
            I => \N__55916\
        );

    \I__12310\ : InMux
    port map (
            O => \N__55949\,
            I => \N__55913\
        );

    \I__12309\ : LocalMux
    port map (
            O => \N__55946\,
            I => \N__55904\
        );

    \I__12308\ : Span4Mux_h
    port map (
            O => \N__55941\,
            I => \N__55904\
        );

    \I__12307\ : Span4Mux_v
    port map (
            O => \N__55938\,
            I => \N__55904\
        );

    \I__12306\ : LocalMux
    port map (
            O => \N__55931\,
            I => \N__55904\
        );

    \I__12305\ : LocalMux
    port map (
            O => \N__55928\,
            I => \N__55901\
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__55925\,
            I => \N__55898\
        );

    \I__12303\ : Span4Mux_h
    port map (
            O => \N__55922\,
            I => \N__55893\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__55919\,
            I => \N__55893\
        );

    \I__12301\ : Span4Mux_h
    port map (
            O => \N__55916\,
            I => \N__55888\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__55913\,
            I => \N__55888\
        );

    \I__12299\ : Span4Mux_h
    port map (
            O => \N__55904\,
            I => \N__55882\
        );

    \I__12298\ : Span4Mux_v
    port map (
            O => \N__55901\,
            I => \N__55879\
        );

    \I__12297\ : Span4Mux_v
    port map (
            O => \N__55898\,
            I => \N__55876\
        );

    \I__12296\ : Span4Mux_h
    port map (
            O => \N__55893\,
            I => \N__55872\
        );

    \I__12295\ : Span4Mux_v
    port map (
            O => \N__55888\,
            I => \N__55869\
        );

    \I__12294\ : InMux
    port map (
            O => \N__55887\,
            I => \N__55862\
        );

    \I__12293\ : InMux
    port map (
            O => \N__55886\,
            I => \N__55862\
        );

    \I__12292\ : InMux
    port map (
            O => \N__55885\,
            I => \N__55862\
        );

    \I__12291\ : Span4Mux_h
    port map (
            O => \N__55882\,
            I => \N__55859\
        );

    \I__12290\ : Span4Mux_v
    port map (
            O => \N__55879\,
            I => \N__55854\
        );

    \I__12289\ : Span4Mux_h
    port map (
            O => \N__55876\,
            I => \N__55854\
        );

    \I__12288\ : InMux
    port map (
            O => \N__55875\,
            I => \N__55851\
        );

    \I__12287\ : Span4Mux_v
    port map (
            O => \N__55872\,
            I => \N__55848\
        );

    \I__12286\ : Odrv4
    port map (
            O => \N__55869\,
            I => \ALU.status_19_6\
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__55862\,
            I => \ALU.status_19_6\
        );

    \I__12284\ : Odrv4
    port map (
            O => \N__55859\,
            I => \ALU.status_19_6\
        );

    \I__12283\ : Odrv4
    port map (
            O => \N__55854\,
            I => \ALU.status_19_6\
        );

    \I__12282\ : LocalMux
    port map (
            O => \N__55851\,
            I => \ALU.status_19_6\
        );

    \I__12281\ : Odrv4
    port map (
            O => \N__55848\,
            I => \ALU.status_19_6\
        );

    \I__12280\ : CascadeMux
    port map (
            O => \N__55835\,
            I => \N__55832\
        );

    \I__12279\ : InMux
    port map (
            O => \N__55832\,
            I => \N__55829\
        );

    \I__12278\ : LocalMux
    port map (
            O => \N__55829\,
            I => \N__55826\
        );

    \I__12277\ : Odrv4
    port map (
            O => \N__55826\,
            I => \ALU.aluOut_i_7\
        );

    \I__12276\ : CascadeMux
    port map (
            O => \N__55823\,
            I => \N__55818\
        );

    \I__12275\ : InMux
    port map (
            O => \N__55822\,
            I => \N__55813\
        );

    \I__12274\ : InMux
    port map (
            O => \N__55821\,
            I => \N__55808\
        );

    \I__12273\ : InMux
    port map (
            O => \N__55818\,
            I => \N__55805\
        );

    \I__12272\ : InMux
    port map (
            O => \N__55817\,
            I => \N__55802\
        );

    \I__12271\ : CascadeMux
    port map (
            O => \N__55816\,
            I => \N__55796\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__55813\,
            I => \N__55793\
        );

    \I__12269\ : InMux
    port map (
            O => \N__55812\,
            I => \N__55788\
        );

    \I__12268\ : InMux
    port map (
            O => \N__55811\,
            I => \N__55788\
        );

    \I__12267\ : LocalMux
    port map (
            O => \N__55808\,
            I => \N__55783\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__55805\,
            I => \N__55783\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__55802\,
            I => \N__55780\
        );

    \I__12264\ : InMux
    port map (
            O => \N__55801\,
            I => \N__55777\
        );

    \I__12263\ : InMux
    port map (
            O => \N__55800\,
            I => \N__55772\
        );

    \I__12262\ : InMux
    port map (
            O => \N__55799\,
            I => \N__55772\
        );

    \I__12261\ : InMux
    port map (
            O => \N__55796\,
            I => \N__55769\
        );

    \I__12260\ : Span4Mux_v
    port map (
            O => \N__55793\,
            I => \N__55764\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__55788\,
            I => \N__55761\
        );

    \I__12258\ : Span4Mux_v
    port map (
            O => \N__55783\,
            I => \N__55752\
        );

    \I__12257\ : Span4Mux_v
    port map (
            O => \N__55780\,
            I => \N__55752\
        );

    \I__12256\ : LocalMux
    port map (
            O => \N__55777\,
            I => \N__55752\
        );

    \I__12255\ : LocalMux
    port map (
            O => \N__55772\,
            I => \N__55752\
        );

    \I__12254\ : LocalMux
    port map (
            O => \N__55769\,
            I => \N__55749\
        );

    \I__12253\ : InMux
    port map (
            O => \N__55768\,
            I => \N__55746\
        );

    \I__12252\ : InMux
    port map (
            O => \N__55767\,
            I => \N__55743\
        );

    \I__12251\ : Sp12to4
    port map (
            O => \N__55764\,
            I => \N__55740\
        );

    \I__12250\ : Span4Mux_h
    port map (
            O => \N__55761\,
            I => \N__55737\
        );

    \I__12249\ : Span4Mux_h
    port map (
            O => \N__55752\,
            I => \N__55734\
        );

    \I__12248\ : Span4Mux_h
    port map (
            O => \N__55749\,
            I => \N__55727\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__55746\,
            I => \N__55727\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__55743\,
            I => \N__55727\
        );

    \I__12245\ : Span12Mux_h
    port map (
            O => \N__55740\,
            I => \N__55721\
        );

    \I__12244\ : Span4Mux_v
    port map (
            O => \N__55737\,
            I => \N__55716\
        );

    \I__12243\ : Span4Mux_v
    port map (
            O => \N__55734\,
            I => \N__55716\
        );

    \I__12242\ : Span4Mux_v
    port map (
            O => \N__55727\,
            I => \N__55713\
        );

    \I__12241\ : InMux
    port map (
            O => \N__55726\,
            I => \N__55706\
        );

    \I__12240\ : InMux
    port map (
            O => \N__55725\,
            I => \N__55706\
        );

    \I__12239\ : InMux
    port map (
            O => \N__55724\,
            I => \N__55706\
        );

    \I__12238\ : Odrv12
    port map (
            O => \N__55721\,
            I => \ALU.status_19_7\
        );

    \I__12237\ : Odrv4
    port map (
            O => \N__55716\,
            I => \ALU.status_19_7\
        );

    \I__12236\ : Odrv4
    port map (
            O => \N__55713\,
            I => \ALU.status_19_7\
        );

    \I__12235\ : LocalMux
    port map (
            O => \N__55706\,
            I => \ALU.status_19_7\
        );

    \I__12234\ : CascadeMux
    port map (
            O => \N__55697\,
            I => \N__55694\
        );

    \I__12233\ : InMux
    port map (
            O => \N__55694\,
            I => \N__55691\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__55691\,
            I => \ALU.aluOut_i_8\
        );

    \I__12231\ : CascadeMux
    port map (
            O => \N__55688\,
            I => \N__55682\
        );

    \I__12230\ : InMux
    port map (
            O => \N__55687\,
            I => \N__55678\
        );

    \I__12229\ : CascadeMux
    port map (
            O => \N__55686\,
            I => \N__55675\
        );

    \I__12228\ : CascadeMux
    port map (
            O => \N__55685\,
            I => \N__55671\
        );

    \I__12227\ : InMux
    port map (
            O => \N__55682\,
            I => \N__55665\
        );

    \I__12226\ : InMux
    port map (
            O => \N__55681\,
            I => \N__55665\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__55678\,
            I => \N__55662\
        );

    \I__12224\ : InMux
    port map (
            O => \N__55675\,
            I => \N__55657\
        );

    \I__12223\ : InMux
    port map (
            O => \N__55674\,
            I => \N__55654\
        );

    \I__12222\ : InMux
    port map (
            O => \N__55671\,
            I => \N__55651\
        );

    \I__12221\ : CascadeMux
    port map (
            O => \N__55670\,
            I => \N__55648\
        );

    \I__12220\ : LocalMux
    port map (
            O => \N__55665\,
            I => \N__55644\
        );

    \I__12219\ : Span12Mux_s8_v
    port map (
            O => \N__55662\,
            I => \N__55641\
        );

    \I__12218\ : InMux
    port map (
            O => \N__55661\,
            I => \N__55638\
        );

    \I__12217\ : InMux
    port map (
            O => \N__55660\,
            I => \N__55635\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__55657\,
            I => \N__55628\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__55654\,
            I => \N__55628\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__55651\,
            I => \N__55628\
        );

    \I__12213\ : InMux
    port map (
            O => \N__55648\,
            I => \N__55625\
        );

    \I__12212\ : InMux
    port map (
            O => \N__55647\,
            I => \N__55622\
        );

    \I__12211\ : Span4Mux_v
    port map (
            O => \N__55644\,
            I => \N__55619\
        );

    \I__12210\ : Span12Mux_h
    port map (
            O => \N__55641\,
            I => \N__55612\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__55638\,
            I => \N__55612\
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__55635\,
            I => \N__55612\
        );

    \I__12207\ : Span4Mux_h
    port map (
            O => \N__55628\,
            I => \N__55609\
        );

    \I__12206\ : LocalMux
    port map (
            O => \N__55625\,
            I => \ALU.status_19_8\
        );

    \I__12205\ : LocalMux
    port map (
            O => \N__55622\,
            I => \ALU.status_19_8\
        );

    \I__12204\ : Odrv4
    port map (
            O => \N__55619\,
            I => \ALU.status_19_8\
        );

    \I__12203\ : Odrv12
    port map (
            O => \N__55612\,
            I => \ALU.status_19_8\
        );

    \I__12202\ : Odrv4
    port map (
            O => \N__55609\,
            I => \ALU.status_19_8\
        );

    \I__12201\ : CascadeMux
    port map (
            O => \N__55598\,
            I => \N__55595\
        );

    \I__12200\ : InMux
    port map (
            O => \N__55595\,
            I => \N__55592\
        );

    \I__12199\ : LocalMux
    port map (
            O => \N__55592\,
            I => \ALU.aluOut_i_9\
        );

    \I__12198\ : InMux
    port map (
            O => \N__55589\,
            I => \N__55586\
        );

    \I__12197\ : LocalMux
    port map (
            O => \N__55586\,
            I => \N__55582\
        );

    \I__12196\ : InMux
    port map (
            O => \N__55585\,
            I => \N__55579\
        );

    \I__12195\ : Span4Mux_v
    port map (
            O => \N__55582\,
            I => \N__55573\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__55579\,
            I => \N__55570\
        );

    \I__12193\ : InMux
    port map (
            O => \N__55578\,
            I => \N__55565\
        );

    \I__12192\ : InMux
    port map (
            O => \N__55577\,
            I => \N__55565\
        );

    \I__12191\ : InMux
    port map (
            O => \N__55576\,
            I => \N__55562\
        );

    \I__12190\ : Sp12to4
    port map (
            O => \N__55573\,
            I => \N__55559\
        );

    \I__12189\ : Span4Mux_h
    port map (
            O => \N__55570\,
            I => \N__55555\
        );

    \I__12188\ : LocalMux
    port map (
            O => \N__55565\,
            I => \N__55550\
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__55562\,
            I => \N__55550\
        );

    \I__12186\ : Span12Mux_h
    port map (
            O => \N__55559\,
            I => \N__55543\
        );

    \I__12185\ : InMux
    port map (
            O => \N__55558\,
            I => \N__55540\
        );

    \I__12184\ : Span4Mux_v
    port map (
            O => \N__55555\,
            I => \N__55535\
        );

    \I__12183\ : Span4Mux_h
    port map (
            O => \N__55550\,
            I => \N__55535\
        );

    \I__12182\ : InMux
    port map (
            O => \N__55549\,
            I => \N__55526\
        );

    \I__12181\ : InMux
    port map (
            O => \N__55548\,
            I => \N__55526\
        );

    \I__12180\ : InMux
    port map (
            O => \N__55547\,
            I => \N__55526\
        );

    \I__12179\ : InMux
    port map (
            O => \N__55546\,
            I => \N__55526\
        );

    \I__12178\ : Odrv12
    port map (
            O => \N__55543\,
            I => \ALU.status_19_9\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__55540\,
            I => \ALU.status_19_9\
        );

    \I__12176\ : Odrv4
    port map (
            O => \N__55535\,
            I => \ALU.status_19_9\
        );

    \I__12175\ : LocalMux
    port map (
            O => \N__55526\,
            I => \ALU.status_19_9\
        );

    \I__12174\ : CascadeMux
    port map (
            O => \N__55517\,
            I => \N__55514\
        );

    \I__12173\ : InMux
    port map (
            O => \N__55514\,
            I => \N__55511\
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__55511\,
            I => \N__55508\
        );

    \I__12171\ : Odrv4
    port map (
            O => \N__55508\,
            I => \ALU.aluOut_i_10\
        );

    \I__12170\ : CascadeMux
    port map (
            O => \N__55505\,
            I => \N__55502\
        );

    \I__12169\ : InMux
    port map (
            O => \N__55502\,
            I => \N__55499\
        );

    \I__12168\ : LocalMux
    port map (
            O => \N__55499\,
            I => \N__55496\
        );

    \I__12167\ : Span4Mux_v
    port map (
            O => \N__55496\,
            I => \N__55493\
        );

    \I__12166\ : Sp12to4
    port map (
            O => \N__55493\,
            I => \N__55490\
        );

    \I__12165\ : Span12Mux_h
    port map (
            O => \N__55490\,
            I => \N__55487\
        );

    \I__12164\ : Odrv12
    port map (
            O => \N__55487\,
            I => \PROM.ROMDATA.m158\
        );

    \I__12163\ : CascadeMux
    port map (
            O => \N__55484\,
            I => \PROM.ROMDATA.m158_cascade_\
        );

    \I__12162\ : InMux
    port map (
            O => \N__55481\,
            I => \N__55478\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__55478\,
            I => \PROM.ROMDATA.m196_ns\
        );

    \I__12160\ : InMux
    port map (
            O => \N__55475\,
            I => \N__55467\
        );

    \I__12159\ : InMux
    port map (
            O => \N__55474\,
            I => \N__55462\
        );

    \I__12158\ : InMux
    port map (
            O => \N__55473\,
            I => \N__55457\
        );

    \I__12157\ : InMux
    port map (
            O => \N__55472\,
            I => \N__55457\
        );

    \I__12156\ : InMux
    port map (
            O => \N__55471\,
            I => \N__55448\
        );

    \I__12155\ : InMux
    port map (
            O => \N__55470\,
            I => \N__55445\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__55467\,
            I => \N__55441\
        );

    \I__12153\ : InMux
    port map (
            O => \N__55466\,
            I => \N__55436\
        );

    \I__12152\ : InMux
    port map (
            O => \N__55465\,
            I => \N__55436\
        );

    \I__12151\ : LocalMux
    port map (
            O => \N__55462\,
            I => \N__55431\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__55457\,
            I => \N__55431\
        );

    \I__12149\ : InMux
    port map (
            O => \N__55456\,
            I => \N__55424\
        );

    \I__12148\ : InMux
    port map (
            O => \N__55455\,
            I => \N__55424\
        );

    \I__12147\ : InMux
    port map (
            O => \N__55454\,
            I => \N__55424\
        );

    \I__12146\ : InMux
    port map (
            O => \N__55453\,
            I => \N__55418\
        );

    \I__12145\ : InMux
    port map (
            O => \N__55452\,
            I => \N__55413\
        );

    \I__12144\ : InMux
    port map (
            O => \N__55451\,
            I => \N__55413\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__55448\,
            I => \N__55408\
        );

    \I__12142\ : LocalMux
    port map (
            O => \N__55445\,
            I => \N__55408\
        );

    \I__12141\ : InMux
    port map (
            O => \N__55444\,
            I => \N__55405\
        );

    \I__12140\ : Span4Mux_v
    port map (
            O => \N__55441\,
            I => \N__55400\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__55436\,
            I => \N__55400\
        );

    \I__12138\ : Span4Mux_h
    port map (
            O => \N__55431\,
            I => \N__55396\
        );

    \I__12137\ : LocalMux
    port map (
            O => \N__55424\,
            I => \N__55393\
        );

    \I__12136\ : InMux
    port map (
            O => \N__55423\,
            I => \N__55386\
        );

    \I__12135\ : InMux
    port map (
            O => \N__55422\,
            I => \N__55386\
        );

    \I__12134\ : InMux
    port map (
            O => \N__55421\,
            I => \N__55386\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__55418\,
            I => \N__55381\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__55413\,
            I => \N__55381\
        );

    \I__12131\ : Span4Mux_h
    port map (
            O => \N__55408\,
            I => \N__55376\
        );

    \I__12130\ : LocalMux
    port map (
            O => \N__55405\,
            I => \N__55376\
        );

    \I__12129\ : Span4Mux_h
    port map (
            O => \N__55400\,
            I => \N__55373\
        );

    \I__12128\ : InMux
    port map (
            O => \N__55399\,
            I => \N__55370\
        );

    \I__12127\ : Span4Mux_h
    port map (
            O => \N__55396\,
            I => \N__55365\
        );

    \I__12126\ : Span4Mux_h
    port map (
            O => \N__55393\,
            I => \N__55365\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__55386\,
            I => \N__55360\
        );

    \I__12124\ : Span4Mux_v
    port map (
            O => \N__55381\,
            I => \N__55360\
        );

    \I__12123\ : Span4Mux_h
    port map (
            O => \N__55376\,
            I => \N__55357\
        );

    \I__12122\ : Span4Mux_h
    port map (
            O => \N__55373\,
            I => \N__55354\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__55370\,
            I => \N__55351\
        );

    \I__12120\ : Span4Mux_v
    port map (
            O => \N__55365\,
            I => \N__55346\
        );

    \I__12119\ : Span4Mux_h
    port map (
            O => \N__55360\,
            I => \N__55346\
        );

    \I__12118\ : Span4Mux_h
    port map (
            O => \N__55357\,
            I => \N__55343\
        );

    \I__12117\ : Odrv4
    port map (
            O => \N__55354\,
            I => \PROM_ROMDATA_dintern_6ro\
        );

    \I__12116\ : Odrv12
    port map (
            O => \N__55351\,
            I => \PROM_ROMDATA_dintern_6ro\
        );

    \I__12115\ : Odrv4
    port map (
            O => \N__55346\,
            I => \PROM_ROMDATA_dintern_6ro\
        );

    \I__12114\ : Odrv4
    port map (
            O => \N__55343\,
            I => \PROM_ROMDATA_dintern_6ro\
        );

    \I__12113\ : InMux
    port map (
            O => \N__55334\,
            I => \N__55330\
        );

    \I__12112\ : InMux
    port map (
            O => \N__55333\,
            I => \N__55327\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__55330\,
            I => \N__55324\
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__55327\,
            I => \N__55321\
        );

    \I__12109\ : Span4Mux_v
    port map (
            O => \N__55324\,
            I => \N__55318\
        );

    \I__12108\ : Span12Mux_v
    port map (
            O => \N__55321\,
            I => \N__55315\
        );

    \I__12107\ : Span4Mux_h
    port map (
            O => \N__55318\,
            I => \N__55312\
        );

    \I__12106\ : Span12Mux_h
    port map (
            O => \N__55315\,
            I => \N__55309\
        );

    \I__12105\ : Span4Mux_h
    port map (
            O => \N__55312\,
            I => \N__55306\
        );

    \I__12104\ : Odrv12
    port map (
            O => \N__55309\,
            I => \CONTROL.ctrlOut_4\
        );

    \I__12103\ : Odrv4
    port map (
            O => \N__55306\,
            I => \CONTROL.ctrlOut_4\
        );

    \I__12102\ : InMux
    port map (
            O => \N__55301\,
            I => \N__55298\
        );

    \I__12101\ : LocalMux
    port map (
            O => \N__55298\,
            I => \N__55295\
        );

    \I__12100\ : Span4Mux_h
    port map (
            O => \N__55295\,
            I => \N__55291\
        );

    \I__12099\ : InMux
    port map (
            O => \N__55294\,
            I => \N__55288\
        );

    \I__12098\ : Odrv4
    port map (
            O => \N__55291\,
            I => \CONTROL.dout_reto_4\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__55288\,
            I => \CONTROL.dout_reto_4\
        );

    \I__12096\ : CascadeMux
    port map (
            O => \N__55283\,
            I => \N__55280\
        );

    \I__12095\ : InMux
    port map (
            O => \N__55280\,
            I => \N__55277\
        );

    \I__12094\ : LocalMux
    port map (
            O => \N__55277\,
            I => \ALU.aluOut_i_0\
        );

    \I__12093\ : CascadeMux
    port map (
            O => \N__55274\,
            I => \N__55271\
        );

    \I__12092\ : InMux
    port map (
            O => \N__55271\,
            I => \N__55268\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__55268\,
            I => \ALU.aluOut_i_1\
        );

    \I__12090\ : CascadeMux
    port map (
            O => \N__55265\,
            I => \N__55262\
        );

    \I__12089\ : InMux
    port map (
            O => \N__55262\,
            I => \N__55259\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__55259\,
            I => \ALU.aluOut_i_2\
        );

    \I__12087\ : CascadeMux
    port map (
            O => \N__55256\,
            I => \PROM.ROMDATA.m183_cascade_\
        );

    \I__12086\ : InMux
    port map (
            O => \N__55253\,
            I => \N__55250\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__55250\,
            I => \PROM.ROMDATA.m185_bm\
        );

    \I__12084\ : CascadeMux
    port map (
            O => \N__55247\,
            I => \PROM.ROMDATA.N_525_mux_cascade_\
        );

    \I__12083\ : InMux
    port map (
            O => \N__55244\,
            I => \N__55241\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__55241\,
            I => \PROM.ROMDATA.i4_mux\
        );

    \I__12081\ : InMux
    port map (
            O => \N__55238\,
            I => \N__55235\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__55235\,
            I => \N__55232\
        );

    \I__12079\ : Span4Mux_h
    port map (
            O => \N__55232\,
            I => \N__55229\
        );

    \I__12078\ : Odrv4
    port map (
            O => \N__55229\,
            I => \PROM.ROMDATA.m103\
        );

    \I__12077\ : InMux
    port map (
            O => \N__55226\,
            I => \N__55223\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__55223\,
            I => \N__55218\
        );

    \I__12075\ : InMux
    port map (
            O => \N__55222\,
            I => \N__55215\
        );

    \I__12074\ : InMux
    port map (
            O => \N__55221\,
            I => \N__55212\
        );

    \I__12073\ : Odrv12
    port map (
            O => \N__55218\,
            I => \PROM.ROMDATA.m226\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__55215\,
            I => \PROM.ROMDATA.m226\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__55212\,
            I => \PROM.ROMDATA.m226\
        );

    \I__12070\ : CascadeMux
    port map (
            O => \N__55205\,
            I => \N__55202\
        );

    \I__12069\ : InMux
    port map (
            O => \N__55202\,
            I => \N__55199\
        );

    \I__12068\ : LocalMux
    port map (
            O => \N__55199\,
            I => \PROM.ROMDATA.m92_am_1\
        );

    \I__12067\ : InMux
    port map (
            O => \N__55196\,
            I => \N__55193\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__55193\,
            I => \N__55190\
        );

    \I__12065\ : Span4Mux_h
    port map (
            O => \N__55190\,
            I => \N__55187\
        );

    \I__12064\ : Odrv4
    port map (
            O => \N__55187\,
            I => \PROM.ROMDATA.m55\
        );

    \I__12063\ : InMux
    port map (
            O => \N__55184\,
            I => \N__55180\
        );

    \I__12062\ : InMux
    port map (
            O => \N__55183\,
            I => \N__55177\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__55180\,
            I => \N__55174\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__55177\,
            I => \CONTROL.programCounter_1_reto_4\
        );

    \I__12059\ : Odrv4
    port map (
            O => \N__55174\,
            I => \CONTROL.programCounter_1_reto_4\
        );

    \I__12058\ : InMux
    port map (
            O => \N__55169\,
            I => \N__55164\
        );

    \I__12057\ : InMux
    port map (
            O => \N__55168\,
            I => \N__55159\
        );

    \I__12056\ : InMux
    port map (
            O => \N__55167\,
            I => \N__55159\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__55164\,
            I => \N__55156\
        );

    \I__12054\ : LocalMux
    port map (
            O => \N__55159\,
            I => \N__55152\
        );

    \I__12053\ : Span4Mux_h
    port map (
            O => \N__55156\,
            I => \N__55149\
        );

    \I__12052\ : InMux
    port map (
            O => \N__55155\,
            I => \N__55146\
        );

    \I__12051\ : Odrv12
    port map (
            O => \N__55152\,
            I => \CONTROL_addrstack_reto_4\
        );

    \I__12050\ : Odrv4
    port map (
            O => \N__55149\,
            I => \CONTROL_addrstack_reto_4\
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__55146\,
            I => \CONTROL_addrstack_reto_4\
        );

    \I__12048\ : InMux
    port map (
            O => \N__55139\,
            I => \N__55134\
        );

    \I__12047\ : InMux
    port map (
            O => \N__55138\,
            I => \N__55131\
        );

    \I__12046\ : InMux
    port map (
            O => \N__55137\,
            I => \N__55128\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__55134\,
            I => \N__55125\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__55131\,
            I => \N__55115\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__55128\,
            I => \N__55112\
        );

    \I__12042\ : Span4Mux_h
    port map (
            O => \N__55125\,
            I => \N__55109\
        );

    \I__12041\ : InMux
    port map (
            O => \N__55124\,
            I => \N__55104\
        );

    \I__12040\ : InMux
    port map (
            O => \N__55123\,
            I => \N__55104\
        );

    \I__12039\ : InMux
    port map (
            O => \N__55122\,
            I => \N__55099\
        );

    \I__12038\ : InMux
    port map (
            O => \N__55121\,
            I => \N__55099\
        );

    \I__12037\ : InMux
    port map (
            O => \N__55120\,
            I => \N__55092\
        );

    \I__12036\ : InMux
    port map (
            O => \N__55119\,
            I => \N__55092\
        );

    \I__12035\ : InMux
    port map (
            O => \N__55118\,
            I => \N__55092\
        );

    \I__12034\ : Odrv4
    port map (
            O => \N__55115\,
            I => \CONTROL.programCounter11_reto_fast\
        );

    \I__12033\ : Odrv4
    port map (
            O => \N__55112\,
            I => \CONTROL.programCounter11_reto_fast\
        );

    \I__12032\ : Odrv4
    port map (
            O => \N__55109\,
            I => \CONTROL.programCounter11_reto_fast\
        );

    \I__12031\ : LocalMux
    port map (
            O => \N__55104\,
            I => \CONTROL.programCounter11_reto_fast\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__55099\,
            I => \CONTROL.programCounter11_reto_fast\
        );

    \I__12029\ : LocalMux
    port map (
            O => \N__55092\,
            I => \CONTROL.programCounter11_reto_fast\
        );

    \I__12028\ : InMux
    port map (
            O => \N__55079\,
            I => \N__55074\
        );

    \I__12027\ : InMux
    port map (
            O => \N__55078\,
            I => \N__55071\
        );

    \I__12026\ : InMux
    port map (
            O => \N__55077\,
            I => \N__55068\
        );

    \I__12025\ : LocalMux
    port map (
            O => \N__55074\,
            I => \N__55065\
        );

    \I__12024\ : LocalMux
    port map (
            O => \N__55071\,
            I => \N__55059\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__55068\,
            I => \N__55059\
        );

    \I__12022\ : Span4Mux_v
    port map (
            O => \N__55065\,
            I => \N__55050\
        );

    \I__12021\ : InMux
    port map (
            O => \N__55064\,
            I => \N__55047\
        );

    \I__12020\ : Span4Mux_v
    port map (
            O => \N__55059\,
            I => \N__55044\
        );

    \I__12019\ : InMux
    port map (
            O => \N__55058\,
            I => \N__55041\
        );

    \I__12018\ : InMux
    port map (
            O => \N__55057\,
            I => \N__55036\
        );

    \I__12017\ : InMux
    port map (
            O => \N__55056\,
            I => \N__55036\
        );

    \I__12016\ : InMux
    port map (
            O => \N__55055\,
            I => \N__55033\
        );

    \I__12015\ : InMux
    port map (
            O => \N__55054\,
            I => \N__55028\
        );

    \I__12014\ : InMux
    port map (
            O => \N__55053\,
            I => \N__55028\
        );

    \I__12013\ : Odrv4
    port map (
            O => \N__55050\,
            I => \CONTROL.un1_programCounter9_reto_fast\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__55047\,
            I => \CONTROL.un1_programCounter9_reto_fast\
        );

    \I__12011\ : Odrv4
    port map (
            O => \N__55044\,
            I => \CONTROL.un1_programCounter9_reto_fast\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__55041\,
            I => \CONTROL.un1_programCounter9_reto_fast\
        );

    \I__12009\ : LocalMux
    port map (
            O => \N__55036\,
            I => \CONTROL.un1_programCounter9_reto_fast\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__55033\,
            I => \CONTROL.un1_programCounter9_reto_fast\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__55028\,
            I => \CONTROL.un1_programCounter9_reto_fast\
        );

    \I__12006\ : CascadeMux
    port map (
            O => \N__55013\,
            I => \CONTROL.programCounter_ret_1_RNINC8IZ0Z_4_cascade_\
        );

    \I__12005\ : InMux
    port map (
            O => \N__55010\,
            I => \N__55007\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__55007\,
            I => \N__55004\
        );

    \I__12003\ : Span4Mux_h
    port map (
            O => \N__55004\,
            I => \N__55001\
        );

    \I__12002\ : Odrv4
    port map (
            O => \N__55001\,
            I => \CONTROL.programCounter_ret_19_RNIGQ8JZ0Z_4\
        );

    \I__12001\ : InMux
    port map (
            O => \N__54998\,
            I => \N__54995\
        );

    \I__12000\ : LocalMux
    port map (
            O => \N__54995\,
            I => \PROM.ROMDATA.m143\
        );

    \I__11999\ : CascadeMux
    port map (
            O => \N__54992\,
            I => \progRomAddress_4_cascade_\
        );

    \I__11998\ : InMux
    port map (
            O => \N__54989\,
            I => \N__54986\
        );

    \I__11997\ : LocalMux
    port map (
            O => \N__54986\,
            I => \N__54983\
        );

    \I__11996\ : Odrv4
    port map (
            O => \N__54983\,
            I => \PROM.ROMDATA.m145\
        );

    \I__11995\ : InMux
    port map (
            O => \N__54980\,
            I => \N__54977\
        );

    \I__11994\ : LocalMux
    port map (
            O => \N__54977\,
            I => \N__54974\
        );

    \I__11993\ : Span12Mux_s11_h
    port map (
            O => \N__54974\,
            I => \N__54971\
        );

    \I__11992\ : Odrv12
    port map (
            O => \N__54971\,
            I => \PROM.ROMDATA.m90\
        );

    \I__11991\ : InMux
    port map (
            O => \N__54968\,
            I => \N__54965\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__54965\,
            I => \N__54962\
        );

    \I__11989\ : Span4Mux_h
    port map (
            O => \N__54962\,
            I => \N__54959\
        );

    \I__11988\ : Odrv4
    port map (
            O => \N__54959\,
            I => \PROM.ROMDATA.m92_bm\
        );

    \I__11987\ : InMux
    port map (
            O => \N__54956\,
            I => \N__54953\
        );

    \I__11986\ : LocalMux
    port map (
            O => \N__54953\,
            I => \N__54950\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__54950\,
            I => \N__54947\
        );

    \I__11984\ : Odrv4
    port map (
            O => \N__54947\,
            I => \PROM.ROMDATA.m11_am\
        );

    \I__11983\ : CascadeMux
    port map (
            O => \N__54944\,
            I => \PROM.ROMDATA.m19_ns_1_cascade_\
        );

    \I__11982\ : InMux
    port map (
            O => \N__54941\,
            I => \N__54938\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__54938\,
            I => \PROM.ROMDATA.m18_am\
        );

    \I__11980\ : InMux
    port map (
            O => \N__54935\,
            I => \N__54932\
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__54932\,
            I => \N__54929\
        );

    \I__11978\ : Span4Mux_v
    port map (
            O => \N__54929\,
            I => \N__54926\
        );

    \I__11977\ : Odrv4
    port map (
            O => \N__54926\,
            I => \PROM.ROMDATA.m19_ns\
        );

    \I__11976\ : CascadeMux
    port map (
            O => \N__54923\,
            I => \N__54919\
        );

    \I__11975\ : InMux
    port map (
            O => \N__54922\,
            I => \N__54916\
        );

    \I__11974\ : InMux
    port map (
            O => \N__54919\,
            I => \N__54913\
        );

    \I__11973\ : LocalMux
    port map (
            O => \N__54916\,
            I => \N__54908\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__54913\,
            I => \N__54908\
        );

    \I__11971\ : Span4Mux_v
    port map (
            O => \N__54908\,
            I => \N__54905\
        );

    \I__11970\ : Odrv4
    port map (
            O => \N__54905\,
            I => \PROM.ROMDATA.m33\
        );

    \I__11969\ : InMux
    port map (
            O => \N__54902\,
            I => \N__54898\
        );

    \I__11968\ : InMux
    port map (
            O => \N__54901\,
            I => \N__54895\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__54898\,
            I => \CONTROL.dout_reto_1\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__54895\,
            I => \CONTROL.dout_reto_1\
        );

    \I__11965\ : InMux
    port map (
            O => \N__54890\,
            I => \N__54884\
        );

    \I__11964\ : InMux
    port map (
            O => \N__54889\,
            I => \N__54884\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__54884\,
            I => \N__54881\
        );

    \I__11962\ : Span4Mux_v
    port map (
            O => \N__54881\,
            I => \N__54878\
        );

    \I__11961\ : Odrv4
    port map (
            O => \N__54878\,
            I => \CONTROL.programCounter_1_reto_1\
        );

    \I__11960\ : CascadeMux
    port map (
            O => \N__54875\,
            I => \CONTROL.programCounter_ret_1_RNIH68IZ0Z_1_cascade_\
        );

    \I__11959\ : InMux
    port map (
            O => \N__54872\,
            I => \N__54869\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__54869\,
            I => \CONTROL.programCounter_ret_19_RNIAK8JZ0Z_1\
        );

    \I__11957\ : CascadeMux
    port map (
            O => \N__54866\,
            I => \progRomAddress_1_cascade_\
        );

    \I__11956\ : InMux
    port map (
            O => \N__54863\,
            I => \N__54860\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__54860\,
            I => \PROM.ROMDATA.m437_ns\
        );

    \I__11954\ : InMux
    port map (
            O => \N__54857\,
            I => \N__54854\
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__54854\,
            I => \PROM.ROMDATA.m312_bm\
        );

    \I__11952\ : InMux
    port map (
            O => \N__54851\,
            I => \N__54848\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__54848\,
            I => \N__54845\
        );

    \I__11950\ : Span4Mux_h
    port map (
            O => \N__54845\,
            I => \N__54842\
        );

    \I__11949\ : Span4Mux_h
    port map (
            O => \N__54842\,
            I => \N__54839\
        );

    \I__11948\ : Odrv4
    port map (
            O => \N__54839\,
            I => \PROM.ROMDATA.m312_am\
        );

    \I__11947\ : InMux
    port map (
            O => \N__54836\,
            I => \N__54833\
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__54833\,
            I => \PROM.ROMDATA.m437_ns_1\
        );

    \I__11945\ : InMux
    port map (
            O => \N__54830\,
            I => \N__54827\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__54827\,
            I => \PROM.ROMDATA.m11_bm\
        );

    \I__11943\ : CascadeMux
    port map (
            O => \N__54824\,
            I => \PROM.ROMDATA.m18_bm_cascade_\
        );

    \I__11942\ : InMux
    port map (
            O => \N__54821\,
            I => \N__54818\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__54818\,
            I => \N__54815\
        );

    \I__11940\ : Span12Mux_v
    port map (
            O => \N__54815\,
            I => \N__54811\
        );

    \I__11939\ : InMux
    port map (
            O => \N__54814\,
            I => \N__54808\
        );

    \I__11938\ : Odrv12
    port map (
            O => \N__54811\,
            I => \CONTROL.ctrlOut_2\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__54808\,
            I => \CONTROL.ctrlOut_2\
        );

    \I__11936\ : InMux
    port map (
            O => \N__54803\,
            I => \N__54799\
        );

    \I__11935\ : InMux
    port map (
            O => \N__54802\,
            I => \N__54796\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__54799\,
            I => \N__54791\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__54796\,
            I => \N__54791\
        );

    \I__11932\ : Span4Mux_h
    port map (
            O => \N__54791\,
            I => \N__54788\
        );

    \I__11931\ : Span4Mux_v
    port map (
            O => \N__54788\,
            I => \N__54785\
        );

    \I__11930\ : Odrv4
    port map (
            O => \N__54785\,
            I => \CONTROL.dout_reto_2\
        );

    \I__11929\ : InMux
    port map (
            O => \N__54782\,
            I => \N__54779\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__54779\,
            I => \N__54776\
        );

    \I__11927\ : Span12Mux_v
    port map (
            O => \N__54776\,
            I => \N__54773\
        );

    \I__11926\ : Odrv12
    port map (
            O => \N__54773\,
            I => \CONTROL.N_136_0\
        );

    \I__11925\ : InMux
    port map (
            O => \N__54770\,
            I => \N__54767\
        );

    \I__11924\ : LocalMux
    port map (
            O => \N__54767\,
            I => \N__54763\
        );

    \I__11923\ : InMux
    port map (
            O => \N__54766\,
            I => \N__54760\
        );

    \I__11922\ : Span4Mux_v
    port map (
            O => \N__54763\,
            I => \N__54757\
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__54760\,
            I => \CONTROL.N_86_0\
        );

    \I__11920\ : Odrv4
    port map (
            O => \N__54757\,
            I => \CONTROL.N_86_0\
        );

    \I__11919\ : CascadeMux
    port map (
            O => \N__54752\,
            I => \N__54747\
        );

    \I__11918\ : InMux
    port map (
            O => \N__54751\,
            I => \N__54741\
        );

    \I__11917\ : InMux
    port map (
            O => \N__54750\,
            I => \N__54741\
        );

    \I__11916\ : InMux
    port map (
            O => \N__54747\,
            I => \N__54738\
        );

    \I__11915\ : InMux
    port map (
            O => \N__54746\,
            I => \N__54735\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__54741\,
            I => \N__54732\
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__54738\,
            I => \N__54729\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__54735\,
            I => \N__54726\
        );

    \I__11911\ : Span4Mux_v
    port map (
            O => \N__54732\,
            I => \N__54723\
        );

    \I__11910\ : Span4Mux_h
    port map (
            O => \N__54729\,
            I => \N__54720\
        );

    \I__11909\ : Span4Mux_v
    port map (
            O => \N__54726\,
            I => \N__54716\
        );

    \I__11908\ : Span4Mux_h
    port map (
            O => \N__54723\,
            I => \N__54711\
        );

    \I__11907\ : Span4Mux_v
    port map (
            O => \N__54720\,
            I => \N__54711\
        );

    \I__11906\ : InMux
    port map (
            O => \N__54719\,
            I => \N__54708\
        );

    \I__11905\ : Span4Mux_h
    port map (
            O => \N__54716\,
            I => \N__54702\
        );

    \I__11904\ : Span4Mux_h
    port map (
            O => \N__54711\,
            I => \N__54702\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__54708\,
            I => \N__54699\
        );

    \I__11902\ : InMux
    port map (
            O => \N__54707\,
            I => \N__54696\
        );

    \I__11901\ : Odrv4
    port map (
            O => \N__54702\,
            I => \CONTROL.N_98_0\
        );

    \I__11900\ : Odrv4
    port map (
            O => \N__54699\,
            I => \CONTROL.N_98_0\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__54696\,
            I => \CONTROL.N_98_0\
        );

    \I__11898\ : InMux
    port map (
            O => \N__54689\,
            I => \N__54682\
        );

    \I__11897\ : InMux
    port map (
            O => \N__54688\,
            I => \N__54674\
        );

    \I__11896\ : InMux
    port map (
            O => \N__54687\,
            I => \N__54671\
        );

    \I__11895\ : InMux
    port map (
            O => \N__54686\,
            I => \N__54665\
        );

    \I__11894\ : InMux
    port map (
            O => \N__54685\,
            I => \N__54662\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__54682\,
            I => \N__54648\
        );

    \I__11892\ : InMux
    port map (
            O => \N__54681\,
            I => \N__54641\
        );

    \I__11891\ : InMux
    port map (
            O => \N__54680\,
            I => \N__54641\
        );

    \I__11890\ : InMux
    port map (
            O => \N__54679\,
            I => \N__54641\
        );

    \I__11889\ : InMux
    port map (
            O => \N__54678\,
            I => \N__54636\
        );

    \I__11888\ : InMux
    port map (
            O => \N__54677\,
            I => \N__54636\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__54674\,
            I => \N__54627\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__54671\,
            I => \N__54627\
        );

    \I__11885\ : InMux
    port map (
            O => \N__54670\,
            I => \N__54620\
        );

    \I__11884\ : InMux
    port map (
            O => \N__54669\,
            I => \N__54620\
        );

    \I__11883\ : InMux
    port map (
            O => \N__54668\,
            I => \N__54620\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__54665\,
            I => \N__54615\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__54662\,
            I => \N__54615\
        );

    \I__11880\ : InMux
    port map (
            O => \N__54661\,
            I => \N__54612\
        );

    \I__11879\ : InMux
    port map (
            O => \N__54660\,
            I => \N__54609\
        );

    \I__11878\ : InMux
    port map (
            O => \N__54659\,
            I => \N__54602\
        );

    \I__11877\ : InMux
    port map (
            O => \N__54658\,
            I => \N__54602\
        );

    \I__11876\ : InMux
    port map (
            O => \N__54657\,
            I => \N__54602\
        );

    \I__11875\ : InMux
    port map (
            O => \N__54656\,
            I => \N__54599\
        );

    \I__11874\ : InMux
    port map (
            O => \N__54655\,
            I => \N__54596\
        );

    \I__11873\ : InMux
    port map (
            O => \N__54654\,
            I => \N__54593\
        );

    \I__11872\ : InMux
    port map (
            O => \N__54653\,
            I => \N__54588\
        );

    \I__11871\ : InMux
    port map (
            O => \N__54652\,
            I => \N__54588\
        );

    \I__11870\ : CascadeMux
    port map (
            O => \N__54651\,
            I => \N__54576\
        );

    \I__11869\ : Span4Mux_v
    port map (
            O => \N__54648\,
            I => \N__54563\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__54641\,
            I => \N__54563\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__54636\,
            I => \N__54560\
        );

    \I__11866\ : InMux
    port map (
            O => \N__54635\,
            I => \N__54553\
        );

    \I__11865\ : InMux
    port map (
            O => \N__54634\,
            I => \N__54553\
        );

    \I__11864\ : InMux
    port map (
            O => \N__54633\,
            I => \N__54553\
        );

    \I__11863\ : InMux
    port map (
            O => \N__54632\,
            I => \N__54550\
        );

    \I__11862\ : Span4Mux_h
    port map (
            O => \N__54627\,
            I => \N__54545\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__54620\,
            I => \N__54545\
        );

    \I__11860\ : Span4Mux_h
    port map (
            O => \N__54615\,
            I => \N__54536\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__54612\,
            I => \N__54531\
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__54609\,
            I => \N__54531\
        );

    \I__11857\ : LocalMux
    port map (
            O => \N__54602\,
            I => \N__54528\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__54599\,
            I => \N__54519\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__54596\,
            I => \N__54519\
        );

    \I__11854\ : LocalMux
    port map (
            O => \N__54593\,
            I => \N__54519\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__54588\,
            I => \N__54519\
        );

    \I__11852\ : InMux
    port map (
            O => \N__54587\,
            I => \N__54514\
        );

    \I__11851\ : InMux
    port map (
            O => \N__54586\,
            I => \N__54514\
        );

    \I__11850\ : InMux
    port map (
            O => \N__54585\,
            I => \N__54511\
        );

    \I__11849\ : InMux
    port map (
            O => \N__54584\,
            I => \N__54506\
        );

    \I__11848\ : InMux
    port map (
            O => \N__54583\,
            I => \N__54506\
        );

    \I__11847\ : InMux
    port map (
            O => \N__54582\,
            I => \N__54501\
        );

    \I__11846\ : InMux
    port map (
            O => \N__54581\,
            I => \N__54501\
        );

    \I__11845\ : InMux
    port map (
            O => \N__54580\,
            I => \N__54494\
        );

    \I__11844\ : InMux
    port map (
            O => \N__54579\,
            I => \N__54494\
        );

    \I__11843\ : InMux
    port map (
            O => \N__54576\,
            I => \N__54494\
        );

    \I__11842\ : InMux
    port map (
            O => \N__54575\,
            I => \N__54491\
        );

    \I__11841\ : InMux
    port map (
            O => \N__54574\,
            I => \N__54486\
        );

    \I__11840\ : InMux
    port map (
            O => \N__54573\,
            I => \N__54486\
        );

    \I__11839\ : InMux
    port map (
            O => \N__54572\,
            I => \N__54477\
        );

    \I__11838\ : InMux
    port map (
            O => \N__54571\,
            I => \N__54477\
        );

    \I__11837\ : InMux
    port map (
            O => \N__54570\,
            I => \N__54477\
        );

    \I__11836\ : InMux
    port map (
            O => \N__54569\,
            I => \N__54477\
        );

    \I__11835\ : InMux
    port map (
            O => \N__54568\,
            I => \N__54474\
        );

    \I__11834\ : Span4Mux_h
    port map (
            O => \N__54563\,
            I => \N__54469\
        );

    \I__11833\ : Span4Mux_v
    port map (
            O => \N__54560\,
            I => \N__54469\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__54553\,
            I => \N__54466\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__54550\,
            I => \N__54461\
        );

    \I__11830\ : Span4Mux_h
    port map (
            O => \N__54545\,
            I => \N__54461\
        );

    \I__11829\ : InMux
    port map (
            O => \N__54544\,
            I => \N__54458\
        );

    \I__11828\ : InMux
    port map (
            O => \N__54543\,
            I => \N__54453\
        );

    \I__11827\ : InMux
    port map (
            O => \N__54542\,
            I => \N__54453\
        );

    \I__11826\ : InMux
    port map (
            O => \N__54541\,
            I => \N__54446\
        );

    \I__11825\ : InMux
    port map (
            O => \N__54540\,
            I => \N__54446\
        );

    \I__11824\ : InMux
    port map (
            O => \N__54539\,
            I => \N__54446\
        );

    \I__11823\ : Span4Mux_v
    port map (
            O => \N__54536\,
            I => \N__54435\
        );

    \I__11822\ : Span4Mux_v
    port map (
            O => \N__54531\,
            I => \N__54435\
        );

    \I__11821\ : Span4Mux_h
    port map (
            O => \N__54528\,
            I => \N__54435\
        );

    \I__11820\ : Span4Mux_v
    port map (
            O => \N__54519\,
            I => \N__54435\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__54514\,
            I => \N__54435\
        );

    \I__11818\ : LocalMux
    port map (
            O => \N__54511\,
            I => \N__54426\
        );

    \I__11817\ : LocalMux
    port map (
            O => \N__54506\,
            I => \N__54426\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__54501\,
            I => \N__54426\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__54494\,
            I => \N__54426\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__54491\,
            I => \controlWord_4\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__54486\,
            I => \controlWord_4\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__54477\,
            I => \controlWord_4\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__54474\,
            I => \controlWord_4\
        );

    \I__11810\ : Odrv4
    port map (
            O => \N__54469\,
            I => \controlWord_4\
        );

    \I__11809\ : Odrv4
    port map (
            O => \N__54466\,
            I => \controlWord_4\
        );

    \I__11808\ : Odrv4
    port map (
            O => \N__54461\,
            I => \controlWord_4\
        );

    \I__11807\ : LocalMux
    port map (
            O => \N__54458\,
            I => \controlWord_4\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__54453\,
            I => \controlWord_4\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__54446\,
            I => \controlWord_4\
        );

    \I__11804\ : Odrv4
    port map (
            O => \N__54435\,
            I => \controlWord_4\
        );

    \I__11803\ : Odrv4
    port map (
            O => \N__54426\,
            I => \controlWord_4\
        );

    \I__11802\ : InMux
    port map (
            O => \N__54401\,
            I => \N__54398\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__54398\,
            I => \PROM.ROMDATA.m320_am\
        );

    \I__11800\ : InMux
    port map (
            O => \N__54395\,
            I => \N__54392\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__54392\,
            I => \PROM.ROMDATA.m150\
        );

    \I__11798\ : CascadeMux
    port map (
            O => \N__54389\,
            I => \N__54386\
        );

    \I__11797\ : InMux
    port map (
            O => \N__54386\,
            I => \N__54383\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__54383\,
            I => \N__54380\
        );

    \I__11795\ : Span12Mux_v
    port map (
            O => \N__54380\,
            I => \N__54377\
        );

    \I__11794\ : Odrv12
    port map (
            O => \N__54377\,
            I => \PROM.ROMDATA.N_558_mux\
        );

    \I__11793\ : CascadeMux
    port map (
            O => \N__54374\,
            I => \PROM.ROMDATA.m49_cascade_\
        );

    \I__11792\ : InMux
    port map (
            O => \N__54371\,
            I => \N__54368\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__54368\,
            I => \PROM.ROMDATA.m229_1\
        );

    \I__11790\ : CascadeMux
    port map (
            O => \N__54365\,
            I => \PROM.ROMDATA.m228_bm_cascade_\
        );

    \I__11789\ : InMux
    port map (
            O => \N__54362\,
            I => \N__54359\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__54359\,
            I => \N__54352\
        );

    \I__11787\ : InMux
    port map (
            O => \N__54358\,
            I => \N__54343\
        );

    \I__11786\ : InMux
    port map (
            O => \N__54357\,
            I => \N__54343\
        );

    \I__11785\ : InMux
    port map (
            O => \N__54356\,
            I => \N__54343\
        );

    \I__11784\ : InMux
    port map (
            O => \N__54355\,
            I => \N__54343\
        );

    \I__11783\ : Span4Mux_h
    port map (
            O => \N__54352\,
            I => \N__54338\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__54343\,
            I => \N__54338\
        );

    \I__11781\ : Span4Mux_h
    port map (
            O => \N__54338\,
            I => \N__54335\
        );

    \I__11780\ : Span4Mux_h
    port map (
            O => \N__54335\,
            I => \N__54332\
        );

    \I__11779\ : Odrv4
    port map (
            O => \N__54332\,
            I => \PROM.ROMDATA.m229\
        );

    \I__11778\ : InMux
    port map (
            O => \N__54329\,
            I => \N__54323\
        );

    \I__11777\ : InMux
    port map (
            O => \N__54328\,
            I => \N__54323\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__54323\,
            I => \N__54320\
        );

    \I__11775\ : Odrv12
    port map (
            O => \N__54320\,
            I => \ALU.dZ0Z_15\
        );

    \I__11774\ : InMux
    port map (
            O => \N__54317\,
            I => \N__54314\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__54314\,
            I => \N__54311\
        );

    \I__11772\ : Odrv12
    port map (
            O => \N__54311\,
            I => \ALU.dout_6_ns_1_15\
        );

    \I__11771\ : CascadeMux
    port map (
            O => \N__54308\,
            I => \N__54305\
        );

    \I__11770\ : InMux
    port map (
            O => \N__54305\,
            I => \N__54300\
        );

    \I__11769\ : InMux
    port map (
            O => \N__54304\,
            I => \N__54289\
        );

    \I__11768\ : InMux
    port map (
            O => \N__54303\,
            I => \N__54286\
        );

    \I__11767\ : LocalMux
    port map (
            O => \N__54300\,
            I => \N__54281\
        );

    \I__11766\ : InMux
    port map (
            O => \N__54299\,
            I => \N__54276\
        );

    \I__11765\ : InMux
    port map (
            O => \N__54298\,
            I => \N__54276\
        );

    \I__11764\ : InMux
    port map (
            O => \N__54297\,
            I => \N__54271\
        );

    \I__11763\ : InMux
    port map (
            O => \N__54296\,
            I => \N__54271\
        );

    \I__11762\ : InMux
    port map (
            O => \N__54295\,
            I => \N__54266\
        );

    \I__11761\ : InMux
    port map (
            O => \N__54294\,
            I => \N__54266\
        );

    \I__11760\ : InMux
    port map (
            O => \N__54293\,
            I => \N__54261\
        );

    \I__11759\ : InMux
    port map (
            O => \N__54292\,
            I => \N__54261\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__54289\,
            I => \N__54258\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__54286\,
            I => \N__54255\
        );

    \I__11756\ : InMux
    port map (
            O => \N__54285\,
            I => \N__54250\
        );

    \I__11755\ : InMux
    port map (
            O => \N__54284\,
            I => \N__54250\
        );

    \I__11754\ : Span4Mux_h
    port map (
            O => \N__54281\,
            I => \N__54244\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__54276\,
            I => \N__54244\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__54271\,
            I => \N__54237\
        );

    \I__11751\ : LocalMux
    port map (
            O => \N__54266\,
            I => \N__54237\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__54261\,
            I => \N__54237\
        );

    \I__11749\ : Span4Mux_h
    port map (
            O => \N__54258\,
            I => \N__54231\
        );

    \I__11748\ : Span4Mux_h
    port map (
            O => \N__54255\,
            I => \N__54228\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__54250\,
            I => \N__54225\
        );

    \I__11746\ : InMux
    port map (
            O => \N__54249\,
            I => \N__54222\
        );

    \I__11745\ : Span4Mux_h
    port map (
            O => \N__54244\,
            I => \N__54217\
        );

    \I__11744\ : Span4Mux_h
    port map (
            O => \N__54237\,
            I => \N__54217\
        );

    \I__11743\ : InMux
    port map (
            O => \N__54236\,
            I => \N__54212\
        );

    \I__11742\ : InMux
    port map (
            O => \N__54235\,
            I => \N__54212\
        );

    \I__11741\ : InMux
    port map (
            O => \N__54234\,
            I => \N__54209\
        );

    \I__11740\ : Odrv4
    port map (
            O => \N__54231\,
            I => \aluOperand1_1_rep2\
        );

    \I__11739\ : Odrv4
    port map (
            O => \N__54228\,
            I => \aluOperand1_1_rep2\
        );

    \I__11738\ : Odrv4
    port map (
            O => \N__54225\,
            I => \aluOperand1_1_rep2\
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__54222\,
            I => \aluOperand1_1_rep2\
        );

    \I__11736\ : Odrv4
    port map (
            O => \N__54217\,
            I => \aluOperand1_1_rep2\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__54212\,
            I => \aluOperand1_1_rep2\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__54209\,
            I => \aluOperand1_1_rep2\
        );

    \I__11733\ : InMux
    port map (
            O => \N__54194\,
            I => \N__54191\
        );

    \I__11732\ : LocalMux
    port map (
            O => \N__54191\,
            I => \N__54188\
        );

    \I__11731\ : Span12Mux_v
    port map (
            O => \N__54188\,
            I => \N__54183\
        );

    \I__11730\ : InMux
    port map (
            O => \N__54187\,
            I => \N__54178\
        );

    \I__11729\ : InMux
    port map (
            O => \N__54186\,
            I => \N__54178\
        );

    \I__11728\ : Span12Mux_v
    port map (
            O => \N__54183\,
            I => \N__54175\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__54178\,
            I => \N__54172\
        );

    \I__11726\ : Span12Mux_h
    port map (
            O => \N__54175\,
            I => \N__54169\
        );

    \I__11725\ : Span4Mux_v
    port map (
            O => \N__54172\,
            I => \N__54166\
        );

    \I__11724\ : Odrv12
    port map (
            O => \N__54169\,
            I => h_15
        );

    \I__11723\ : Odrv4
    port map (
            O => \N__54166\,
            I => h_15
        );

    \I__11722\ : InMux
    port map (
            O => \N__54161\,
            I => \N__54158\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__54158\,
            I => \N__54155\
        );

    \I__11720\ : Span4Mux_h
    port map (
            O => \N__54155\,
            I => \N__54152\
        );

    \I__11719\ : Span4Mux_h
    port map (
            O => \N__54152\,
            I => \N__54149\
        );

    \I__11718\ : Odrv4
    port map (
            O => \N__54149\,
            I => \ALU.N_1100\
        );

    \I__11717\ : CascadeMux
    port map (
            O => \N__54146\,
            I => \ALU.N_1148_cascade_\
        );

    \I__11716\ : InMux
    port map (
            O => \N__54143\,
            I => \N__54135\
        );

    \I__11715\ : InMux
    port map (
            O => \N__54142\,
            I => \N__54131\
        );

    \I__11714\ : InMux
    port map (
            O => \N__54141\,
            I => \N__54125\
        );

    \I__11713\ : InMux
    port map (
            O => \N__54140\,
            I => \N__54122\
        );

    \I__11712\ : InMux
    port map (
            O => \N__54139\,
            I => \N__54119\
        );

    \I__11711\ : InMux
    port map (
            O => \N__54138\,
            I => \N__54115\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__54135\,
            I => \N__54107\
        );

    \I__11709\ : InMux
    port map (
            O => \N__54134\,
            I => \N__54104\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__54131\,
            I => \N__54101\
        );

    \I__11707\ : InMux
    port map (
            O => \N__54130\,
            I => \N__54098\
        );

    \I__11706\ : InMux
    port map (
            O => \N__54129\,
            I => \N__54093\
        );

    \I__11705\ : InMux
    port map (
            O => \N__54128\,
            I => \N__54093\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__54125\,
            I => \N__54090\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__54122\,
            I => \N__54085\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__54119\,
            I => \N__54085\
        );

    \I__11701\ : InMux
    port map (
            O => \N__54118\,
            I => \N__54082\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__54115\,
            I => \N__54079\
        );

    \I__11699\ : InMux
    port map (
            O => \N__54114\,
            I => \N__54074\
        );

    \I__11698\ : InMux
    port map (
            O => \N__54113\,
            I => \N__54074\
        );

    \I__11697\ : InMux
    port map (
            O => \N__54112\,
            I => \N__54069\
        );

    \I__11696\ : InMux
    port map (
            O => \N__54111\,
            I => \N__54069\
        );

    \I__11695\ : InMux
    port map (
            O => \N__54110\,
            I => \N__54066\
        );

    \I__11694\ : Span4Mux_h
    port map (
            O => \N__54107\,
            I => \N__54063\
        );

    \I__11693\ : LocalMux
    port map (
            O => \N__54104\,
            I => \N__54056\
        );

    \I__11692\ : Span4Mux_v
    port map (
            O => \N__54101\,
            I => \N__54047\
        );

    \I__11691\ : LocalMux
    port map (
            O => \N__54098\,
            I => \N__54047\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__54093\,
            I => \N__54047\
        );

    \I__11689\ : Span4Mux_h
    port map (
            O => \N__54090\,
            I => \N__54047\
        );

    \I__11688\ : Span4Mux_h
    port map (
            O => \N__54085\,
            I => \N__54042\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__54082\,
            I => \N__54042\
        );

    \I__11686\ : Span4Mux_v
    port map (
            O => \N__54079\,
            I => \N__54034\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__54074\,
            I => \N__54034\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__54069\,
            I => \N__54034\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__54066\,
            I => \N__54029\
        );

    \I__11682\ : Span4Mux_v
    port map (
            O => \N__54063\,
            I => \N__54029\
        );

    \I__11681\ : InMux
    port map (
            O => \N__54062\,
            I => \N__54022\
        );

    \I__11680\ : InMux
    port map (
            O => \N__54061\,
            I => \N__54022\
        );

    \I__11679\ : InMux
    port map (
            O => \N__54060\,
            I => \N__54022\
        );

    \I__11678\ : InMux
    port map (
            O => \N__54059\,
            I => \N__54019\
        );

    \I__11677\ : Span4Mux_v
    port map (
            O => \N__54056\,
            I => \N__54012\
        );

    \I__11676\ : Span4Mux_h
    port map (
            O => \N__54047\,
            I => \N__54012\
        );

    \I__11675\ : Span4Mux_h
    port map (
            O => \N__54042\,
            I => \N__54012\
        );

    \I__11674\ : InMux
    port map (
            O => \N__54041\,
            I => \N__54009\
        );

    \I__11673\ : Span4Mux_h
    port map (
            O => \N__54034\,
            I => \N__54006\
        );

    \I__11672\ : Span4Mux_v
    port map (
            O => \N__54029\,
            I => \N__54001\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__54022\,
            I => \N__54001\
        );

    \I__11670\ : LocalMux
    port map (
            O => \N__54019\,
            I => \aluOperand1_0\
        );

    \I__11669\ : Odrv4
    port map (
            O => \N__54012\,
            I => \aluOperand1_0\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__54009\,
            I => \aluOperand1_0\
        );

    \I__11667\ : Odrv4
    port map (
            O => \N__54006\,
            I => \aluOperand1_0\
        );

    \I__11666\ : Odrv4
    port map (
            O => \N__54001\,
            I => \aluOperand1_0\
        );

    \I__11665\ : InMux
    port map (
            O => \N__53990\,
            I => \N__53987\
        );

    \I__11664\ : LocalMux
    port map (
            O => \N__53987\,
            I => \ALU.N_1260\
        );

    \I__11663\ : InMux
    port map (
            O => \N__53984\,
            I => \N__53981\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__53981\,
            I => \N__53978\
        );

    \I__11661\ : Span4Mux_h
    port map (
            O => \N__53978\,
            I => \N__53975\
        );

    \I__11660\ : Span4Mux_h
    port map (
            O => \N__53975\,
            I => \N__53972\
        );

    \I__11659\ : Odrv4
    port map (
            O => \N__53972\,
            I => \ALU.N_1212\
        );

    \I__11658\ : CascadeMux
    port map (
            O => \N__53969\,
            I => \N__53958\
        );

    \I__11657\ : InMux
    port map (
            O => \N__53968\,
            I => \N__53953\
        );

    \I__11656\ : InMux
    port map (
            O => \N__53967\,
            I => \N__53946\
        );

    \I__11655\ : InMux
    port map (
            O => \N__53966\,
            I => \N__53946\
        );

    \I__11654\ : InMux
    port map (
            O => \N__53965\,
            I => \N__53943\
        );

    \I__11653\ : InMux
    port map (
            O => \N__53964\,
            I => \N__53931\
        );

    \I__11652\ : InMux
    port map (
            O => \N__53963\,
            I => \N__53931\
        );

    \I__11651\ : InMux
    port map (
            O => \N__53962\,
            I => \N__53924\
        );

    \I__11650\ : InMux
    port map (
            O => \N__53961\,
            I => \N__53924\
        );

    \I__11649\ : InMux
    port map (
            O => \N__53958\,
            I => \N__53924\
        );

    \I__11648\ : InMux
    port map (
            O => \N__53957\,
            I => \N__53919\
        );

    \I__11647\ : InMux
    port map (
            O => \N__53956\,
            I => \N__53919\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__53953\,
            I => \N__53916\
        );

    \I__11645\ : InMux
    port map (
            O => \N__53952\,
            I => \N__53911\
        );

    \I__11644\ : InMux
    port map (
            O => \N__53951\,
            I => \N__53911\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__53946\,
            I => \N__53904\
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__53943\,
            I => \N__53904\
        );

    \I__11641\ : InMux
    port map (
            O => \N__53942\,
            I => \N__53899\
        );

    \I__11640\ : InMux
    port map (
            O => \N__53941\,
            I => \N__53899\
        );

    \I__11639\ : CascadeMux
    port map (
            O => \N__53940\,
            I => \N__53895\
        );

    \I__11638\ : InMux
    port map (
            O => \N__53939\,
            I => \N__53890\
        );

    \I__11637\ : InMux
    port map (
            O => \N__53938\,
            I => \N__53890\
        );

    \I__11636\ : InMux
    port map (
            O => \N__53937\,
            I => \N__53882\
        );

    \I__11635\ : InMux
    port map (
            O => \N__53936\,
            I => \N__53882\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__53931\,
            I => \N__53879\
        );

    \I__11633\ : LocalMux
    port map (
            O => \N__53924\,
            I => \N__53876\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__53919\,
            I => \N__53873\
        );

    \I__11631\ : Span4Mux_v
    port map (
            O => \N__53916\,
            I => \N__53870\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__53911\,
            I => \N__53867\
        );

    \I__11629\ : InMux
    port map (
            O => \N__53910\,
            I => \N__53862\
        );

    \I__11628\ : InMux
    port map (
            O => \N__53909\,
            I => \N__53862\
        );

    \I__11627\ : Span4Mux_h
    port map (
            O => \N__53904\,
            I => \N__53856\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__53899\,
            I => \N__53853\
        );

    \I__11625\ : InMux
    port map (
            O => \N__53898\,
            I => \N__53848\
        );

    \I__11624\ : InMux
    port map (
            O => \N__53895\,
            I => \N__53848\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__53890\,
            I => \N__53845\
        );

    \I__11622\ : InMux
    port map (
            O => \N__53889\,
            I => \N__53842\
        );

    \I__11621\ : InMux
    port map (
            O => \N__53888\,
            I => \N__53837\
        );

    \I__11620\ : InMux
    port map (
            O => \N__53887\,
            I => \N__53837\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__53882\,
            I => \N__53828\
        );

    \I__11618\ : Span4Mux_v
    port map (
            O => \N__53879\,
            I => \N__53828\
        );

    \I__11617\ : Span4Mux_h
    port map (
            O => \N__53876\,
            I => \N__53828\
        );

    \I__11616\ : Span4Mux_v
    port map (
            O => \N__53873\,
            I => \N__53828\
        );

    \I__11615\ : Span4Mux_h
    port map (
            O => \N__53870\,
            I => \N__53823\
        );

    \I__11614\ : Span4Mux_v
    port map (
            O => \N__53867\,
            I => \N__53823\
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__53862\,
            I => \N__53820\
        );

    \I__11612\ : InMux
    port map (
            O => \N__53861\,
            I => \N__53817\
        );

    \I__11611\ : InMux
    port map (
            O => \N__53860\,
            I => \N__53812\
        );

    \I__11610\ : InMux
    port map (
            O => \N__53859\,
            I => \N__53812\
        );

    \I__11609\ : Span4Mux_h
    port map (
            O => \N__53856\,
            I => \N__53805\
        );

    \I__11608\ : Span4Mux_h
    port map (
            O => \N__53853\,
            I => \N__53805\
        );

    \I__11607\ : LocalMux
    port map (
            O => \N__53848\,
            I => \N__53805\
        );

    \I__11606\ : Span4Mux_h
    port map (
            O => \N__53845\,
            I => \N__53796\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__53842\,
            I => \N__53796\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__53837\,
            I => \N__53796\
        );

    \I__11603\ : Span4Mux_h
    port map (
            O => \N__53828\,
            I => \N__53796\
        );

    \I__11602\ : Odrv4
    port map (
            O => \N__53823\,
            I => \aluOperand2_0\
        );

    \I__11601\ : Odrv12
    port map (
            O => \N__53820\,
            I => \aluOperand2_0\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__53817\,
            I => \aluOperand2_0\
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__53812\,
            I => \aluOperand2_0\
        );

    \I__11598\ : Odrv4
    port map (
            O => \N__53805\,
            I => \aluOperand2_0\
        );

    \I__11597\ : Odrv4
    port map (
            O => \N__53796\,
            I => \aluOperand2_0\
        );

    \I__11596\ : InMux
    port map (
            O => \N__53783\,
            I => \N__53780\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__53780\,
            I => \N__53777\
        );

    \I__11594\ : Span4Mux_v
    port map (
            O => \N__53777\,
            I => \N__53774\
        );

    \I__11593\ : Sp12to4
    port map (
            O => \N__53774\,
            I => \N__53771\
        );

    \I__11592\ : Span12Mux_h
    port map (
            O => \N__53771\,
            I => \N__53768\
        );

    \I__11591\ : Odrv12
    port map (
            O => \N__53768\,
            I => \ALU.combOperand2_d_bmZ0Z_15\
        );

    \I__11590\ : CascadeMux
    port map (
            O => \N__53765\,
            I => \ALU.c_RNI8VV95Z0Z_15_cascade_\
        );

    \I__11589\ : InMux
    port map (
            O => \N__53762\,
            I => \N__53759\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__53759\,
            I => \N__53754\
        );

    \I__11587\ : InMux
    port map (
            O => \N__53758\,
            I => \N__53749\
        );

    \I__11586\ : InMux
    port map (
            O => \N__53757\,
            I => \N__53749\
        );

    \I__11585\ : Odrv4
    port map (
            O => \N__53754\,
            I => \ALU.c_RNIJTKD7Z0Z_15\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__53749\,
            I => \ALU.c_RNIJTKD7Z0Z_15\
        );

    \I__11583\ : CascadeMux
    port map (
            O => \N__53744\,
            I => \PROM.ROMDATA.m320_bm_cascade_\
        );

    \I__11582\ : InMux
    port map (
            O => \N__53741\,
            I => \N__53738\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__53738\,
            I => \PROM.ROMDATA.m410_am\
        );

    \I__11580\ : CascadeMux
    port map (
            O => \N__53735\,
            I => \PROM.ROMDATA.m413_am_cascade_\
        );

    \I__11579\ : CascadeMux
    port map (
            O => \N__53732\,
            I => \ALU.status_e_0_RNO_0Z0Z_2_cascade_\
        );

    \I__11578\ : CascadeMux
    port map (
            O => \N__53729\,
            I => \ALU.N_570_cascade_\
        );

    \I__11577\ : InMux
    port map (
            O => \N__53726\,
            I => \N__53723\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__53723\,
            I => \ALU.status_e_0_RNO_1Z0Z_2\
        );

    \I__11575\ : InMux
    port map (
            O => \N__53720\,
            I => \N__53714\
        );

    \I__11574\ : InMux
    port map (
            O => \N__53719\,
            I => \N__53709\
        );

    \I__11573\ : InMux
    port map (
            O => \N__53718\,
            I => \N__53709\
        );

    \I__11572\ : CascadeMux
    port map (
            O => \N__53717\,
            I => \N__53706\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__53714\,
            I => \N__53701\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__53709\,
            I => \N__53698\
        );

    \I__11569\ : InMux
    port map (
            O => \N__53706\,
            I => \N__53691\
        );

    \I__11568\ : InMux
    port map (
            O => \N__53705\,
            I => \N__53691\
        );

    \I__11567\ : InMux
    port map (
            O => \N__53704\,
            I => \N__53691\
        );

    \I__11566\ : Span4Mux_v
    port map (
            O => \N__53701\,
            I => \N__53682\
        );

    \I__11565\ : Span4Mux_v
    port map (
            O => \N__53698\,
            I => \N__53682\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__53691\,
            I => \N__53682\
        );

    \I__11563\ : InMux
    port map (
            O => \N__53690\,
            I => \N__53677\
        );

    \I__11562\ : InMux
    port map (
            O => \N__53689\,
            I => \N__53677\
        );

    \I__11561\ : Span4Mux_v
    port map (
            O => \N__53682\,
            I => \N__53674\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__53677\,
            I => \aluStatus_2\
        );

    \I__11559\ : Odrv4
    port map (
            O => \N__53674\,
            I => \aluStatus_2\
        );

    \I__11558\ : InMux
    port map (
            O => \N__53669\,
            I => \N__53663\
        );

    \I__11557\ : InMux
    port map (
            O => \N__53668\,
            I => \N__53658\
        );

    \I__11556\ : InMux
    port map (
            O => \N__53667\,
            I => \N__53653\
        );

    \I__11555\ : InMux
    port map (
            O => \N__53666\,
            I => \N__53653\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__53663\,
            I => \N__53650\
        );

    \I__11553\ : InMux
    port map (
            O => \N__53662\,
            I => \N__53645\
        );

    \I__11552\ : InMux
    port map (
            O => \N__53661\,
            I => \N__53645\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__53658\,
            I => \N__53642\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__53653\,
            I => \N__53639\
        );

    \I__11549\ : Span4Mux_h
    port map (
            O => \N__53650\,
            I => \N__53636\
        );

    \I__11548\ : LocalMux
    port map (
            O => \N__53645\,
            I => \PROM_ROMDATA_dintern_9ro\
        );

    \I__11547\ : Odrv12
    port map (
            O => \N__53642\,
            I => \PROM_ROMDATA_dintern_9ro\
        );

    \I__11546\ : Odrv4
    port map (
            O => \N__53639\,
            I => \PROM_ROMDATA_dintern_9ro\
        );

    \I__11545\ : Odrv4
    port map (
            O => \N__53636\,
            I => \PROM_ROMDATA_dintern_9ro\
        );

    \I__11544\ : InMux
    port map (
            O => \N__53627\,
            I => \N__53624\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__53624\,
            I => \N__53621\
        );

    \I__11542\ : Span4Mux_v
    port map (
            O => \N__53621\,
            I => \N__53618\
        );

    \I__11541\ : Span4Mux_h
    port map (
            O => \N__53618\,
            I => \N__53615\
        );

    \I__11540\ : Odrv4
    port map (
            O => \N__53615\,
            I => \CONTROL.g3Z0Z_0\
        );

    \I__11539\ : InMux
    port map (
            O => \N__53612\,
            I => \N__53608\
        );

    \I__11538\ : InMux
    port map (
            O => \N__53611\,
            I => \N__53605\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__53608\,
            I => \N__53602\
        );

    \I__11536\ : LocalMux
    port map (
            O => \N__53605\,
            I => \N__53599\
        );

    \I__11535\ : Span12Mux_h
    port map (
            O => \N__53602\,
            I => \N__53596\
        );

    \I__11534\ : Span4Mux_v
    port map (
            O => \N__53599\,
            I => \N__53593\
        );

    \I__11533\ : Odrv12
    port map (
            O => \N__53596\,
            I => \ALU.bZ0Z_15\
        );

    \I__11532\ : Odrv4
    port map (
            O => \N__53593\,
            I => \ALU.bZ0Z_15\
        );

    \I__11531\ : InMux
    port map (
            O => \N__53588\,
            I => \N__53585\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__53585\,
            I => \N__53580\
        );

    \I__11529\ : InMux
    port map (
            O => \N__53584\,
            I => \N__53575\
        );

    \I__11528\ : InMux
    port map (
            O => \N__53583\,
            I => \N__53575\
        );

    \I__11527\ : Span4Mux_v
    port map (
            O => \N__53580\,
            I => \N__53567\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__53575\,
            I => \N__53564\
        );

    \I__11525\ : InMux
    port map (
            O => \N__53574\,
            I => \N__53561\
        );

    \I__11524\ : InMux
    port map (
            O => \N__53573\,
            I => \N__53558\
        );

    \I__11523\ : InMux
    port map (
            O => \N__53572\,
            I => \N__53555\
        );

    \I__11522\ : InMux
    port map (
            O => \N__53571\,
            I => \N__53550\
        );

    \I__11521\ : InMux
    port map (
            O => \N__53570\,
            I => \N__53550\
        );

    \I__11520\ : Span4Mux_h
    port map (
            O => \N__53567\,
            I => \N__53545\
        );

    \I__11519\ : Span4Mux_v
    port map (
            O => \N__53564\,
            I => \N__53545\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__53561\,
            I => \aluOperand2_fast_2\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__53558\,
            I => \aluOperand2_fast_2\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__53555\,
            I => \aluOperand2_fast_2\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__53550\,
            I => \aluOperand2_fast_2\
        );

    \I__11514\ : Odrv4
    port map (
            O => \N__53545\,
            I => \aluOperand2_fast_2\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__53534\,
            I => \N__53531\
        );

    \I__11512\ : InMux
    port map (
            O => \N__53531\,
            I => \N__53527\
        );

    \I__11511\ : CascadeMux
    port map (
            O => \N__53530\,
            I => \N__53524\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__53527\,
            I => \N__53521\
        );

    \I__11509\ : InMux
    port map (
            O => \N__53524\,
            I => \N__53518\
        );

    \I__11508\ : Span4Mux_h
    port map (
            O => \N__53521\,
            I => \N__53514\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__53518\,
            I => \N__53511\
        );

    \I__11506\ : CascadeMux
    port map (
            O => \N__53517\,
            I => \N__53508\
        );

    \I__11505\ : Span4Mux_v
    port map (
            O => \N__53514\,
            I => \N__53505\
        );

    \I__11504\ : Span4Mux_v
    port map (
            O => \N__53511\,
            I => \N__53502\
        );

    \I__11503\ : InMux
    port map (
            O => \N__53508\,
            I => \N__53499\
        );

    \I__11502\ : Sp12to4
    port map (
            O => \N__53505\,
            I => \N__53496\
        );

    \I__11501\ : Sp12to4
    port map (
            O => \N__53502\,
            I => \N__53493\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__53499\,
            I => \N__53490\
        );

    \I__11499\ : Span12Mux_v
    port map (
            O => \N__53496\,
            I => \N__53485\
        );

    \I__11498\ : Span12Mux_h
    port map (
            O => \N__53493\,
            I => \N__53485\
        );

    \I__11497\ : Odrv4
    port map (
            O => \N__53490\,
            I => f_15
        );

    \I__11496\ : Odrv12
    port map (
            O => \N__53485\,
            I => f_15
        );

    \I__11495\ : InMux
    port map (
            O => \N__53480\,
            I => \N__53474\
        );

    \I__11494\ : InMux
    port map (
            O => \N__53479\,
            I => \N__53471\
        );

    \I__11493\ : InMux
    port map (
            O => \N__53478\,
            I => \N__53468\
        );

    \I__11492\ : InMux
    port map (
            O => \N__53477\,
            I => \N__53463\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__53474\,
            I => \N__53458\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__53471\,
            I => \N__53458\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__53468\,
            I => \N__53455\
        );

    \I__11488\ : InMux
    port map (
            O => \N__53467\,
            I => \N__53450\
        );

    \I__11487\ : InMux
    port map (
            O => \N__53466\,
            I => \N__53450\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__53463\,
            I => \N__53445\
        );

    \I__11485\ : Span4Mux_v
    port map (
            O => \N__53458\,
            I => \N__53445\
        );

    \I__11484\ : Odrv12
    port map (
            O => \N__53455\,
            I => \aluOperand2_fast_1\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__53450\,
            I => \aluOperand2_fast_1\
        );

    \I__11482\ : Odrv4
    port map (
            O => \N__53445\,
            I => \aluOperand2_fast_1\
        );

    \I__11481\ : CascadeMux
    port map (
            O => \N__53438\,
            I => \ALU.operand2_6_ns_1_15_cascade_\
        );

    \I__11480\ : InMux
    port map (
            O => \N__53435\,
            I => \N__53431\
        );

    \I__11479\ : InMux
    port map (
            O => \N__53434\,
            I => \N__53426\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__53431\,
            I => \N__53422\
        );

    \I__11477\ : InMux
    port map (
            O => \N__53430\,
            I => \N__53417\
        );

    \I__11476\ : InMux
    port map (
            O => \N__53429\,
            I => \N__53417\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__53426\,
            I => \N__53414\
        );

    \I__11474\ : InMux
    port map (
            O => \N__53425\,
            I => \N__53411\
        );

    \I__11473\ : Span4Mux_h
    port map (
            O => \N__53422\,
            I => \N__53407\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__53417\,
            I => \N__53402\
        );

    \I__11471\ : Span4Mux_h
    port map (
            O => \N__53414\,
            I => \N__53395\
        );

    \I__11470\ : LocalMux
    port map (
            O => \N__53411\,
            I => \N__53395\
        );

    \I__11469\ : InMux
    port map (
            O => \N__53410\,
            I => \N__53392\
        );

    \I__11468\ : Span4Mux_h
    port map (
            O => \N__53407\,
            I => \N__53389\
        );

    \I__11467\ : InMux
    port map (
            O => \N__53406\,
            I => \N__53384\
        );

    \I__11466\ : InMux
    port map (
            O => \N__53405\,
            I => \N__53384\
        );

    \I__11465\ : Span4Mux_h
    port map (
            O => \N__53402\,
            I => \N__53381\
        );

    \I__11464\ : InMux
    port map (
            O => \N__53401\,
            I => \N__53376\
        );

    \I__11463\ : InMux
    port map (
            O => \N__53400\,
            I => \N__53376\
        );

    \I__11462\ : Odrv4
    port map (
            O => \N__53395\,
            I => \aluOperand2_1_rep1\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__53392\,
            I => \aluOperand2_1_rep1\
        );

    \I__11460\ : Odrv4
    port map (
            O => \N__53389\,
            I => \aluOperand2_1_rep1\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__53384\,
            I => \aluOperand2_1_rep1\
        );

    \I__11458\ : Odrv4
    port map (
            O => \N__53381\,
            I => \aluOperand2_1_rep1\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__53376\,
            I => \aluOperand2_1_rep1\
        );

    \I__11456\ : CascadeMux
    port map (
            O => \N__53363\,
            I => \ALU.status_14_0_0_cascade_\
        );

    \I__11455\ : CascadeMux
    port map (
            O => \N__53360\,
            I => \N__53357\
        );

    \I__11454\ : InMux
    port map (
            O => \N__53357\,
            I => \N__53354\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__53354\,
            I => \N__53351\
        );

    \I__11452\ : Span4Mux_v
    port map (
            O => \N__53351\,
            I => \N__53348\
        );

    \I__11451\ : Odrv4
    port map (
            O => \N__53348\,
            I => \ALU.status_14_5_0\
        );

    \I__11450\ : CascadeMux
    port map (
            O => \N__53345\,
            I => \ALU.status_14_7_0_cascade_\
        );

    \I__11449\ : InMux
    port map (
            O => \N__53342\,
            I => \N__53339\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__53339\,
            I => \N__53336\
        );

    \I__11447\ : Odrv4
    port map (
            O => \N__53336\,
            I => \ALU.status_14_13_0\
        );

    \I__11446\ : InMux
    port map (
            O => \N__53333\,
            I => \N__53329\
        );

    \I__11445\ : InMux
    port map (
            O => \N__53332\,
            I => \N__53326\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__53329\,
            I => \N__53323\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__53326\,
            I => \N__53320\
        );

    \I__11442\ : Span4Mux_h
    port map (
            O => \N__53323\,
            I => \N__53317\
        );

    \I__11441\ : Span4Mux_v
    port map (
            O => \N__53320\,
            I => \N__53314\
        );

    \I__11440\ : Odrv4
    port map (
            O => \N__53317\,
            I => \ALU.N_979\
        );

    \I__11439\ : Odrv4
    port map (
            O => \N__53314\,
            I => \ALU.N_979\
        );

    \I__11438\ : CascadeMux
    port map (
            O => \N__53309\,
            I => \ALU.N_979_cascade_\
        );

    \I__11437\ : InMux
    port map (
            O => \N__53306\,
            I => \N__53285\
        );

    \I__11436\ : InMux
    port map (
            O => \N__53305\,
            I => \N__53282\
        );

    \I__11435\ : InMux
    port map (
            O => \N__53304\,
            I => \N__53275\
        );

    \I__11434\ : InMux
    port map (
            O => \N__53303\,
            I => \N__53275\
        );

    \I__11433\ : InMux
    port map (
            O => \N__53302\,
            I => \N__53275\
        );

    \I__11432\ : CascadeMux
    port map (
            O => \N__53301\,
            I => \N__53272\
        );

    \I__11431\ : InMux
    port map (
            O => \N__53300\,
            I => \N__53267\
        );

    \I__11430\ : InMux
    port map (
            O => \N__53299\,
            I => \N__53267\
        );

    \I__11429\ : InMux
    port map (
            O => \N__53298\,
            I => \N__53264\
        );

    \I__11428\ : InMux
    port map (
            O => \N__53297\,
            I => \N__53259\
        );

    \I__11427\ : InMux
    port map (
            O => \N__53296\,
            I => \N__53259\
        );

    \I__11426\ : InMux
    port map (
            O => \N__53295\,
            I => \N__53250\
        );

    \I__11425\ : InMux
    port map (
            O => \N__53294\,
            I => \N__53250\
        );

    \I__11424\ : InMux
    port map (
            O => \N__53293\,
            I => \N__53250\
        );

    \I__11423\ : InMux
    port map (
            O => \N__53292\,
            I => \N__53250\
        );

    \I__11422\ : CascadeMux
    port map (
            O => \N__53291\,
            I => \N__53246\
        );

    \I__11421\ : InMux
    port map (
            O => \N__53290\,
            I => \N__53242\
        );

    \I__11420\ : InMux
    port map (
            O => \N__53289\,
            I => \N__53239\
        );

    \I__11419\ : CascadeMux
    port map (
            O => \N__53288\,
            I => \N__53234\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__53285\,
            I => \N__53226\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__53282\,
            I => \N__53226\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__53275\,
            I => \N__53223\
        );

    \I__11415\ : InMux
    port map (
            O => \N__53272\,
            I => \N__53220\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__53267\,
            I => \N__53217\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__53264\,
            I => \N__53209\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__53259\,
            I => \N__53209\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__53250\,
            I => \N__53209\
        );

    \I__11410\ : CascadeMux
    port map (
            O => \N__53249\,
            I => \N__53206\
        );

    \I__11409\ : InMux
    port map (
            O => \N__53246\,
            I => \N__53201\
        );

    \I__11408\ : InMux
    port map (
            O => \N__53245\,
            I => \N__53198\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__53242\,
            I => \N__53195\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__53239\,
            I => \N__53192\
        );

    \I__11405\ : InMux
    port map (
            O => \N__53238\,
            I => \N__53187\
        );

    \I__11404\ : InMux
    port map (
            O => \N__53237\,
            I => \N__53187\
        );

    \I__11403\ : InMux
    port map (
            O => \N__53234\,
            I => \N__53184\
        );

    \I__11402\ : InMux
    port map (
            O => \N__53233\,
            I => \N__53181\
        );

    \I__11401\ : InMux
    port map (
            O => \N__53232\,
            I => \N__53178\
        );

    \I__11400\ : InMux
    port map (
            O => \N__53231\,
            I => \N__53174\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__53226\,
            I => \N__53171\
        );

    \I__11398\ : Span4Mux_v
    port map (
            O => \N__53223\,
            I => \N__53166\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__53220\,
            I => \N__53166\
        );

    \I__11396\ : Span4Mux_v
    port map (
            O => \N__53217\,
            I => \N__53162\
        );

    \I__11395\ : InMux
    port map (
            O => \N__53216\,
            I => \N__53158\
        );

    \I__11394\ : Span4Mux_v
    port map (
            O => \N__53209\,
            I => \N__53155\
        );

    \I__11393\ : InMux
    port map (
            O => \N__53206\,
            I => \N__53152\
        );

    \I__11392\ : InMux
    port map (
            O => \N__53205\,
            I => \N__53147\
        );

    \I__11391\ : InMux
    port map (
            O => \N__53204\,
            I => \N__53147\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__53201\,
            I => \N__53141\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__53198\,
            I => \N__53138\
        );

    \I__11388\ : Span4Mux_h
    port map (
            O => \N__53195\,
            I => \N__53133\
        );

    \I__11387\ : Span4Mux_h
    port map (
            O => \N__53192\,
            I => \N__53133\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__53187\,
            I => \N__53130\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__53184\,
            I => \N__53127\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__53181\,
            I => \N__53122\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__53178\,
            I => \N__53122\
        );

    \I__11382\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53119\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__53174\,
            I => \N__53112\
        );

    \I__11380\ : Span4Mux_h
    port map (
            O => \N__53171\,
            I => \N__53112\
        );

    \I__11379\ : Span4Mux_v
    port map (
            O => \N__53166\,
            I => \N__53112\
        );

    \I__11378\ : InMux
    port map (
            O => \N__53165\,
            I => \N__53109\
        );

    \I__11377\ : Span4Mux_h
    port map (
            O => \N__53162\,
            I => \N__53106\
        );

    \I__11376\ : InMux
    port map (
            O => \N__53161\,
            I => \N__53103\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__53158\,
            I => \N__53094\
        );

    \I__11374\ : Span4Mux_h
    port map (
            O => \N__53155\,
            I => \N__53094\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__53152\,
            I => \N__53094\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__53147\,
            I => \N__53094\
        );

    \I__11371\ : InMux
    port map (
            O => \N__53146\,
            I => \N__53089\
        );

    \I__11370\ : InMux
    port map (
            O => \N__53145\,
            I => \N__53089\
        );

    \I__11369\ : InMux
    port map (
            O => \N__53144\,
            I => \N__53086\
        );

    \I__11368\ : Span4Mux_h
    port map (
            O => \N__53141\,
            I => \N__53079\
        );

    \I__11367\ : Span4Mux_h
    port map (
            O => \N__53138\,
            I => \N__53079\
        );

    \I__11366\ : Span4Mux_v
    port map (
            O => \N__53133\,
            I => \N__53079\
        );

    \I__11365\ : Span4Mux_h
    port map (
            O => \N__53130\,
            I => \N__53072\
        );

    \I__11364\ : Span4Mux_v
    port map (
            O => \N__53127\,
            I => \N__53072\
        );

    \I__11363\ : Span4Mux_h
    port map (
            O => \N__53122\,
            I => \N__53072\
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__53119\,
            I => \N__53067\
        );

    \I__11361\ : Sp12to4
    port map (
            O => \N__53112\,
            I => \N__53067\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__53109\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11359\ : Odrv4
    port map (
            O => \N__53106\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__53103\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11357\ : Odrv4
    port map (
            O => \N__53094\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__53089\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__53086\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11354\ : Odrv4
    port map (
            O => \N__53079\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11353\ : Odrv4
    port map (
            O => \N__53072\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11352\ : Odrv12
    port map (
            O => \N__53067\,
            I => \ALU.combOperand2_a0_0Z0Z_6\
        );

    \I__11351\ : InMux
    port map (
            O => \N__53048\,
            I => \N__53045\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__53045\,
            I => \N__53042\
        );

    \I__11349\ : Span4Mux_v
    port map (
            O => \N__53042\,
            I => \N__53039\
        );

    \I__11348\ : Odrv4
    port map (
            O => \N__53039\,
            I => \ALU.status_RNO_22Z0Z_0\
        );

    \I__11347\ : InMux
    port map (
            O => \N__53036\,
            I => \N__53033\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__53033\,
            I => \ALU.status_14_6_0\
        );

    \I__11345\ : InMux
    port map (
            O => \N__53030\,
            I => \N__53027\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__53027\,
            I => \N__53024\
        );

    \I__11343\ : Sp12to4
    port map (
            O => \N__53024\,
            I => \N__53021\
        );

    \I__11342\ : Span12Mux_v
    port map (
            O => \N__53021\,
            I => \N__53018\
        );

    \I__11341\ : Span12Mux_h
    port map (
            O => \N__53018\,
            I => \N__53015\
        );

    \I__11340\ : Odrv12
    port map (
            O => \N__53015\,
            I => \ALU.status_17_I_21_c_RNOZ0\
        );

    \I__11339\ : InMux
    port map (
            O => \N__53012\,
            I => \N__53003\
        );

    \I__11338\ : InMux
    port map (
            O => \N__53011\,
            I => \N__53000\
        );

    \I__11337\ : InMux
    port map (
            O => \N__53010\,
            I => \N__52997\
        );

    \I__11336\ : InMux
    port map (
            O => \N__53009\,
            I => \N__52994\
        );

    \I__11335\ : InMux
    port map (
            O => \N__53008\,
            I => \N__52991\
        );

    \I__11334\ : InMux
    port map (
            O => \N__53007\,
            I => \N__52988\
        );

    \I__11333\ : InMux
    port map (
            O => \N__53006\,
            I => \N__52984\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__53003\,
            I => \N__52981\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__53000\,
            I => \N__52974\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__52997\,
            I => \N__52974\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__52994\,
            I => \N__52974\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__52991\,
            I => \N__52971\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__52988\,
            I => \N__52968\
        );

    \I__11326\ : InMux
    port map (
            O => \N__52987\,
            I => \N__52965\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__52984\,
            I => \N__52958\
        );

    \I__11324\ : Span4Mux_h
    port map (
            O => \N__52981\,
            I => \N__52958\
        );

    \I__11323\ : Span4Mux_v
    port map (
            O => \N__52974\,
            I => \N__52958\
        );

    \I__11322\ : Span4Mux_h
    port map (
            O => \N__52971\,
            I => \N__52953\
        );

    \I__11321\ : Span4Mux_h
    port map (
            O => \N__52968\,
            I => \N__52953\
        );

    \I__11320\ : LocalMux
    port map (
            O => \N__52965\,
            I => \N__52950\
        );

    \I__11319\ : Span4Mux_h
    port map (
            O => \N__52958\,
            I => \N__52947\
        );

    \I__11318\ : Span4Mux_h
    port map (
            O => \N__52953\,
            I => \N__52942\
        );

    \I__11317\ : Span4Mux_h
    port map (
            O => \N__52950\,
            I => \N__52942\
        );

    \I__11316\ : Odrv4
    port map (
            O => \N__52947\,
            I => \ALU.mult_15\
        );

    \I__11315\ : Odrv4
    port map (
            O => \N__52942\,
            I => \ALU.mult_15\
        );

    \I__11314\ : InMux
    port map (
            O => \N__52937\,
            I => \N__52928\
        );

    \I__11313\ : InMux
    port map (
            O => \N__52936\,
            I => \N__52925\
        );

    \I__11312\ : InMux
    port map (
            O => \N__52935\,
            I => \N__52922\
        );

    \I__11311\ : InMux
    port map (
            O => \N__52934\,
            I => \N__52919\
        );

    \I__11310\ : InMux
    port map (
            O => \N__52933\,
            I => \N__52916\
        );

    \I__11309\ : InMux
    port map (
            O => \N__52932\,
            I => \N__52913\
        );

    \I__11308\ : InMux
    port map (
            O => \N__52931\,
            I => \N__52910\
        );

    \I__11307\ : LocalMux
    port map (
            O => \N__52928\,
            I => \N__52905\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__52925\,
            I => \N__52905\
        );

    \I__11305\ : LocalMux
    port map (
            O => \N__52922\,
            I => \N__52902\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__52919\,
            I => \ALU.a_15_1_15\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__52916\,
            I => \ALU.a_15_1_15\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__52913\,
            I => \ALU.a_15_1_15\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__52910\,
            I => \ALU.a_15_1_15\
        );

    \I__11300\ : Odrv4
    port map (
            O => \N__52905\,
            I => \ALU.a_15_1_15\
        );

    \I__11299\ : Odrv4
    port map (
            O => \N__52902\,
            I => \ALU.a_15_1_15\
        );

    \I__11298\ : CascadeMux
    port map (
            O => \N__52889\,
            I => \N__52886\
        );

    \I__11297\ : InMux
    port map (
            O => \N__52886\,
            I => \N__52883\
        );

    \I__11296\ : LocalMux
    port map (
            O => \N__52883\,
            I => \N__52880\
        );

    \I__11295\ : Span4Mux_v
    port map (
            O => \N__52880\,
            I => \N__52875\
        );

    \I__11294\ : InMux
    port map (
            O => \N__52879\,
            I => \N__52872\
        );

    \I__11293\ : InMux
    port map (
            O => \N__52878\,
            I => \N__52867\
        );

    \I__11292\ : Span4Mux_h
    port map (
            O => \N__52875\,
            I => \N__52863\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__52872\,
            I => \N__52860\
        );

    \I__11290\ : InMux
    port map (
            O => \N__52871\,
            I => \N__52857\
        );

    \I__11289\ : InMux
    port map (
            O => \N__52870\,
            I => \N__52853\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__52867\,
            I => \N__52850\
        );

    \I__11287\ : InMux
    port map (
            O => \N__52866\,
            I => \N__52847\
        );

    \I__11286\ : Span4Mux_v
    port map (
            O => \N__52863\,
            I => \N__52844\
        );

    \I__11285\ : Span4Mux_v
    port map (
            O => \N__52860\,
            I => \N__52839\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__52857\,
            I => \N__52839\
        );

    \I__11283\ : InMux
    port map (
            O => \N__52856\,
            I => \N__52836\
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__52853\,
            I => \N__52833\
        );

    \I__11281\ : Span4Mux_v
    port map (
            O => \N__52850\,
            I => \N__52830\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__52847\,
            I => \N__52825\
        );

    \I__11279\ : Span4Mux_h
    port map (
            O => \N__52844\,
            I => \N__52825\
        );

    \I__11278\ : Span4Mux_h
    port map (
            O => \N__52839\,
            I => \N__52822\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__52836\,
            I => \N__52813\
        );

    \I__11276\ : Span4Mux_v
    port map (
            O => \N__52833\,
            I => \N__52813\
        );

    \I__11275\ : Span4Mux_v
    port map (
            O => \N__52830\,
            I => \N__52813\
        );

    \I__11274\ : Span4Mux_v
    port map (
            O => \N__52825\,
            I => \N__52813\
        );

    \I__11273\ : Odrv4
    port map (
            O => \N__52822\,
            I => \ALU.a_15_m1_9\
        );

    \I__11272\ : Odrv4
    port map (
            O => \N__52813\,
            I => \ALU.a_15_m1_9\
        );

    \I__11271\ : InMux
    port map (
            O => \N__52808\,
            I => \N__52802\
        );

    \I__11270\ : CascadeMux
    port map (
            O => \N__52807\,
            I => \N__52798\
        );

    \I__11269\ : InMux
    port map (
            O => \N__52806\,
            I => \N__52795\
        );

    \I__11268\ : InMux
    port map (
            O => \N__52805\,
            I => \N__52792\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__52802\,
            I => \N__52789\
        );

    \I__11266\ : InMux
    port map (
            O => \N__52801\,
            I => \N__52783\
        );

    \I__11265\ : InMux
    port map (
            O => \N__52798\,
            I => \N__52780\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__52795\,
            I => \N__52777\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__52792\,
            I => \N__52772\
        );

    \I__11262\ : Span4Mux_v
    port map (
            O => \N__52789\,
            I => \N__52772\
        );

    \I__11261\ : InMux
    port map (
            O => \N__52788\,
            I => \N__52769\
        );

    \I__11260\ : InMux
    port map (
            O => \N__52787\,
            I => \N__52766\
        );

    \I__11259\ : InMux
    port map (
            O => \N__52786\,
            I => \N__52763\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__52783\,
            I => \N__52754\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__52780\,
            I => \N__52754\
        );

    \I__11256\ : Span4Mux_v
    port map (
            O => \N__52777\,
            I => \N__52754\
        );

    \I__11255\ : Span4Mux_h
    port map (
            O => \N__52772\,
            I => \N__52754\
        );

    \I__11254\ : LocalMux
    port map (
            O => \N__52769\,
            I => \ALU.mult_546_c_RNIJOT4JZ0Z8\
        );

    \I__11253\ : LocalMux
    port map (
            O => \N__52766\,
            I => \ALU.mult_546_c_RNIJOT4JZ0Z8\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__52763\,
            I => \ALU.mult_546_c_RNIJOT4JZ0Z8\
        );

    \I__11251\ : Odrv4
    port map (
            O => \N__52754\,
            I => \ALU.mult_546_c_RNIJOT4JZ0Z8\
        );

    \I__11250\ : InMux
    port map (
            O => \N__52745\,
            I => \N__52741\
        );

    \I__11249\ : InMux
    port map (
            O => \N__52744\,
            I => \N__52738\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__52741\,
            I => \N__52735\
        );

    \I__11247\ : LocalMux
    port map (
            O => \N__52738\,
            I => \N__52732\
        );

    \I__11246\ : Span4Mux_v
    port map (
            O => \N__52735\,
            I => \N__52729\
        );

    \I__11245\ : Span4Mux_v
    port map (
            O => \N__52732\,
            I => \N__52726\
        );

    \I__11244\ : Span4Mux_h
    port map (
            O => \N__52729\,
            I => \N__52723\
        );

    \I__11243\ : Span4Mux_h
    port map (
            O => \N__52726\,
            I => \N__52720\
        );

    \I__11242\ : Span4Mux_h
    port map (
            O => \N__52723\,
            I => \N__52717\
        );

    \I__11241\ : Span4Mux_v
    port map (
            O => \N__52720\,
            I => \N__52714\
        );

    \I__11240\ : Odrv4
    port map (
            O => \N__52717\,
            I => \ALU.dZ0Z_9\
        );

    \I__11239\ : Odrv4
    port map (
            O => \N__52714\,
            I => \ALU.dZ0Z_9\
        );

    \I__11238\ : InMux
    port map (
            O => \N__52709\,
            I => \N__52706\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__52706\,
            I => \N__52702\
        );

    \I__11236\ : InMux
    port map (
            O => \N__52705\,
            I => \N__52699\
        );

    \I__11235\ : Span4Mux_v
    port map (
            O => \N__52702\,
            I => \N__52696\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__52699\,
            I => \ALU.N_835\
        );

    \I__11233\ : Odrv4
    port map (
            O => \N__52696\,
            I => \ALU.N_835\
        );

    \I__11232\ : CascadeMux
    port map (
            O => \N__52691\,
            I => \ALU.d_RNIPFFDD1_0Z0Z_6_cascade_\
        );

    \I__11231\ : CascadeMux
    port map (
            O => \N__52688\,
            I => \ALU.N_863_cascade_\
        );

    \I__11230\ : InMux
    port map (
            O => \N__52685\,
            I => \N__52680\
        );

    \I__11229\ : InMux
    port map (
            O => \N__52684\,
            I => \N__52675\
        );

    \I__11228\ : InMux
    port map (
            O => \N__52683\,
            I => \N__52672\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__52680\,
            I => \N__52669\
        );

    \I__11226\ : InMux
    port map (
            O => \N__52679\,
            I => \N__52666\
        );

    \I__11225\ : InMux
    port map (
            O => \N__52678\,
            I => \N__52663\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__52675\,
            I => \N__52660\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__52672\,
            I => \N__52657\
        );

    \I__11222\ : Span12Mux_h
    port map (
            O => \N__52669\,
            I => \N__52654\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__52666\,
            I => \N__52645\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__52663\,
            I => \N__52645\
        );

    \I__11219\ : Span12Mux_v
    port map (
            O => \N__52660\,
            I => \N__52645\
        );

    \I__11218\ : Span12Mux_h
    port map (
            O => \N__52657\,
            I => \N__52645\
        );

    \I__11217\ : Odrv12
    port map (
            O => \N__52654\,
            I => \ALU.d_RNIN3H0DZ0Z_3\
        );

    \I__11216\ : Odrv12
    port map (
            O => \N__52645\,
            I => \ALU.d_RNIN3H0DZ0Z_3\
        );

    \I__11215\ : CascadeMux
    port map (
            O => \N__52640\,
            I => \ALU.d_RNIGPBNB6Z0Z_2_cascade_\
        );

    \I__11214\ : InMux
    port map (
            O => \N__52637\,
            I => \N__52632\
        );

    \I__11213\ : CascadeMux
    port map (
            O => \N__52636\,
            I => \N__52629\
        );

    \I__11212\ : InMux
    port map (
            O => \N__52635\,
            I => \N__52624\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__52632\,
            I => \N__52620\
        );

    \I__11210\ : InMux
    port map (
            O => \N__52629\,
            I => \N__52616\
        );

    \I__11209\ : InMux
    port map (
            O => \N__52628\,
            I => \N__52613\
        );

    \I__11208\ : InMux
    port map (
            O => \N__52627\,
            I => \N__52609\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__52624\,
            I => \N__52606\
        );

    \I__11206\ : InMux
    port map (
            O => \N__52623\,
            I => \N__52603\
        );

    \I__11205\ : Span4Mux_h
    port map (
            O => \N__52620\,
            I => \N__52600\
        );

    \I__11204\ : InMux
    port map (
            O => \N__52619\,
            I => \N__52597\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__52616\,
            I => \N__52592\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__52613\,
            I => \N__52592\
        );

    \I__11201\ : InMux
    port map (
            O => \N__52612\,
            I => \N__52589\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__52609\,
            I => \N__52586\
        );

    \I__11199\ : Span4Mux_h
    port map (
            O => \N__52606\,
            I => \N__52583\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__52603\,
            I => \N__52580\
        );

    \I__11197\ : Span4Mux_h
    port map (
            O => \N__52600\,
            I => \N__52577\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__52597\,
            I => \N__52572\
        );

    \I__11195\ : Span4Mux_v
    port map (
            O => \N__52592\,
            I => \N__52572\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__52589\,
            I => \N__52565\
        );

    \I__11193\ : Span4Mux_h
    port map (
            O => \N__52586\,
            I => \N__52565\
        );

    \I__11192\ : Span4Mux_v
    port map (
            O => \N__52583\,
            I => \N__52565\
        );

    \I__11191\ : Span4Mux_h
    port map (
            O => \N__52580\,
            I => \N__52562\
        );

    \I__11190\ : Span4Mux_h
    port map (
            O => \N__52577\,
            I => \N__52559\
        );

    \I__11189\ : Span4Mux_h
    port map (
            O => \N__52572\,
            I => \N__52556\
        );

    \I__11188\ : Sp12to4
    port map (
            O => \N__52565\,
            I => \N__52553\
        );

    \I__11187\ : Span4Mux_h
    port map (
            O => \N__52562\,
            I => \N__52548\
        );

    \I__11186\ : Span4Mux_v
    port map (
            O => \N__52559\,
            I => \N__52548\
        );

    \I__11185\ : Odrv4
    port map (
            O => \N__52556\,
            I => \ALU.a_15_m0_5\
        );

    \I__11184\ : Odrv12
    port map (
            O => \N__52553\,
            I => \ALU.a_15_m0_5\
        );

    \I__11183\ : Odrv4
    port map (
            O => \N__52548\,
            I => \ALU.a_15_m0_5\
        );

    \I__11182\ : IoInMux
    port map (
            O => \N__52541\,
            I => \N__52538\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__52538\,
            I => \N__52535\
        );

    \I__11180\ : IoSpan4Mux
    port map (
            O => \N__52535\,
            I => \N__52532\
        );

    \I__11179\ : IoSpan4Mux
    port map (
            O => \N__52532\,
            I => \N__52528\
        );

    \I__11178\ : IoInMux
    port map (
            O => \N__52531\,
            I => \N__52524\
        );

    \I__11177\ : Span4Mux_s2_h
    port map (
            O => \N__52528\,
            I => \N__52521\
        );

    \I__11176\ : InMux
    port map (
            O => \N__52527\,
            I => \N__52518\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__52524\,
            I => \N__52515\
        );

    \I__11174\ : Sp12to4
    port map (
            O => \N__52521\,
            I => \N__52510\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__52518\,
            I => \N__52510\
        );

    \I__11172\ : Span12Mux_s8_h
    port map (
            O => \N__52515\,
            I => \N__52507\
        );

    \I__11171\ : Span12Mux_h
    port map (
            O => \N__52510\,
            I => \N__52504\
        );

    \I__11170\ : Odrv12
    port map (
            O => \N__52507\,
            I => bus_5
        );

    \I__11169\ : Odrv12
    port map (
            O => \N__52504\,
            I => bus_5
        );

    \I__11168\ : InMux
    port map (
            O => \N__52499\,
            I => \N__52496\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__52496\,
            I => \ALU.c_RNINGV0T2Z0Z_15\
        );

    \I__11166\ : InMux
    port map (
            O => \N__52493\,
            I => \N__52490\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__52490\,
            I => \ALU.d_RNIPFFDD1Z0Z_6\
        );

    \I__11164\ : CascadeMux
    port map (
            O => \N__52487\,
            I => \N__52484\
        );

    \I__11163\ : InMux
    port map (
            O => \N__52484\,
            I => \N__52481\
        );

    \I__11162\ : LocalMux
    port map (
            O => \N__52481\,
            I => \N__52478\
        );

    \I__11161\ : Span4Mux_h
    port map (
            O => \N__52478\,
            I => \N__52474\
        );

    \I__11160\ : InMux
    port map (
            O => \N__52477\,
            I => \N__52471\
        );

    \I__11159\ : Span4Mux_h
    port map (
            O => \N__52474\,
            I => \N__52468\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__52471\,
            I => \N__52465\
        );

    \I__11157\ : Span4Mux_v
    port map (
            O => \N__52468\,
            I => \N__52462\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__52465\,
            I => \N__52459\
        );

    \I__11155\ : Span4Mux_v
    port map (
            O => \N__52462\,
            I => \N__52456\
        );

    \I__11154\ : Odrv4
    port map (
            O => \N__52459\,
            I => \ALU.eZ0Z_13\
        );

    \I__11153\ : Odrv4
    port map (
            O => \N__52456\,
            I => \ALU.eZ0Z_13\
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__52451\,
            I => \N__52448\
        );

    \I__11151\ : InMux
    port map (
            O => \N__52448\,
            I => \N__52444\
        );

    \I__11150\ : InMux
    port map (
            O => \N__52447\,
            I => \N__52441\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__52444\,
            I => \N__52438\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__52441\,
            I => \N__52435\
        );

    \I__11147\ : Span4Mux_h
    port map (
            O => \N__52438\,
            I => \N__52432\
        );

    \I__11146\ : Span4Mux_h
    port map (
            O => \N__52435\,
            I => \N__52429\
        );

    \I__11145\ : Span4Mux_h
    port map (
            O => \N__52432\,
            I => \N__52426\
        );

    \I__11144\ : Span4Mux_h
    port map (
            O => \N__52429\,
            I => \N__52423\
        );

    \I__11143\ : Sp12to4
    port map (
            O => \N__52426\,
            I => \N__52420\
        );

    \I__11142\ : Span4Mux_v
    port map (
            O => \N__52423\,
            I => \N__52417\
        );

    \I__11141\ : Odrv12
    port map (
            O => \N__52420\,
            I => \ALU.eZ0Z_14\
        );

    \I__11140\ : Odrv4
    port map (
            O => \N__52417\,
            I => \ALU.eZ0Z_14\
        );

    \I__11139\ : InMux
    port map (
            O => \N__52412\,
            I => \N__52407\
        );

    \I__11138\ : InMux
    port map (
            O => \N__52411\,
            I => \N__52404\
        );

    \I__11137\ : InMux
    port map (
            O => \N__52410\,
            I => \N__52401\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__52407\,
            I => \N__52398\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__52404\,
            I => \N__52395\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__52401\,
            I => \N__52392\
        );

    \I__11133\ : Span4Mux_h
    port map (
            O => \N__52398\,
            I => \N__52389\
        );

    \I__11132\ : Span4Mux_v
    port map (
            O => \N__52395\,
            I => \N__52386\
        );

    \I__11131\ : Span4Mux_v
    port map (
            O => \N__52392\,
            I => \N__52383\
        );

    \I__11130\ : Span4Mux_h
    port map (
            O => \N__52389\,
            I => \N__52380\
        );

    \I__11129\ : Span4Mux_h
    port map (
            O => \N__52386\,
            I => \N__52375\
        );

    \I__11128\ : Span4Mux_v
    port map (
            O => \N__52383\,
            I => \N__52375\
        );

    \I__11127\ : Span4Mux_h
    port map (
            O => \N__52380\,
            I => \N__52372\
        );

    \I__11126\ : Span4Mux_h
    port map (
            O => \N__52375\,
            I => \N__52369\
        );

    \I__11125\ : Span4Mux_v
    port map (
            O => \N__52372\,
            I => \N__52366\
        );

    \I__11124\ : Span4Mux_h
    port map (
            O => \N__52369\,
            I => \N__52363\
        );

    \I__11123\ : Odrv4
    port map (
            O => \N__52366\,
            I => g_12
        );

    \I__11122\ : Odrv4
    port map (
            O => \N__52363\,
            I => g_12
        );

    \I__11121\ : InMux
    port map (
            O => \N__52358\,
            I => \N__52354\
        );

    \I__11120\ : CascadeMux
    port map (
            O => \N__52357\,
            I => \N__52351\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__52354\,
            I => \N__52347\
        );

    \I__11118\ : InMux
    port map (
            O => \N__52351\,
            I => \N__52344\
        );

    \I__11117\ : InMux
    port map (
            O => \N__52350\,
            I => \N__52341\
        );

    \I__11116\ : Span4Mux_v
    port map (
            O => \N__52347\,
            I => \N__52338\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__52344\,
            I => \N__52335\
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__52341\,
            I => \N__52332\
        );

    \I__11113\ : Span4Mux_h
    port map (
            O => \N__52338\,
            I => \N__52329\
        );

    \I__11112\ : Sp12to4
    port map (
            O => \N__52335\,
            I => \N__52326\
        );

    \I__11111\ : Span4Mux_v
    port map (
            O => \N__52332\,
            I => \N__52323\
        );

    \I__11110\ : Span4Mux_h
    port map (
            O => \N__52329\,
            I => \N__52320\
        );

    \I__11109\ : Span12Mux_v
    port map (
            O => \N__52326\,
            I => \N__52315\
        );

    \I__11108\ : Sp12to4
    port map (
            O => \N__52323\,
            I => \N__52315\
        );

    \I__11107\ : Sp12to4
    port map (
            O => \N__52320\,
            I => \N__52312\
        );

    \I__11106\ : Span12Mux_h
    port map (
            O => \N__52315\,
            I => \N__52307\
        );

    \I__11105\ : Span12Mux_s10_h
    port map (
            O => \N__52312\,
            I => \N__52307\
        );

    \I__11104\ : Odrv12
    port map (
            O => \N__52307\,
            I => g_13
        );

    \I__11103\ : InMux
    port map (
            O => \N__52304\,
            I => \N__52301\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__52301\,
            I => \N__52298\
        );

    \I__11101\ : Span4Mux_v
    port map (
            O => \N__52298\,
            I => \N__52295\
        );

    \I__11100\ : Span4Mux_h
    port map (
            O => \N__52295\,
            I => \N__52292\
        );

    \I__11099\ : Span4Mux_h
    port map (
            O => \N__52292\,
            I => \N__52288\
        );

    \I__11098\ : InMux
    port map (
            O => \N__52291\,
            I => \N__52285\
        );

    \I__11097\ : Span4Mux_h
    port map (
            O => \N__52288\,
            I => \N__52281\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__52285\,
            I => \N__52278\
        );

    \I__11095\ : InMux
    port map (
            O => \N__52284\,
            I => \N__52275\
        );

    \I__11094\ : Span4Mux_v
    port map (
            O => \N__52281\,
            I => \N__52270\
        );

    \I__11093\ : Span4Mux_h
    port map (
            O => \N__52278\,
            I => \N__52270\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__52275\,
            I => \N__52267\
        );

    \I__11091\ : Span4Mux_h
    port map (
            O => \N__52270\,
            I => \N__52264\
        );

    \I__11090\ : Span4Mux_h
    port map (
            O => \N__52267\,
            I => \N__52261\
        );

    \I__11089\ : Span4Mux_h
    port map (
            O => \N__52264\,
            I => \N__52258\
        );

    \I__11088\ : Span4Mux_v
    port map (
            O => \N__52261\,
            I => \N__52255\
        );

    \I__11087\ : Span4Mux_v
    port map (
            O => \N__52258\,
            I => \N__52252\
        );

    \I__11086\ : Odrv4
    port map (
            O => \N__52255\,
            I => g_14
        );

    \I__11085\ : Odrv4
    port map (
            O => \N__52252\,
            I => g_14
        );

    \I__11084\ : CascadeMux
    port map (
            O => \N__52247\,
            I => \N__52242\
        );

    \I__11083\ : CascadeMux
    port map (
            O => \N__52246\,
            I => \N__52237\
        );

    \I__11082\ : CascadeMux
    port map (
            O => \N__52245\,
            I => \N__52233\
        );

    \I__11081\ : InMux
    port map (
            O => \N__52242\,
            I => \N__52230\
        );

    \I__11080\ : InMux
    port map (
            O => \N__52241\,
            I => \N__52227\
        );

    \I__11079\ : InMux
    port map (
            O => \N__52240\,
            I => \N__52224\
        );

    \I__11078\ : InMux
    port map (
            O => \N__52237\,
            I => \N__52220\
        );

    \I__11077\ : InMux
    port map (
            O => \N__52236\,
            I => \N__52217\
        );

    \I__11076\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52214\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__52230\,
            I => \N__52211\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__52227\,
            I => \N__52206\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__52224\,
            I => \N__52206\
        );

    \I__11072\ : InMux
    port map (
            O => \N__52223\,
            I => \N__52202\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__52220\,
            I => \N__52199\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__52217\,
            I => \N__52196\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__52214\,
            I => \N__52189\
        );

    \I__11068\ : Span4Mux_h
    port map (
            O => \N__52211\,
            I => \N__52189\
        );

    \I__11067\ : Span4Mux_v
    port map (
            O => \N__52206\,
            I => \N__52189\
        );

    \I__11066\ : InMux
    port map (
            O => \N__52205\,
            I => \N__52186\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__52202\,
            I => \N__52183\
        );

    \I__11064\ : Span4Mux_h
    port map (
            O => \N__52199\,
            I => \N__52178\
        );

    \I__11063\ : Span4Mux_v
    port map (
            O => \N__52196\,
            I => \N__52178\
        );

    \I__11062\ : Span4Mux_h
    port map (
            O => \N__52189\,
            I => \N__52175\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__52186\,
            I => \ALU.a_15_ns_1_1\
        );

    \I__11060\ : Odrv4
    port map (
            O => \N__52183\,
            I => \ALU.a_15_ns_1_1\
        );

    \I__11059\ : Odrv4
    port map (
            O => \N__52178\,
            I => \ALU.a_15_ns_1_1\
        );

    \I__11058\ : Odrv4
    port map (
            O => \N__52175\,
            I => \ALU.a_15_ns_1_1\
        );

    \I__11057\ : InMux
    port map (
            O => \N__52166\,
            I => \N__52162\
        );

    \I__11056\ : InMux
    port map (
            O => \N__52165\,
            I => \N__52159\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__52162\,
            I => \N__52156\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__52159\,
            I => \N__52153\
        );

    \I__11053\ : Span4Mux_v
    port map (
            O => \N__52156\,
            I => \N__52150\
        );

    \I__11052\ : Span4Mux_v
    port map (
            O => \N__52153\,
            I => \N__52147\
        );

    \I__11051\ : Span4Mux_h
    port map (
            O => \N__52150\,
            I => \N__52144\
        );

    \I__11050\ : Span4Mux_h
    port map (
            O => \N__52147\,
            I => \N__52141\
        );

    \I__11049\ : Span4Mux_h
    port map (
            O => \N__52144\,
            I => \N__52138\
        );

    \I__11048\ : Span4Mux_h
    port map (
            O => \N__52141\,
            I => \N__52135\
        );

    \I__11047\ : Span4Mux_v
    port map (
            O => \N__52138\,
            I => \N__52132\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__52135\,
            I => \N__52129\
        );

    \I__11045\ : Odrv4
    port map (
            O => \N__52132\,
            I => \ALU.dZ0Z_1\
        );

    \I__11044\ : Odrv4
    port map (
            O => \N__52129\,
            I => \ALU.dZ0Z_1\
        );

    \I__11043\ : InMux
    port map (
            O => \N__52124\,
            I => \N__52119\
        );

    \I__11042\ : InMux
    port map (
            O => \N__52123\,
            I => \N__52114\
        );

    \I__11041\ : InMux
    port map (
            O => \N__52122\,
            I => \N__52111\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__52119\,
            I => \N__52108\
        );

    \I__11039\ : InMux
    port map (
            O => \N__52118\,
            I => \N__52105\
        );

    \I__11038\ : InMux
    port map (
            O => \N__52117\,
            I => \N__52102\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__52114\,
            I => \N__52097\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__52111\,
            I => \N__52097\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__52108\,
            I => \N__52093\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__52105\,
            I => \N__52090\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__52102\,
            I => \N__52087\
        );

    \I__11032\ : Span4Mux_v
    port map (
            O => \N__52097\,
            I => \N__52084\
        );

    \I__11031\ : InMux
    port map (
            O => \N__52096\,
            I => \N__52081\
        );

    \I__11030\ : Span4Mux_h
    port map (
            O => \N__52093\,
            I => \N__52077\
        );

    \I__11029\ : Span4Mux_v
    port map (
            O => \N__52090\,
            I => \N__52072\
        );

    \I__11028\ : Span4Mux_v
    port map (
            O => \N__52087\,
            I => \N__52072\
        );

    \I__11027\ : Sp12to4
    port map (
            O => \N__52084\,
            I => \N__52067\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__52081\,
            I => \N__52067\
        );

    \I__11025\ : InMux
    port map (
            O => \N__52080\,
            I => \N__52064\
        );

    \I__11024\ : Odrv4
    port map (
            O => \N__52077\,
            I => \ALU.d_RNINUGCF4Z0Z_0\
        );

    \I__11023\ : Odrv4
    port map (
            O => \N__52072\,
            I => \ALU.d_RNINUGCF4Z0Z_0\
        );

    \I__11022\ : Odrv12
    port map (
            O => \N__52067\,
            I => \ALU.d_RNINUGCF4Z0Z_0\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__52064\,
            I => \ALU.d_RNINUGCF4Z0Z_0\
        );

    \I__11020\ : InMux
    port map (
            O => \N__52055\,
            I => \N__52046\
        );

    \I__11019\ : InMux
    port map (
            O => \N__52054\,
            I => \N__52043\
        );

    \I__11018\ : InMux
    port map (
            O => \N__52053\,
            I => \N__52040\
        );

    \I__11017\ : InMux
    port map (
            O => \N__52052\,
            I => \N__52037\
        );

    \I__11016\ : InMux
    port map (
            O => \N__52051\,
            I => \N__52034\
        );

    \I__11015\ : InMux
    port map (
            O => \N__52050\,
            I => \N__52030\
        );

    \I__11014\ : InMux
    port map (
            O => \N__52049\,
            I => \N__52027\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__52046\,
            I => \N__52024\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__52043\,
            I => \N__52021\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__52040\,
            I => \N__52014\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__52037\,
            I => \N__52014\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__52034\,
            I => \N__52014\
        );

    \I__11008\ : InMux
    port map (
            O => \N__52033\,
            I => \N__52011\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__52030\,
            I => \N__52008\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__52027\,
            I => \N__52005\
        );

    \I__11005\ : Span4Mux_h
    port map (
            O => \N__52024\,
            I => \N__52002\
        );

    \I__11004\ : Span4Mux_v
    port map (
            O => \N__52021\,
            I => \N__51999\
        );

    \I__11003\ : Span4Mux_v
    port map (
            O => \N__52014\,
            I => \N__51996\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__52011\,
            I => \N__51989\
        );

    \I__11001\ : Span4Mux_h
    port map (
            O => \N__52008\,
            I => \N__51989\
        );

    \I__11000\ : Span4Mux_v
    port map (
            O => \N__52005\,
            I => \N__51989\
        );

    \I__10999\ : Span4Mux_v
    port map (
            O => \N__52002\,
            I => \N__51986\
        );

    \I__10998\ : Span4Mux_v
    port map (
            O => \N__51999\,
            I => \N__51981\
        );

    \I__10997\ : Span4Mux_v
    port map (
            O => \N__51996\,
            I => \N__51981\
        );

    \I__10996\ : Span4Mux_v
    port map (
            O => \N__51989\,
            I => \N__51978\
        );

    \I__10995\ : Odrv4
    port map (
            O => \N__51986\,
            I => \ALU.rshift_0\
        );

    \I__10994\ : Odrv4
    port map (
            O => \N__51981\,
            I => \ALU.rshift_0\
        );

    \I__10993\ : Odrv4
    port map (
            O => \N__51978\,
            I => \ALU.rshift_0\
        );

    \I__10992\ : InMux
    port map (
            O => \N__51971\,
            I => \N__51968\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__51968\,
            I => \N__51964\
        );

    \I__10990\ : InMux
    port map (
            O => \N__51967\,
            I => \N__51961\
        );

    \I__10989\ : Span4Mux_v
    port map (
            O => \N__51964\,
            I => \N__51958\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__51961\,
            I => \N__51955\
        );

    \I__10987\ : Span4Mux_h
    port map (
            O => \N__51958\,
            I => \N__51952\
        );

    \I__10986\ : Span4Mux_v
    port map (
            O => \N__51955\,
            I => \N__51949\
        );

    \I__10985\ : Span4Mux_h
    port map (
            O => \N__51952\,
            I => \N__51946\
        );

    \I__10984\ : Span4Mux_h
    port map (
            O => \N__51949\,
            I => \N__51941\
        );

    \I__10983\ : Span4Mux_v
    port map (
            O => \N__51946\,
            I => \N__51941\
        );

    \I__10982\ : Odrv4
    port map (
            O => \N__51941\,
            I => \ALU.dZ0Z_0\
        );

    \I__10981\ : CascadeMux
    port map (
            O => \N__51938\,
            I => \N__51934\
        );

    \I__10980\ : InMux
    port map (
            O => \N__51937\,
            I => \N__51926\
        );

    \I__10979\ : InMux
    port map (
            O => \N__51934\,
            I => \N__51923\
        );

    \I__10978\ : CascadeMux
    port map (
            O => \N__51933\,
            I => \N__51920\
        );

    \I__10977\ : InMux
    port map (
            O => \N__51932\,
            I => \N__51917\
        );

    \I__10976\ : InMux
    port map (
            O => \N__51931\,
            I => \N__51914\
        );

    \I__10975\ : InMux
    port map (
            O => \N__51930\,
            I => \N__51911\
        );

    \I__10974\ : InMux
    port map (
            O => \N__51929\,
            I => \N__51908\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__51926\,
            I => \N__51905\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__51923\,
            I => \N__51901\
        );

    \I__10971\ : InMux
    port map (
            O => \N__51920\,
            I => \N__51898\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__51917\,
            I => \N__51893\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__51914\,
            I => \N__51893\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__51911\,
            I => \N__51886\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__51908\,
            I => \N__51886\
        );

    \I__10966\ : Span4Mux_v
    port map (
            O => \N__51905\,
            I => \N__51886\
        );

    \I__10965\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51883\
        );

    \I__10964\ : Span4Mux_h
    port map (
            O => \N__51901\,
            I => \N__51880\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__51898\,
            I => \N__51875\
        );

    \I__10962\ : Span4Mux_v
    port map (
            O => \N__51893\,
            I => \N__51875\
        );

    \I__10961\ : Span4Mux_v
    port map (
            O => \N__51886\,
            I => \N__51872\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__51883\,
            I => \ALU.a_15_m0_7\
        );

    \I__10959\ : Odrv4
    port map (
            O => \N__51880\,
            I => \ALU.a_15_m0_7\
        );

    \I__10958\ : Odrv4
    port map (
            O => \N__51875\,
            I => \ALU.a_15_m0_7\
        );

    \I__10957\ : Odrv4
    port map (
            O => \N__51872\,
            I => \ALU.a_15_m0_7\
        );

    \I__10956\ : CascadeMux
    port map (
            O => \N__51863\,
            I => \N__51859\
        );

    \I__10955\ : InMux
    port map (
            O => \N__51862\,
            I => \N__51854\
        );

    \I__10954\ : InMux
    port map (
            O => \N__51859\,
            I => \N__51848\
        );

    \I__10953\ : InMux
    port map (
            O => \N__51858\,
            I => \N__51845\
        );

    \I__10952\ : InMux
    port map (
            O => \N__51857\,
            I => \N__51842\
        );

    \I__10951\ : LocalMux
    port map (
            O => \N__51854\,
            I => \N__51839\
        );

    \I__10950\ : InMux
    port map (
            O => \N__51853\,
            I => \N__51836\
        );

    \I__10949\ : InMux
    port map (
            O => \N__51852\,
            I => \N__51833\
        );

    \I__10948\ : InMux
    port map (
            O => \N__51851\,
            I => \N__51830\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__51848\,
            I => \N__51827\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__51845\,
            I => \N__51824\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__51842\,
            I => \N__51819\
        );

    \I__10944\ : Span4Mux_v
    port map (
            O => \N__51839\,
            I => \N__51819\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__51836\,
            I => \ALU.mult_492_c_RNIGN2JECZ0\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__51833\,
            I => \ALU.mult_492_c_RNIGN2JECZ0\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__51830\,
            I => \ALU.mult_492_c_RNIGN2JECZ0\
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__51827\,
            I => \ALU.mult_492_c_RNIGN2JECZ0\
        );

    \I__10939\ : Odrv4
    port map (
            O => \N__51824\,
            I => \ALU.mult_492_c_RNIGN2JECZ0\
        );

    \I__10938\ : Odrv4
    port map (
            O => \N__51819\,
            I => \ALU.mult_492_c_RNIGN2JECZ0\
        );

    \I__10937\ : InMux
    port map (
            O => \N__51806\,
            I => \N__51802\
        );

    \I__10936\ : InMux
    port map (
            O => \N__51805\,
            I => \N__51799\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__51802\,
            I => \N__51794\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__51799\,
            I => \N__51794\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__51794\,
            I => \N__51791\
        );

    \I__10932\ : Odrv4
    port map (
            O => \N__51791\,
            I => \ALU.dZ0Z_7\
        );

    \I__10931\ : CascadeMux
    port map (
            O => \N__51788\,
            I => \N__51785\
        );

    \I__10930\ : InMux
    port map (
            O => \N__51785\,
            I => \N__51780\
        );

    \I__10929\ : InMux
    port map (
            O => \N__51784\,
            I => \N__51772\
        );

    \I__10928\ : InMux
    port map (
            O => \N__51783\,
            I => \N__51769\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__51780\,
            I => \N__51766\
        );

    \I__10926\ : InMux
    port map (
            O => \N__51779\,
            I => \N__51763\
        );

    \I__10925\ : InMux
    port map (
            O => \N__51778\,
            I => \N__51760\
        );

    \I__10924\ : InMux
    port map (
            O => \N__51777\,
            I => \N__51757\
        );

    \I__10923\ : InMux
    port map (
            O => \N__51776\,
            I => \N__51754\
        );

    \I__10922\ : InMux
    port map (
            O => \N__51775\,
            I => \N__51751\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__51772\,
            I => \N__51748\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__51769\,
            I => \N__51743\
        );

    \I__10919\ : Span4Mux_h
    port map (
            O => \N__51766\,
            I => \N__51743\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__51763\,
            I => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__51760\,
            I => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__51757\,
            I => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__51754\,
            I => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__51751\,
            I => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\
        );

    \I__10913\ : Odrv4
    port map (
            O => \N__51748\,
            I => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\
        );

    \I__10912\ : Odrv4
    port map (
            O => \N__51743\,
            I => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\
        );

    \I__10911\ : CascadeMux
    port map (
            O => \N__51728\,
            I => \N__51724\
        );

    \I__10910\ : InMux
    port map (
            O => \N__51727\,
            I => \N__51717\
        );

    \I__10909\ : InMux
    port map (
            O => \N__51724\,
            I => \N__51714\
        );

    \I__10908\ : CascadeMux
    port map (
            O => \N__51723\,
            I => \N__51711\
        );

    \I__10907\ : CascadeMux
    port map (
            O => \N__51722\,
            I => \N__51708\
        );

    \I__10906\ : CascadeMux
    port map (
            O => \N__51721\,
            I => \N__51705\
        );

    \I__10905\ : CascadeMux
    port map (
            O => \N__51720\,
            I => \N__51700\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__51717\,
            I => \N__51695\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__51714\,
            I => \N__51695\
        );

    \I__10902\ : InMux
    port map (
            O => \N__51711\,
            I => \N__51692\
        );

    \I__10901\ : InMux
    port map (
            O => \N__51708\,
            I => \N__51689\
        );

    \I__10900\ : InMux
    port map (
            O => \N__51705\,
            I => \N__51686\
        );

    \I__10899\ : InMux
    port map (
            O => \N__51704\,
            I => \N__51683\
        );

    \I__10898\ : InMux
    port map (
            O => \N__51703\,
            I => \N__51680\
        );

    \I__10897\ : InMux
    port map (
            O => \N__51700\,
            I => \N__51677\
        );

    \I__10896\ : Span4Mux_v
    port map (
            O => \N__51695\,
            I => \N__51674\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__51692\,
            I => \N__51669\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__51689\,
            I => \N__51669\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__51686\,
            I => \N__51660\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__51683\,
            I => \N__51660\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__51680\,
            I => \N__51660\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__51677\,
            I => \N__51660\
        );

    \I__10889\ : Span4Mux_v
    port map (
            O => \N__51674\,
            I => \N__51657\
        );

    \I__10888\ : Span4Mux_v
    port map (
            O => \N__51669\,
            I => \N__51654\
        );

    \I__10887\ : Span12Mux_v
    port map (
            O => \N__51660\,
            I => \N__51649\
        );

    \I__10886\ : Sp12to4
    port map (
            O => \N__51657\,
            I => \N__51649\
        );

    \I__10885\ : Span4Mux_h
    port map (
            O => \N__51654\,
            I => \N__51646\
        );

    \I__10884\ : Span12Mux_s11_h
    port map (
            O => \N__51649\,
            I => \N__51643\
        );

    \I__10883\ : Odrv4
    port map (
            O => \N__51646\,
            I => \ALU.a_15_m3_sZ0Z_13\
        );

    \I__10882\ : Odrv12
    port map (
            O => \N__51643\,
            I => \ALU.a_15_m3_sZ0Z_13\
        );

    \I__10881\ : InMux
    port map (
            O => \N__51638\,
            I => \N__51629\
        );

    \I__10880\ : InMux
    port map (
            O => \N__51637\,
            I => \N__51626\
        );

    \I__10879\ : InMux
    port map (
            O => \N__51636\,
            I => \N__51623\
        );

    \I__10878\ : InMux
    port map (
            O => \N__51635\,
            I => \N__51620\
        );

    \I__10877\ : InMux
    port map (
            O => \N__51634\,
            I => \N__51617\
        );

    \I__10876\ : InMux
    port map (
            O => \N__51633\,
            I => \N__51614\
        );

    \I__10875\ : InMux
    port map (
            O => \N__51632\,
            I => \N__51611\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__51629\,
            I => \N__51608\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__51626\,
            I => \N__51605\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__51623\,
            I => \N__51602\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__51620\,
            I => \ALU.mult_495_c_RNIKOB51JZ0\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__51617\,
            I => \ALU.mult_495_c_RNIKOB51JZ0\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__51614\,
            I => \ALU.mult_495_c_RNIKOB51JZ0\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__51611\,
            I => \ALU.mult_495_c_RNIKOB51JZ0\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__51608\,
            I => \ALU.mult_495_c_RNIKOB51JZ0\
        );

    \I__10866\ : Odrv4
    port map (
            O => \N__51605\,
            I => \ALU.mult_495_c_RNIKOB51JZ0\
        );

    \I__10865\ : Odrv12
    port map (
            O => \N__51602\,
            I => \ALU.mult_495_c_RNIKOB51JZ0\
        );

    \I__10864\ : InMux
    port map (
            O => \N__51587\,
            I => \N__51584\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__51584\,
            I => \N__51581\
        );

    \I__10862\ : Span4Mux_h
    port map (
            O => \N__51581\,
            I => \N__51577\
        );

    \I__10861\ : InMux
    port map (
            O => \N__51580\,
            I => \N__51574\
        );

    \I__10860\ : Span4Mux_h
    port map (
            O => \N__51577\,
            I => \N__51571\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__51574\,
            I => \N__51568\
        );

    \I__10858\ : Span4Mux_h
    port map (
            O => \N__51571\,
            I => \N__51565\
        );

    \I__10857\ : Span12Mux_h
    port map (
            O => \N__51568\,
            I => \N__51562\
        );

    \I__10856\ : Span4Mux_v
    port map (
            O => \N__51565\,
            I => \N__51559\
        );

    \I__10855\ : Odrv12
    port map (
            O => \N__51562\,
            I => \ALU.dZ0Z_8\
        );

    \I__10854\ : Odrv4
    port map (
            O => \N__51559\,
            I => \ALU.dZ0Z_8\
        );

    \I__10853\ : CascadeMux
    port map (
            O => \N__51554\,
            I => \ALU.c_RNIV5AOKZ0Z_13_cascade_\
        );

    \I__10852\ : CascadeMux
    port map (
            O => \N__51551\,
            I => \ALU.c_RNIO5N04A_0Z0Z_13_cascade_\
        );

    \I__10851\ : InMux
    port map (
            O => \N__51548\,
            I => \N__51545\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__51545\,
            I => \N__51542\
        );

    \I__10849\ : Span4Mux_v
    port map (
            O => \N__51542\,
            I => \N__51538\
        );

    \I__10848\ : InMux
    port map (
            O => \N__51541\,
            I => \N__51535\
        );

    \I__10847\ : Span4Mux_v
    port map (
            O => \N__51538\,
            I => \N__51532\
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__51535\,
            I => \N__51529\
        );

    \I__10845\ : Sp12to4
    port map (
            O => \N__51532\,
            I => \N__51526\
        );

    \I__10844\ : Span4Mux_v
    port map (
            O => \N__51529\,
            I => \N__51523\
        );

    \I__10843\ : Span12Mux_h
    port map (
            O => \N__51526\,
            I => \N__51520\
        );

    \I__10842\ : Odrv4
    port map (
            O => \N__51523\,
            I => \ALU.bZ0Z_13\
        );

    \I__10841\ : Odrv12
    port map (
            O => \N__51520\,
            I => \ALU.bZ0Z_13\
        );

    \I__10840\ : InMux
    port map (
            O => \N__51515\,
            I => \N__51512\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__51512\,
            I => \ALU.c_RNIV5AOKZ0Z_13\
        );

    \I__10838\ : CascadeMux
    port map (
            O => \N__51509\,
            I => \N__51506\
        );

    \I__10837\ : InMux
    port map (
            O => \N__51506\,
            I => \N__51503\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__51503\,
            I => \N__51499\
        );

    \I__10835\ : InMux
    port map (
            O => \N__51502\,
            I => \N__51496\
        );

    \I__10834\ : Odrv4
    port map (
            O => \N__51499\,
            I => \ALU.d_RNIRFBHE9Z0Z_0\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__51496\,
            I => \ALU.d_RNIRFBHE9Z0Z_0\
        );

    \I__10832\ : InMux
    port map (
            O => \N__51491\,
            I => \N__51487\
        );

    \I__10831\ : InMux
    port map (
            O => \N__51490\,
            I => \N__51484\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__51487\,
            I => \N__51481\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__51484\,
            I => \N__51478\
        );

    \I__10828\ : Span4Mux_h
    port map (
            O => \N__51481\,
            I => \N__51475\
        );

    \I__10827\ : Span12Mux_v
    port map (
            O => \N__51478\,
            I => \N__51472\
        );

    \I__10826\ : Span4Mux_v
    port map (
            O => \N__51475\,
            I => \N__51469\
        );

    \I__10825\ : Span12Mux_h
    port map (
            O => \N__51472\,
            I => \N__51466\
        );

    \I__10824\ : Odrv4
    port map (
            O => \N__51469\,
            I => \ALU.log_1_4\
        );

    \I__10823\ : Odrv12
    port map (
            O => \N__51466\,
            I => \ALU.log_1_4\
        );

    \I__10822\ : CascadeMux
    port map (
            O => \N__51461\,
            I => \ALU.N_16_0_cascade_\
        );

    \I__10821\ : InMux
    port map (
            O => \N__51458\,
            I => \N__51455\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__51455\,
            I => \N__51452\
        );

    \I__10819\ : Span4Mux_h
    port map (
            O => \N__51452\,
            I => \N__51449\
        );

    \I__10818\ : Span4Mux_h
    port map (
            O => \N__51449\,
            I => \N__51446\
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__51446\,
            I => \ALU.status_8_8_0\
        );

    \I__10816\ : InMux
    port map (
            O => \N__51443\,
            I => \N__51440\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__51440\,
            I => \ALU.log_1_9\
        );

    \I__10814\ : InMux
    port map (
            O => \N__51437\,
            I => \N__51434\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__51434\,
            I => \N__51431\
        );

    \I__10812\ : Span4Mux_h
    port map (
            O => \N__51431\,
            I => \N__51428\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__51428\,
            I => \N__51425\
        );

    \I__10810\ : Odrv4
    port map (
            O => \N__51425\,
            I => \ALU.d_RNI7KS2IZ0Z_9\
        );

    \I__10809\ : CascadeMux
    port map (
            O => \N__51422\,
            I => \N__51418\
        );

    \I__10808\ : CascadeMux
    port map (
            O => \N__51421\,
            I => \N__51415\
        );

    \I__10807\ : InMux
    port map (
            O => \N__51418\,
            I => \N__51412\
        );

    \I__10806\ : InMux
    port map (
            O => \N__51415\,
            I => \N__51409\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__51412\,
            I => \N__51406\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__51409\,
            I => \N__51403\
        );

    \I__10803\ : Span4Mux_h
    port map (
            O => \N__51406\,
            I => \N__51400\
        );

    \I__10802\ : Span4Mux_v
    port map (
            O => \N__51403\,
            I => \N__51397\
        );

    \I__10801\ : Span4Mux_h
    port map (
            O => \N__51400\,
            I => \N__51394\
        );

    \I__10800\ : Span4Mux_h
    port map (
            O => \N__51397\,
            I => \N__51391\
        );

    \I__10799\ : Span4Mux_v
    port map (
            O => \N__51394\,
            I => \N__51388\
        );

    \I__10798\ : Span4Mux_h
    port map (
            O => \N__51391\,
            I => \N__51385\
        );

    \I__10797\ : Span4Mux_h
    port map (
            O => \N__51388\,
            I => \N__51382\
        );

    \I__10796\ : Odrv4
    port map (
            O => \N__51385\,
            I => \ALU.eZ0Z_12\
        );

    \I__10795\ : Odrv4
    port map (
            O => \N__51382\,
            I => \ALU.eZ0Z_12\
        );

    \I__10794\ : CascadeMux
    port map (
            O => \N__51377\,
            I => \PROM.ROMDATA.m58_cascade_\
        );

    \I__10793\ : InMux
    port map (
            O => \N__51374\,
            I => \N__51371\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__51371\,
            I => \PROM.ROMDATA.m64_am\
        );

    \I__10791\ : InMux
    port map (
            O => \N__51368\,
            I => \N__51365\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__51365\,
            I => \N__51362\
        );

    \I__10789\ : Odrv4
    port map (
            O => \N__51362\,
            I => \PROM.ROMDATA.m45\
        );

    \I__10788\ : InMux
    port map (
            O => \N__51359\,
            I => \N__51356\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__51356\,
            I => \N__51353\
        );

    \I__10786\ : Span4Mux_h
    port map (
            O => \N__51353\,
            I => \N__51350\
        );

    \I__10785\ : Span4Mux_v
    port map (
            O => \N__51350\,
            I => \N__51347\
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__51347\,
            I => \ALU.log_1_7\
        );

    \I__10783\ : InMux
    port map (
            O => \N__51344\,
            I => \N__51341\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__51341\,
            I => \N__51338\
        );

    \I__10781\ : Span4Mux_h
    port map (
            O => \N__51338\,
            I => \N__51335\
        );

    \I__10780\ : Span4Mux_h
    port map (
            O => \N__51335\,
            I => \N__51331\
        );

    \I__10779\ : InMux
    port map (
            O => \N__51334\,
            I => \N__51328\
        );

    \I__10778\ : Odrv4
    port map (
            O => \N__51331\,
            I => \ALU.log_1_5\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__51328\,
            I => \ALU.log_1_5\
        );

    \I__10776\ : CascadeMux
    port map (
            O => \N__51323\,
            I => \N__51319\
        );

    \I__10775\ : InMux
    port map (
            O => \N__51322\,
            I => \N__51316\
        );

    \I__10774\ : InMux
    port map (
            O => \N__51319\,
            I => \N__51313\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__51316\,
            I => \N__51310\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__51313\,
            I => \N__51307\
        );

    \I__10771\ : Span4Mux_v
    port map (
            O => \N__51310\,
            I => \N__51304\
        );

    \I__10770\ : Span4Mux_h
    port map (
            O => \N__51307\,
            I => \N__51301\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__51304\,
            I => \ALU.log_1_11\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__51301\,
            I => \ALU.log_1_11\
        );

    \I__10767\ : InMux
    port map (
            O => \N__51296\,
            I => \N__51292\
        );

    \I__10766\ : InMux
    port map (
            O => \N__51295\,
            I => \N__51289\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__51292\,
            I => \N__51286\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__51289\,
            I => \N__51283\
        );

    \I__10763\ : Span4Mux_v
    port map (
            O => \N__51286\,
            I => \N__51280\
        );

    \I__10762\ : Span4Mux_v
    port map (
            O => \N__51283\,
            I => \N__51277\
        );

    \I__10761\ : Span4Mux_v
    port map (
            O => \N__51280\,
            I => \N__51272\
        );

    \I__10760\ : Span4Mux_v
    port map (
            O => \N__51277\,
            I => \N__51272\
        );

    \I__10759\ : Sp12to4
    port map (
            O => \N__51272\,
            I => \N__51269\
        );

    \I__10758\ : Span12Mux_h
    port map (
            O => \N__51269\,
            I => \N__51266\
        );

    \I__10757\ : Odrv12
    port map (
            O => \N__51266\,
            I => \ALU.log_1_10\
        );

    \I__10756\ : InMux
    port map (
            O => \N__51263\,
            I => \N__51259\
        );

    \I__10755\ : InMux
    port map (
            O => \N__51262\,
            I => \N__51256\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__51259\,
            I => \N__51253\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__51256\,
            I => \N__51248\
        );

    \I__10752\ : Span12Mux_v
    port map (
            O => \N__51253\,
            I => \N__51248\
        );

    \I__10751\ : Span12Mux_h
    port map (
            O => \N__51248\,
            I => \N__51245\
        );

    \I__10750\ : Odrv12
    port map (
            O => \N__51245\,
            I => \ALU.N_22_0\
        );

    \I__10749\ : InMux
    port map (
            O => \N__51242\,
            I => \N__51239\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__51239\,
            I => \N__51235\
        );

    \I__10747\ : InMux
    port map (
            O => \N__51238\,
            I => \N__51232\
        );

    \I__10746\ : Span4Mux_h
    port map (
            O => \N__51235\,
            I => \N__51229\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__51232\,
            I => \N__51226\
        );

    \I__10744\ : Span4Mux_v
    port map (
            O => \N__51229\,
            I => \N__51223\
        );

    \I__10743\ : Span4Mux_v
    port map (
            O => \N__51226\,
            I => \N__51220\
        );

    \I__10742\ : Span4Mux_h
    port map (
            O => \N__51223\,
            I => \N__51217\
        );

    \I__10741\ : Span4Mux_h
    port map (
            O => \N__51220\,
            I => \N__51214\
        );

    \I__10740\ : Span4Mux_v
    port map (
            O => \N__51217\,
            I => \N__51211\
        );

    \I__10739\ : Odrv4
    port map (
            O => \N__51214\,
            I => \ALU.N_20_0\
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__51211\,
            I => \ALU.N_20_0\
        );

    \I__10737\ : CascadeMux
    port map (
            O => \N__51206\,
            I => \ALU.status_8_10_0_cascade_\
        );

    \I__10736\ : InMux
    port map (
            O => \N__51203\,
            I => \N__51200\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__51200\,
            I => \N__51197\
        );

    \I__10734\ : Span4Mux_h
    port map (
            O => \N__51197\,
            I => \N__51194\
        );

    \I__10733\ : Span4Mux_h
    port map (
            O => \N__51194\,
            I => \N__51191\
        );

    \I__10732\ : Odrv4
    port map (
            O => \N__51191\,
            I => \ALU.status_8_13_0\
        );

    \I__10731\ : InMux
    port map (
            O => \N__51188\,
            I => \N__51185\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__51185\,
            I => \ALU.status_8_3_1_0\
        );

    \I__10729\ : CascadeMux
    port map (
            O => \N__51182\,
            I => \ALU.log_1_15_cascade_\
        );

    \I__10728\ : InMux
    port map (
            O => \N__51179\,
            I => \N__51176\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__51176\,
            I => \ALU.status_8_13_1_0\
        );

    \I__10726\ : CascadeMux
    port map (
            O => \N__51173\,
            I => \PROM.ROMDATA.m191_cascade_\
        );

    \I__10725\ : InMux
    port map (
            O => \N__51170\,
            I => \N__51167\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__51167\,
            I => \PROM.ROMDATA.m193\
        );

    \I__10723\ : InMux
    port map (
            O => \N__51164\,
            I => \N__51161\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__51161\,
            I => \PROM.ROMDATA.m195_bm\
        );

    \I__10721\ : InMux
    port map (
            O => \N__51158\,
            I => \N__51155\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__51155\,
            I => \N__51152\
        );

    \I__10719\ : Span4Mux_v
    port map (
            O => \N__51152\,
            I => \N__51149\
        );

    \I__10718\ : Span4Mux_h
    port map (
            O => \N__51149\,
            I => \N__51145\
        );

    \I__10717\ : InMux
    port map (
            O => \N__51148\,
            I => \N__51142\
        );

    \I__10716\ : Span4Mux_h
    port map (
            O => \N__51145\,
            I => \N__51139\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__51142\,
            I => \N__51136\
        );

    \I__10714\ : Span4Mux_v
    port map (
            O => \N__51139\,
            I => \N__51133\
        );

    \I__10713\ : Span4Mux_h
    port map (
            O => \N__51136\,
            I => \N__51130\
        );

    \I__10712\ : Odrv4
    port map (
            O => \N__51133\,
            I => \CONTROL.programCounter_1_3\
        );

    \I__10711\ : Odrv4
    port map (
            O => \N__51130\,
            I => \CONTROL.programCounter_1_3\
        );

    \I__10710\ : InMux
    port map (
            O => \N__51125\,
            I => \N__51122\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__51122\,
            I => \N__51118\
        );

    \I__10708\ : InMux
    port map (
            O => \N__51121\,
            I => \N__51115\
        );

    \I__10707\ : Span4Mux_h
    port map (
            O => \N__51118\,
            I => \N__51110\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__51115\,
            I => \N__51110\
        );

    \I__10705\ : Odrv4
    port map (
            O => \N__51110\,
            I => \CONTROL.programCounter_1_reto_3\
        );

    \I__10704\ : InMux
    port map (
            O => \N__51107\,
            I => \N__51104\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__51104\,
            I => \N__51101\
        );

    \I__10702\ : Odrv12
    port map (
            O => \N__51101\,
            I => \PROM.ROMDATA.m92_am\
        );

    \I__10701\ : CascadeMux
    port map (
            O => \N__51098\,
            I => \PROM.ROMDATA.m62_cascade_\
        );

    \I__10700\ : InMux
    port map (
            O => \N__51095\,
            I => \N__51092\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__51092\,
            I => \N__51089\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__51089\,
            I => \PROM.ROMDATA.m53_am\
        );

    \I__10697\ : CascadeMux
    port map (
            O => \N__51086\,
            I => \N__51083\
        );

    \I__10696\ : InMux
    port map (
            O => \N__51083\,
            I => \N__51080\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__51080\,
            I => \N__51077\
        );

    \I__10694\ : Odrv4
    port map (
            O => \N__51077\,
            I => \PROM.ROMDATA.m53_bm\
        );

    \I__10693\ : InMux
    port map (
            O => \N__51074\,
            I => \N__51071\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__51071\,
            I => \PROM.ROMDATA.m64_bm\
        );

    \I__10691\ : CascadeMux
    port map (
            O => \N__51068\,
            I => \PROM.ROMDATA.m65_ns_1_cascade_\
        );

    \I__10690\ : InMux
    port map (
            O => \N__51065\,
            I => \N__51059\
        );

    \I__10689\ : InMux
    port map (
            O => \N__51064\,
            I => \N__51059\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__51059\,
            I => \N__51056\
        );

    \I__10687\ : Span4Mux_h
    port map (
            O => \N__51056\,
            I => \N__51053\
        );

    \I__10686\ : Odrv4
    port map (
            O => \N__51053\,
            I => m65_ns
        );

    \I__10685\ : CascadeMux
    port map (
            O => \N__51050\,
            I => \PROM.ROMDATA.m80_am_cascade_\
        );

    \I__10684\ : InMux
    port map (
            O => \N__51047\,
            I => \N__51044\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__51044\,
            I => \N__51041\
        );

    \I__10682\ : Span4Mux_v
    port map (
            O => \N__51041\,
            I => \N__51038\
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__51038\,
            I => \PROM.ROMDATA.m93_ns_1\
        );

    \I__10680\ : InMux
    port map (
            O => \N__51035\,
            I => \N__51032\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__51032\,
            I => \CONTROL.programCounter_ret_1_RNIJ88IZ0Z_2\
        );

    \I__10678\ : InMux
    port map (
            O => \N__51029\,
            I => \N__51026\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__51026\,
            I => \CONTROL.programCounter_ret_19_RNICM8JZ0Z_2\
        );

    \I__10676\ : CascadeMux
    port map (
            O => \N__51023\,
            I => \progRomAddress_2_cascade_\
        );

    \I__10675\ : InMux
    port map (
            O => \N__51020\,
            I => \N__51017\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__51017\,
            I => \N__51014\
        );

    \I__10673\ : Span4Mux_v
    port map (
            O => \N__51014\,
            I => \N__51011\
        );

    \I__10672\ : Odrv4
    port map (
            O => \N__51011\,
            I => \PROM.ROMDATA.m195_am\
        );

    \I__10671\ : CascadeMux
    port map (
            O => \N__51008\,
            I => \PROM.ROMDATA.m196_ns_1_cascade_\
        );

    \I__10670\ : InMux
    port map (
            O => \N__51005\,
            I => \N__51002\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__51002\,
            I => \N__50999\
        );

    \I__10668\ : Odrv4
    port map (
            O => \N__50999\,
            I => \PROM.ROMDATA.m179\
        );

    \I__10667\ : InMux
    port map (
            O => \N__50996\,
            I => \N__50993\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__50993\,
            I => \PROM.ROMDATA.m185_am\
        );

    \I__10665\ : InMux
    port map (
            O => \N__50990\,
            I => \N__50987\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__50987\,
            I => \N__50983\
        );

    \I__10663\ : InMux
    port map (
            O => \N__50986\,
            I => \N__50980\
        );

    \I__10662\ : Span4Mux_h
    port map (
            O => \N__50983\,
            I => \N__50977\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__50980\,
            I => \N__50974\
        );

    \I__10660\ : Odrv4
    port map (
            O => \N__50977\,
            I => \CONTROL.dout_reto_0\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__50974\,
            I => \CONTROL.dout_reto_0\
        );

    \I__10658\ : InMux
    port map (
            O => \N__50969\,
            I => \N__50966\
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__50966\,
            I => \N__50963\
        );

    \I__10656\ : Span4Mux_h
    port map (
            O => \N__50963\,
            I => \N__50959\
        );

    \I__10655\ : InMux
    port map (
            O => \N__50962\,
            I => \N__50956\
        );

    \I__10654\ : Sp12to4
    port map (
            O => \N__50959\,
            I => \N__50952\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__50956\,
            I => \N__50949\
        );

    \I__10652\ : InMux
    port map (
            O => \N__50955\,
            I => \N__50944\
        );

    \I__10651\ : Span12Mux_v
    port map (
            O => \N__50952\,
            I => \N__50941\
        );

    \I__10650\ : Span4Mux_h
    port map (
            O => \N__50949\,
            I => \N__50938\
        );

    \I__10649\ : InMux
    port map (
            O => \N__50948\,
            I => \N__50935\
        );

    \I__10648\ : InMux
    port map (
            O => \N__50947\,
            I => \N__50932\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__50944\,
            I => \CONTROL_addrstack_reto_0\
        );

    \I__10646\ : Odrv12
    port map (
            O => \N__50941\,
            I => \CONTROL_addrstack_reto_0\
        );

    \I__10645\ : Odrv4
    port map (
            O => \N__50938\,
            I => \CONTROL_addrstack_reto_0\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__50935\,
            I => \CONTROL_addrstack_reto_0\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__50932\,
            I => \CONTROL_addrstack_reto_0\
        );

    \I__10642\ : CascadeMux
    port map (
            O => \N__50921\,
            I => \N__50918\
        );

    \I__10641\ : InMux
    port map (
            O => \N__50918\,
            I => \N__50915\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__50915\,
            I => \N__50912\
        );

    \I__10639\ : Span4Mux_v
    port map (
            O => \N__50912\,
            I => \N__50909\
        );

    \I__10638\ : Odrv4
    port map (
            O => \N__50909\,
            I => \PROM.ROMDATA.m248_ns_1\
        );

    \I__10637\ : InMux
    port map (
            O => \N__50906\,
            I => \N__50900\
        );

    \I__10636\ : InMux
    port map (
            O => \N__50905\,
            I => \N__50893\
        );

    \I__10635\ : InMux
    port map (
            O => \N__50904\,
            I => \N__50893\
        );

    \I__10634\ : InMux
    port map (
            O => \N__50903\,
            I => \N__50890\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__50900\,
            I => \N__50887\
        );

    \I__10632\ : InMux
    port map (
            O => \N__50899\,
            I => \N__50884\
        );

    \I__10631\ : InMux
    port map (
            O => \N__50898\,
            I => \N__50881\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__50893\,
            I => \N__50876\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__50890\,
            I => \N__50876\
        );

    \I__10628\ : Span4Mux_v
    port map (
            O => \N__50887\,
            I => \N__50873\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__50884\,
            I => \N__50866\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__50881\,
            I => \N__50866\
        );

    \I__10625\ : Span4Mux_h
    port map (
            O => \N__50876\,
            I => \N__50863\
        );

    \I__10624\ : Span4Mux_h
    port map (
            O => \N__50873\,
            I => \N__50860\
        );

    \I__10623\ : InMux
    port map (
            O => \N__50872\,
            I => \N__50855\
        );

    \I__10622\ : InMux
    port map (
            O => \N__50871\,
            I => \N__50855\
        );

    \I__10621\ : Span4Mux_v
    port map (
            O => \N__50866\,
            I => \N__50850\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__50863\,
            I => \N__50850\
        );

    \I__10619\ : Odrv4
    port map (
            O => \N__50860\,
            I => \CONTROL.incrementZ0Z_0\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__50855\,
            I => \CONTROL.incrementZ0Z_0\
        );

    \I__10617\ : Odrv4
    port map (
            O => \N__50850\,
            I => \CONTROL.incrementZ0Z_0\
        );

    \I__10616\ : CascadeMux
    port map (
            O => \N__50843\,
            I => \N__50838\
        );

    \I__10615\ : CascadeMux
    port map (
            O => \N__50842\,
            I => \N__50831\
        );

    \I__10614\ : InMux
    port map (
            O => \N__50841\,
            I => \N__50827\
        );

    \I__10613\ : InMux
    port map (
            O => \N__50838\,
            I => \N__50822\
        );

    \I__10612\ : InMux
    port map (
            O => \N__50837\,
            I => \N__50822\
        );

    \I__10611\ : InMux
    port map (
            O => \N__50836\,
            I => \N__50819\
        );

    \I__10610\ : InMux
    port map (
            O => \N__50835\,
            I => \N__50816\
        );

    \I__10609\ : InMux
    port map (
            O => \N__50834\,
            I => \N__50813\
        );

    \I__10608\ : InMux
    port map (
            O => \N__50831\,
            I => \N__50808\
        );

    \I__10607\ : InMux
    port map (
            O => \N__50830\,
            I => \N__50808\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__50827\,
            I => \N__50805\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__50822\,
            I => \N__50800\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__50819\,
            I => \N__50800\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__50816\,
            I => \N__50797\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__50813\,
            I => \N__50794\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__50808\,
            I => \N__50791\
        );

    \I__10600\ : Span4Mux_v
    port map (
            O => \N__50805\,
            I => \N__50788\
        );

    \I__10599\ : Span4Mux_v
    port map (
            O => \N__50800\,
            I => \N__50785\
        );

    \I__10598\ : Span4Mux_v
    port map (
            O => \N__50797\,
            I => \N__50782\
        );

    \I__10597\ : Span4Mux_h
    port map (
            O => \N__50794\,
            I => \N__50775\
        );

    \I__10596\ : Span4Mux_v
    port map (
            O => \N__50791\,
            I => \N__50775\
        );

    \I__10595\ : Span4Mux_h
    port map (
            O => \N__50788\,
            I => \N__50775\
        );

    \I__10594\ : Span4Mux_h
    port map (
            O => \N__50785\,
            I => \N__50772\
        );

    \I__10593\ : Span4Mux_h
    port map (
            O => \N__50782\,
            I => \N__50767\
        );

    \I__10592\ : Span4Mux_v
    port map (
            O => \N__50775\,
            I => \N__50767\
        );

    \I__10591\ : Span4Mux_h
    port map (
            O => \N__50772\,
            I => \N__50764\
        );

    \I__10590\ : Odrv4
    port map (
            O => \N__50767\,
            I => \CONTROL.incrementZ0Z_1\
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__50764\,
            I => \CONTROL.incrementZ0Z_1\
        );

    \I__10588\ : InMux
    port map (
            O => \N__50759\,
            I => \N__50756\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__50756\,
            I => \N__50753\
        );

    \I__10586\ : Span4Mux_h
    port map (
            O => \N__50753\,
            I => \N__50750\
        );

    \I__10585\ : Odrv4
    port map (
            O => \N__50750\,
            I => \PROM.ROMDATA.m284_1\
        );

    \I__10584\ : InMux
    port map (
            O => \N__50747\,
            I => \N__50744\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__50744\,
            I => \CONTROL.programCounter_ret_19_RNI8I8JZ0Z_0\
        );

    \I__10582\ : InMux
    port map (
            O => \N__50741\,
            I => \N__50738\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__50738\,
            I => \CONTROL.programCounter_ret_1_RNIF48IZ0Z_0\
        );

    \I__10580\ : CascadeMux
    port map (
            O => \N__50735\,
            I => \progRomAddress_0_cascade_\
        );

    \I__10579\ : CascadeMux
    port map (
            O => \N__50732\,
            I => \PROM.ROMDATA.m72_cascade_\
        );

    \I__10578\ : InMux
    port map (
            O => \N__50729\,
            I => \N__50726\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__50726\,
            I => \PROM.ROMDATA.m74\
        );

    \I__10576\ : CascadeMux
    port map (
            O => \N__50723\,
            I => \PROM.ROMDATA.m169_cascade_\
        );

    \I__10575\ : InMux
    port map (
            O => \N__50720\,
            I => \N__50717\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__50717\,
            I => \N__50714\
        );

    \I__10573\ : Span4Mux_h
    port map (
            O => \N__50714\,
            I => \N__50710\
        );

    \I__10572\ : InMux
    port map (
            O => \N__50713\,
            I => \N__50707\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__50710\,
            I => \N__50704\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__50707\,
            I => \N__50701\
        );

    \I__10569\ : Odrv4
    port map (
            O => \N__50704\,
            I => \PROM.ROMDATA.m270_am\
        );

    \I__10568\ : Odrv12
    port map (
            O => \N__50701\,
            I => \PROM.ROMDATA.m270_am\
        );

    \I__10567\ : CascadeMux
    port map (
            O => \N__50696\,
            I => \PROM.ROMDATA.m13_cascade_\
        );

    \I__10566\ : InMux
    port map (
            O => \N__50693\,
            I => \N__50690\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__50690\,
            I => \PROM.ROMDATA.m188\
        );

    \I__10564\ : CascadeMux
    port map (
            O => \N__50687\,
            I => \N__50684\
        );

    \I__10563\ : InMux
    port map (
            O => \N__50684\,
            I => \N__50681\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__50681\,
            I => \PROM.ROMDATA.m13\
        );

    \I__10561\ : InMux
    port map (
            O => \N__50678\,
            I => \N__50675\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__50675\,
            I => \PROM.ROMDATA.m263\
        );

    \I__10559\ : InMux
    port map (
            O => \N__50672\,
            I => \N__50669\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__50669\,
            I => \N__50666\
        );

    \I__10557\ : Span4Mux_v
    port map (
            O => \N__50666\,
            I => \N__50663\
        );

    \I__10556\ : Span4Mux_h
    port map (
            O => \N__50663\,
            I => \N__50659\
        );

    \I__10555\ : InMux
    port map (
            O => \N__50662\,
            I => \N__50656\
        );

    \I__10554\ : Odrv4
    port map (
            O => \N__50659\,
            I => \CONTROL.ctrlOut_1\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__50656\,
            I => \CONTROL.ctrlOut_1\
        );

    \I__10552\ : CascadeMux
    port map (
            O => \N__50651\,
            I => \PROM.ROMDATA.m150_cascade_\
        );

    \I__10551\ : CascadeMux
    port map (
            O => \N__50648\,
            I => \PROM.ROMDATA.m228_am_cascade_\
        );

    \I__10550\ : CascadeMux
    port map (
            O => \N__50645\,
            I => \N__50642\
        );

    \I__10549\ : InMux
    port map (
            O => \N__50642\,
            I => \N__50639\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__50639\,
            I => \N__50636\
        );

    \I__10547\ : Odrv4
    port map (
            O => \N__50636\,
            I => \PROM.ROMDATA.m25\
        );

    \I__10546\ : InMux
    port map (
            O => \N__50633\,
            I => \N__50630\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__50630\,
            I => \N__50627\
        );

    \I__10544\ : Span4Mux_v
    port map (
            O => \N__50627\,
            I => \N__50624\
        );

    \I__10543\ : Odrv4
    port map (
            O => \N__50624\,
            I => \PROM.ROMDATA.m280\
        );

    \I__10542\ : CascadeMux
    port map (
            O => \N__50621\,
            I => \N__50617\
        );

    \I__10541\ : InMux
    port map (
            O => \N__50620\,
            I => \N__50612\
        );

    \I__10540\ : InMux
    port map (
            O => \N__50617\,
            I => \N__50612\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__50612\,
            I => \N__50609\
        );

    \I__10538\ : Span4Mux_v
    port map (
            O => \N__50609\,
            I => \N__50606\
        );

    \I__10537\ : Span4Mux_h
    port map (
            O => \N__50606\,
            I => \N__50603\
        );

    \I__10536\ : Span4Mux_h
    port map (
            O => \N__50603\,
            I => \N__50600\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__50600\,
            I => \N__50597\
        );

    \I__10534\ : Span4Mux_v
    port map (
            O => \N__50597\,
            I => \N__50594\
        );

    \I__10533\ : Odrv4
    port map (
            O => \N__50594\,
            I => \PROM.ROMDATA.m438\
        );

    \I__10532\ : InMux
    port map (
            O => \N__50591\,
            I => \N__50587\
        );

    \I__10531\ : InMux
    port map (
            O => \N__50590\,
            I => \N__50584\
        );

    \I__10530\ : LocalMux
    port map (
            O => \N__50587\,
            I => \PROM.ROMDATA.m173\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__50584\,
            I => \PROM.ROMDATA.m173\
        );

    \I__10528\ : InMux
    port map (
            O => \N__50579\,
            I => \N__50576\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__50576\,
            I => \N__50573\
        );

    \I__10526\ : Span4Mux_v
    port map (
            O => \N__50573\,
            I => \N__50569\
        );

    \I__10525\ : InMux
    port map (
            O => \N__50572\,
            I => \N__50566\
        );

    \I__10524\ : Odrv4
    port map (
            O => \N__50569\,
            I => \PROM.ROMDATA.m23\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__50566\,
            I => \PROM.ROMDATA.m23\
        );

    \I__10522\ : InMux
    port map (
            O => \N__50561\,
            I => \N__50558\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__50558\,
            I => \N__50555\
        );

    \I__10520\ : Span4Mux_v
    port map (
            O => \N__50555\,
            I => \N__50552\
        );

    \I__10519\ : Span4Mux_h
    port map (
            O => \N__50552\,
            I => \N__50549\
        );

    \I__10518\ : Span4Mux_h
    port map (
            O => \N__50549\,
            I => \N__50546\
        );

    \I__10517\ : Odrv4
    port map (
            O => \N__50546\,
            I => \PROM_ROMDATA_dintern_31_0__g1\
        );

    \I__10516\ : CascadeMux
    port map (
            O => \N__50543\,
            I => \N__50538\
        );

    \I__10515\ : InMux
    port map (
            O => \N__50542\,
            I => \N__50532\
        );

    \I__10514\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50532\
        );

    \I__10513\ : InMux
    port map (
            O => \N__50538\,
            I => \N__50527\
        );

    \I__10512\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50527\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__50532\,
            I => \N__50524\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__50527\,
            I => \N__50521\
        );

    \I__10509\ : Odrv4
    port map (
            O => \N__50524\,
            I => \ALU.a_15_m2_d_d_sZ0Z_0\
        );

    \I__10508\ : Odrv4
    port map (
            O => \N__50521\,
            I => \ALU.a_15_m2_d_d_sZ0Z_0\
        );

    \I__10507\ : CascadeMux
    port map (
            O => \N__50516\,
            I => \bus_15_cascade_\
        );

    \I__10506\ : InMux
    port map (
            O => \N__50513\,
            I => \N__50507\
        );

    \I__10505\ : InMux
    port map (
            O => \N__50512\,
            I => \N__50507\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__50507\,
            I => \ALU.c_RNIJI6SHZ0Z_15\
        );

    \I__10503\ : InMux
    port map (
            O => \N__50504\,
            I => \N__50501\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__50501\,
            I => \ALU.c_RNID85GQZ0Z_15\
        );

    \I__10501\ : CascadeMux
    port map (
            O => \N__50498\,
            I => \PROM.ROMDATA.m248_ns_cascade_\
        );

    \I__10500\ : CascadeMux
    port map (
            O => \N__50495\,
            I => \N__50491\
        );

    \I__10499\ : CascadeMux
    port map (
            O => \N__50494\,
            I => \N__50488\
        );

    \I__10498\ : InMux
    port map (
            O => \N__50491\,
            I => \N__50477\
        );

    \I__10497\ : InMux
    port map (
            O => \N__50488\,
            I => \N__50477\
        );

    \I__10496\ : InMux
    port map (
            O => \N__50487\,
            I => \N__50477\
        );

    \I__10495\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50477\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__50477\,
            I => \N__50474\
        );

    \I__10493\ : Span4Mux_v
    port map (
            O => \N__50474\,
            I => \N__50471\
        );

    \I__10492\ : Span4Mux_h
    port map (
            O => \N__50471\,
            I => \N__50467\
        );

    \I__10491\ : InMux
    port map (
            O => \N__50470\,
            I => \N__50464\
        );

    \I__10490\ : Span4Mux_v
    port map (
            O => \N__50467\,
            I => \N__50461\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__50464\,
            I => \N__50458\
        );

    \I__10488\ : Span4Mux_h
    port map (
            O => \N__50461\,
            I => \N__50455\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__50458\,
            I => \N__50452\
        );

    \I__10486\ : Odrv4
    port map (
            O => \N__50455\,
            I => \PROM.ROMDATA.m249\
        );

    \I__10485\ : Odrv4
    port map (
            O => \N__50452\,
            I => \PROM.ROMDATA.m249\
        );

    \I__10484\ : InMux
    port map (
            O => \N__50447\,
            I => \N__50444\
        );

    \I__10483\ : LocalMux
    port map (
            O => \N__50444\,
            I => \N__50441\
        );

    \I__10482\ : Odrv4
    port map (
            O => \N__50441\,
            I => \PROM.ROMDATA.m359\
        );

    \I__10481\ : InMux
    port map (
            O => \N__50438\,
            I => \N__50435\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__50435\,
            I => \N__50432\
        );

    \I__10479\ : Span4Mux_v
    port map (
            O => \N__50432\,
            I => \N__50427\
        );

    \I__10478\ : InMux
    port map (
            O => \N__50431\,
            I => \N__50422\
        );

    \I__10477\ : InMux
    port map (
            O => \N__50430\,
            I => \N__50422\
        );

    \I__10476\ : Span4Mux_v
    port map (
            O => \N__50427\,
            I => \N__50417\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__50422\,
            I => \N__50417\
        );

    \I__10474\ : Span4Mux_h
    port map (
            O => \N__50417\,
            I => \N__50414\
        );

    \I__10473\ : Span4Mux_h
    port map (
            O => \N__50414\,
            I => \N__50411\
        );

    \I__10472\ : Span4Mux_h
    port map (
            O => \N__50411\,
            I => \N__50408\
        );

    \I__10471\ : Odrv4
    port map (
            O => \N__50408\,
            I => g_8
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__50405\,
            I => \N__50401\
        );

    \I__10469\ : CascadeMux
    port map (
            O => \N__50404\,
            I => \N__50397\
        );

    \I__10468\ : InMux
    port map (
            O => \N__50401\,
            I => \N__50394\
        );

    \I__10467\ : InMux
    port map (
            O => \N__50400\,
            I => \N__50389\
        );

    \I__10466\ : InMux
    port map (
            O => \N__50397\,
            I => \N__50389\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__50394\,
            I => \N__50386\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__50389\,
            I => \N__50383\
        );

    \I__10463\ : Span4Mux_v
    port map (
            O => \N__50386\,
            I => \N__50380\
        );

    \I__10462\ : Span4Mux_v
    port map (
            O => \N__50383\,
            I => \N__50377\
        );

    \I__10461\ : Span4Mux_h
    port map (
            O => \N__50380\,
            I => \N__50374\
        );

    \I__10460\ : Span4Mux_h
    port map (
            O => \N__50377\,
            I => \N__50371\
        );

    \I__10459\ : Span4Mux_h
    port map (
            O => \N__50374\,
            I => \N__50368\
        );

    \I__10458\ : Span4Mux_h
    port map (
            O => \N__50371\,
            I => \N__50365\
        );

    \I__10457\ : Span4Mux_v
    port map (
            O => \N__50368\,
            I => \N__50362\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__50365\,
            I => \N__50359\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__50362\,
            I => g_15
        );

    \I__10454\ : Odrv4
    port map (
            O => \N__50359\,
            I => g_15
        );

    \I__10453\ : CascadeMux
    port map (
            O => \N__50354\,
            I => \ALU.c_RNID85GQ_0Z0Z_15_cascade_\
        );

    \I__10452\ : InMux
    port map (
            O => \N__50351\,
            I => \N__50348\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__50348\,
            I => \N__50345\
        );

    \I__10450\ : Odrv12
    port map (
            O => \N__50345\,
            I => \ALU.c_RNI9DCRE2Z0Z_15\
        );

    \I__10449\ : InMux
    port map (
            O => \N__50342\,
            I => \N__50338\
        );

    \I__10448\ : InMux
    port map (
            O => \N__50341\,
            I => \N__50334\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__50338\,
            I => \N__50331\
        );

    \I__10446\ : InMux
    port map (
            O => \N__50337\,
            I => \N__50328\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__50334\,
            I => \N__50321\
        );

    \I__10444\ : Span4Mux_v
    port map (
            O => \N__50331\,
            I => \N__50318\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__50328\,
            I => \N__50315\
        );

    \I__10442\ : InMux
    port map (
            O => \N__50327\,
            I => \N__50312\
        );

    \I__10441\ : InMux
    port map (
            O => \N__50326\,
            I => \N__50309\
        );

    \I__10440\ : InMux
    port map (
            O => \N__50325\,
            I => \N__50306\
        );

    \I__10439\ : InMux
    port map (
            O => \N__50324\,
            I => \N__50302\
        );

    \I__10438\ : Span4Mux_v
    port map (
            O => \N__50321\,
            I => \N__50299\
        );

    \I__10437\ : Span4Mux_h
    port map (
            O => \N__50318\,
            I => \N__50293\
        );

    \I__10436\ : Span4Mux_v
    port map (
            O => \N__50315\,
            I => \N__50293\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__50312\,
            I => \N__50290\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__50309\,
            I => \N__50287\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__50306\,
            I => \N__50284\
        );

    \I__10432\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50281\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__50302\,
            I => \N__50277\
        );

    \I__10430\ : Span4Mux_v
    port map (
            O => \N__50299\,
            I => \N__50274\
        );

    \I__10429\ : InMux
    port map (
            O => \N__50298\,
            I => \N__50271\
        );

    \I__10428\ : Span4Mux_h
    port map (
            O => \N__50293\,
            I => \N__50266\
        );

    \I__10427\ : Span4Mux_v
    port map (
            O => \N__50290\,
            I => \N__50266\
        );

    \I__10426\ : Span12Mux_h
    port map (
            O => \N__50287\,
            I => \N__50259\
        );

    \I__10425\ : Sp12to4
    port map (
            O => \N__50284\,
            I => \N__50259\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__50281\,
            I => \N__50259\
        );

    \I__10423\ : InMux
    port map (
            O => \N__50280\,
            I => \N__50256\
        );

    \I__10422\ : Odrv12
    port map (
            O => \N__50277\,
            I => \DROM_ROMDATA_dintern_adflt\
        );

    \I__10421\ : Odrv4
    port map (
            O => \N__50274\,
            I => \DROM_ROMDATA_dintern_adflt\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__50271\,
            I => \DROM_ROMDATA_dintern_adflt\
        );

    \I__10419\ : Odrv4
    port map (
            O => \N__50266\,
            I => \DROM_ROMDATA_dintern_adflt\
        );

    \I__10418\ : Odrv12
    port map (
            O => \N__50259\,
            I => \DROM_ROMDATA_dintern_adflt\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__50256\,
            I => \DROM_ROMDATA_dintern_adflt\
        );

    \I__10416\ : CascadeMux
    port map (
            O => \N__50243\,
            I => \N__50240\
        );

    \I__10415\ : InMux
    port map (
            O => \N__50240\,
            I => \N__50237\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__50237\,
            I => \N__50234\
        );

    \I__10413\ : Span12Mux_v
    port map (
            O => \N__50234\,
            I => \N__50231\
        );

    \I__10412\ : Span12Mux_h
    port map (
            O => \N__50231\,
            I => \N__50228\
        );

    \I__10411\ : Odrv12
    port map (
            O => \N__50228\,
            I => \DROM_ROMDATA_dintern_15ro\
        );

    \I__10410\ : InMux
    port map (
            O => \N__50225\,
            I => \N__50204\
        );

    \I__10409\ : InMux
    port map (
            O => \N__50224\,
            I => \N__50204\
        );

    \I__10408\ : InMux
    port map (
            O => \N__50223\,
            I => \N__50204\
        );

    \I__10407\ : InMux
    port map (
            O => \N__50222\,
            I => \N__50204\
        );

    \I__10406\ : InMux
    port map (
            O => \N__50221\,
            I => \N__50194\
        );

    \I__10405\ : InMux
    port map (
            O => \N__50220\,
            I => \N__50191\
        );

    \I__10404\ : InMux
    port map (
            O => \N__50219\,
            I => \N__50187\
        );

    \I__10403\ : InMux
    port map (
            O => \N__50218\,
            I => \N__50183\
        );

    \I__10402\ : InMux
    port map (
            O => \N__50217\,
            I => \N__50178\
        );

    \I__10401\ : InMux
    port map (
            O => \N__50216\,
            I => \N__50178\
        );

    \I__10400\ : InMux
    port map (
            O => \N__50215\,
            I => \N__50175\
        );

    \I__10399\ : InMux
    port map (
            O => \N__50214\,
            I => \N__50172\
        );

    \I__10398\ : InMux
    port map (
            O => \N__50213\,
            I => \N__50169\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__50204\,
            I => \N__50165\
        );

    \I__10396\ : InMux
    port map (
            O => \N__50203\,
            I => \N__50158\
        );

    \I__10395\ : InMux
    port map (
            O => \N__50202\,
            I => \N__50158\
        );

    \I__10394\ : InMux
    port map (
            O => \N__50201\,
            I => \N__50158\
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__50200\,
            I => \N__50149\
        );

    \I__10392\ : InMux
    port map (
            O => \N__50199\,
            I => \N__50144\
        );

    \I__10391\ : InMux
    port map (
            O => \N__50198\,
            I => \N__50138\
        );

    \I__10390\ : InMux
    port map (
            O => \N__50197\,
            I => \N__50138\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__50194\,
            I => \N__50133\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__50191\,
            I => \N__50133\
        );

    \I__10387\ : InMux
    port map (
            O => \N__50190\,
            I => \N__50128\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__50187\,
            I => \N__50120\
        );

    \I__10385\ : CascadeMux
    port map (
            O => \N__50186\,
            I => \N__50117\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__50183\,
            I => \N__50114\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__50178\,
            I => \N__50108\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__50175\,
            I => \N__50095\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__50172\,
            I => \N__50095\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__50169\,
            I => \N__50095\
        );

    \I__10379\ : InMux
    port map (
            O => \N__50168\,
            I => \N__50092\
        );

    \I__10378\ : Span4Mux_v
    port map (
            O => \N__50165\,
            I => \N__50087\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__50158\,
            I => \N__50087\
        );

    \I__10376\ : InMux
    port map (
            O => \N__50157\,
            I => \N__50084\
        );

    \I__10375\ : InMux
    port map (
            O => \N__50156\,
            I => \N__50077\
        );

    \I__10374\ : InMux
    port map (
            O => \N__50155\,
            I => \N__50077\
        );

    \I__10373\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50077\
        );

    \I__10372\ : InMux
    port map (
            O => \N__50153\,
            I => \N__50074\
        );

    \I__10371\ : InMux
    port map (
            O => \N__50152\,
            I => \N__50071\
        );

    \I__10370\ : InMux
    port map (
            O => \N__50149\,
            I => \N__50068\
        );

    \I__10369\ : InMux
    port map (
            O => \N__50148\,
            I => \N__50063\
        );

    \I__10368\ : InMux
    port map (
            O => \N__50147\,
            I => \N__50063\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__50144\,
            I => \N__50060\
        );

    \I__10366\ : InMux
    port map (
            O => \N__50143\,
            I => \N__50057\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__50138\,
            I => \N__50052\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__50133\,
            I => \N__50052\
        );

    \I__10363\ : InMux
    port map (
            O => \N__50132\,
            I => \N__50047\
        );

    \I__10362\ : InMux
    port map (
            O => \N__50131\,
            I => \N__50047\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__50128\,
            I => \N__50044\
        );

    \I__10360\ : InMux
    port map (
            O => \N__50127\,
            I => \N__50041\
        );

    \I__10359\ : InMux
    port map (
            O => \N__50126\,
            I => \N__50032\
        );

    \I__10358\ : InMux
    port map (
            O => \N__50125\,
            I => \N__50032\
        );

    \I__10357\ : InMux
    port map (
            O => \N__50124\,
            I => \N__50032\
        );

    \I__10356\ : InMux
    port map (
            O => \N__50123\,
            I => \N__50032\
        );

    \I__10355\ : Span4Mux_v
    port map (
            O => \N__50120\,
            I => \N__50029\
        );

    \I__10354\ : InMux
    port map (
            O => \N__50117\,
            I => \N__50026\
        );

    \I__10353\ : Span12Mux_h
    port map (
            O => \N__50114\,
            I => \N__50023\
        );

    \I__10352\ : InMux
    port map (
            O => \N__50113\,
            I => \N__50012\
        );

    \I__10351\ : InMux
    port map (
            O => \N__50112\,
            I => \N__50012\
        );

    \I__10350\ : InMux
    port map (
            O => \N__50111\,
            I => \N__50012\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__50108\,
            I => \N__50000\
        );

    \I__10348\ : InMux
    port map (
            O => \N__50107\,
            I => \N__49991\
        );

    \I__10347\ : InMux
    port map (
            O => \N__50106\,
            I => \N__49991\
        );

    \I__10346\ : InMux
    port map (
            O => \N__50105\,
            I => \N__49991\
        );

    \I__10345\ : InMux
    port map (
            O => \N__50104\,
            I => \N__49991\
        );

    \I__10344\ : InMux
    port map (
            O => \N__50103\,
            I => \N__49986\
        );

    \I__10343\ : InMux
    port map (
            O => \N__50102\,
            I => \N__49986\
        );

    \I__10342\ : Span4Mux_h
    port map (
            O => \N__50095\,
            I => \N__49979\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__50092\,
            I => \N__49979\
        );

    \I__10340\ : Span4Mux_h
    port map (
            O => \N__50087\,
            I => \N__49979\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__50084\,
            I => \N__49974\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__50077\,
            I => \N__49974\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__50074\,
            I => \N__49969\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__50071\,
            I => \N__49969\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__50068\,
            I => \N__49956\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__50063\,
            I => \N__49956\
        );

    \I__10333\ : Span4Mux_h
    port map (
            O => \N__50060\,
            I => \N__49956\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__50057\,
            I => \N__49956\
        );

    \I__10331\ : Span4Mux_v
    port map (
            O => \N__50052\,
            I => \N__49956\
        );

    \I__10330\ : LocalMux
    port map (
            O => \N__50047\,
            I => \N__49956\
        );

    \I__10329\ : Span4Mux_v
    port map (
            O => \N__50044\,
            I => \N__49949\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__50041\,
            I => \N__49949\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__50032\,
            I => \N__49949\
        );

    \I__10326\ : Span4Mux_v
    port map (
            O => \N__50029\,
            I => \N__49939\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__50026\,
            I => \N__49934\
        );

    \I__10324\ : Span12Mux_v
    port map (
            O => \N__50023\,
            I => \N__49934\
        );

    \I__10323\ : InMux
    port map (
            O => \N__50022\,
            I => \N__49925\
        );

    \I__10322\ : InMux
    port map (
            O => \N__50021\,
            I => \N__49925\
        );

    \I__10321\ : InMux
    port map (
            O => \N__50020\,
            I => \N__49925\
        );

    \I__10320\ : InMux
    port map (
            O => \N__50019\,
            I => \N__49925\
        );

    \I__10319\ : LocalMux
    port map (
            O => \N__50012\,
            I => \N__49922\
        );

    \I__10318\ : InMux
    port map (
            O => \N__50011\,
            I => \N__49911\
        );

    \I__10317\ : InMux
    port map (
            O => \N__50010\,
            I => \N__49911\
        );

    \I__10316\ : InMux
    port map (
            O => \N__50009\,
            I => \N__49911\
        );

    \I__10315\ : InMux
    port map (
            O => \N__50008\,
            I => \N__49911\
        );

    \I__10314\ : InMux
    port map (
            O => \N__50007\,
            I => \N__49911\
        );

    \I__10313\ : InMux
    port map (
            O => \N__50006\,
            I => \N__49902\
        );

    \I__10312\ : InMux
    port map (
            O => \N__50005\,
            I => \N__49902\
        );

    \I__10311\ : InMux
    port map (
            O => \N__50004\,
            I => \N__49902\
        );

    \I__10310\ : InMux
    port map (
            O => \N__50003\,
            I => \N__49902\
        );

    \I__10309\ : Span4Mux_v
    port map (
            O => \N__50000\,
            I => \N__49893\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__49991\,
            I => \N__49893\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__49986\,
            I => \N__49893\
        );

    \I__10306\ : Span4Mux_h
    port map (
            O => \N__49979\,
            I => \N__49893\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__49974\,
            I => \N__49888\
        );

    \I__10304\ : Span4Mux_v
    port map (
            O => \N__49969\,
            I => \N__49888\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__49956\,
            I => \N__49883\
        );

    \I__10302\ : Span4Mux_h
    port map (
            O => \N__49949\,
            I => \N__49883\
        );

    \I__10301\ : InMux
    port map (
            O => \N__49948\,
            I => \N__49880\
        );

    \I__10300\ : InMux
    port map (
            O => \N__49947\,
            I => \N__49867\
        );

    \I__10299\ : InMux
    port map (
            O => \N__49946\,
            I => \N__49867\
        );

    \I__10298\ : InMux
    port map (
            O => \N__49945\,
            I => \N__49867\
        );

    \I__10297\ : InMux
    port map (
            O => \N__49944\,
            I => \N__49867\
        );

    \I__10296\ : InMux
    port map (
            O => \N__49943\,
            I => \N__49867\
        );

    \I__10295\ : InMux
    port map (
            O => \N__49942\,
            I => \N__49867\
        );

    \I__10294\ : Odrv4
    port map (
            O => \N__49939\,
            I => \busState_1\
        );

    \I__10293\ : Odrv12
    port map (
            O => \N__49934\,
            I => \busState_1\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__49925\,
            I => \busState_1\
        );

    \I__10291\ : Odrv12
    port map (
            O => \N__49922\,
            I => \busState_1\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__49911\,
            I => \busState_1\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__49902\,
            I => \busState_1\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__49893\,
            I => \busState_1\
        );

    \I__10287\ : Odrv4
    port map (
            O => \N__49888\,
            I => \busState_1\
        );

    \I__10286\ : Odrv4
    port map (
            O => \N__49883\,
            I => \busState_1\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__49880\,
            I => \busState_1\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__49867\,
            I => \busState_1\
        );

    \I__10283\ : CascadeMux
    port map (
            O => \N__49844\,
            I => \N_208_cascade_\
        );

    \I__10282\ : CascadeMux
    port map (
            O => \N__49841\,
            I => \ALU.status_19_14_cascade_\
        );

    \I__10281\ : InMux
    port map (
            O => \N__49838\,
            I => \N__49835\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__49835\,
            I => \N_208\
        );

    \I__10279\ : InMux
    port map (
            O => \N__49832\,
            I => \N__49826\
        );

    \I__10278\ : InMux
    port map (
            O => \N__49831\,
            I => \N__49819\
        );

    \I__10277\ : InMux
    port map (
            O => \N__49830\,
            I => \N__49819\
        );

    \I__10276\ : InMux
    port map (
            O => \N__49829\,
            I => \N__49812\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__49826\,
            I => \N__49807\
        );

    \I__10274\ : InMux
    port map (
            O => \N__49825\,
            I => \N__49803\
        );

    \I__10273\ : CascadeMux
    port map (
            O => \N__49824\,
            I => \N__49799\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__49819\,
            I => \N__49794\
        );

    \I__10271\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49790\
        );

    \I__10270\ : InMux
    port map (
            O => \N__49817\,
            I => \N__49787\
        );

    \I__10269\ : InMux
    port map (
            O => \N__49816\,
            I => \N__49780\
        );

    \I__10268\ : InMux
    port map (
            O => \N__49815\,
            I => \N__49780\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__49812\,
            I => \N__49777\
        );

    \I__10266\ : InMux
    port map (
            O => \N__49811\,
            I => \N__49774\
        );

    \I__10265\ : InMux
    port map (
            O => \N__49810\,
            I => \N__49771\
        );

    \I__10264\ : Span4Mux_v
    port map (
            O => \N__49807\,
            I => \N__49768\
        );

    \I__10263\ : InMux
    port map (
            O => \N__49806\,
            I => \N__49765\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__49803\,
            I => \N__49762\
        );

    \I__10261\ : InMux
    port map (
            O => \N__49802\,
            I => \N__49759\
        );

    \I__10260\ : InMux
    port map (
            O => \N__49799\,
            I => \N__49755\
        );

    \I__10259\ : InMux
    port map (
            O => \N__49798\,
            I => \N__49752\
        );

    \I__10258\ : InMux
    port map (
            O => \N__49797\,
            I => \N__49749\
        );

    \I__10257\ : Span4Mux_h
    port map (
            O => \N__49794\,
            I => \N__49746\
        );

    \I__10256\ : InMux
    port map (
            O => \N__49793\,
            I => \N__49743\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__49790\,
            I => \N__49739\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__49787\,
            I => \N__49736\
        );

    \I__10253\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49733\
        );

    \I__10252\ : InMux
    port map (
            O => \N__49785\,
            I => \N__49730\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__49780\,
            I => \N__49727\
        );

    \I__10250\ : Span4Mux_v
    port map (
            O => \N__49777\,
            I => \N__49724\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__49774\,
            I => \N__49719\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__49771\,
            I => \N__49719\
        );

    \I__10247\ : Span4Mux_h
    port map (
            O => \N__49768\,
            I => \N__49712\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__49765\,
            I => \N__49712\
        );

    \I__10245\ : Span4Mux_v
    port map (
            O => \N__49762\,
            I => \N__49712\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__49759\,
            I => \N__49706\
        );

    \I__10243\ : InMux
    port map (
            O => \N__49758\,
            I => \N__49703\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__49755\,
            I => \N__49700\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__49752\,
            I => \N__49697\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__49749\,
            I => \N__49690\
        );

    \I__10239\ : Span4Mux_h
    port map (
            O => \N__49746\,
            I => \N__49690\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__49743\,
            I => \N__49690\
        );

    \I__10237\ : InMux
    port map (
            O => \N__49742\,
            I => \N__49687\
        );

    \I__10236\ : Span12Mux_v
    port map (
            O => \N__49739\,
            I => \N__49684\
        );

    \I__10235\ : Span12Mux_h
    port map (
            O => \N__49736\,
            I => \N__49681\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__49733\,
            I => \N__49678\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__49730\,
            I => \N__49675\
        );

    \I__10232\ : Span4Mux_v
    port map (
            O => \N__49727\,
            I => \N__49666\
        );

    \I__10231\ : Span4Mux_v
    port map (
            O => \N__49724\,
            I => \N__49666\
        );

    \I__10230\ : Span4Mux_v
    port map (
            O => \N__49719\,
            I => \N__49666\
        );

    \I__10229\ : Span4Mux_h
    port map (
            O => \N__49712\,
            I => \N__49666\
        );

    \I__10228\ : InMux
    port map (
            O => \N__49711\,
            I => \N__49659\
        );

    \I__10227\ : InMux
    port map (
            O => \N__49710\,
            I => \N__49659\
        );

    \I__10226\ : InMux
    port map (
            O => \N__49709\,
            I => \N__49659\
        );

    \I__10225\ : Span4Mux_h
    port map (
            O => \N__49706\,
            I => \N__49652\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__49703\,
            I => \N__49652\
        );

    \I__10223\ : Span4Mux_h
    port map (
            O => \N__49700\,
            I => \N__49652\
        );

    \I__10222\ : Span4Mux_h
    port map (
            O => \N__49697\,
            I => \N__49647\
        );

    \I__10221\ : Span4Mux_h
    port map (
            O => \N__49690\,
            I => \N__49647\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__49687\,
            I => \busState_0\
        );

    \I__10219\ : Odrv12
    port map (
            O => \N__49684\,
            I => \busState_0\
        );

    \I__10218\ : Odrv12
    port map (
            O => \N__49681\,
            I => \busState_0\
        );

    \I__10217\ : Odrv4
    port map (
            O => \N__49678\,
            I => \busState_0\
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__49675\,
            I => \busState_0\
        );

    \I__10215\ : Odrv4
    port map (
            O => \N__49666\,
            I => \busState_0\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__49659\,
            I => \busState_0\
        );

    \I__10213\ : Odrv4
    port map (
            O => \N__49652\,
            I => \busState_0\
        );

    \I__10212\ : Odrv4
    port map (
            O => \N__49647\,
            I => \busState_0\
        );

    \I__10211\ : CascadeMux
    port map (
            O => \N__49628\,
            I => \N__49625\
        );

    \I__10210\ : InMux
    port map (
            O => \N__49625\,
            I => \N__49622\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__49622\,
            I => \N__49619\
        );

    \I__10208\ : Span4Mux_v
    port map (
            O => \N__49619\,
            I => \N__49616\
        );

    \I__10207\ : Span4Mux_v
    port map (
            O => \N__49616\,
            I => \N__49613\
        );

    \I__10206\ : Span4Mux_h
    port map (
            O => \N__49613\,
            I => \N__49610\
        );

    \I__10205\ : Odrv4
    port map (
            O => \N__49610\,
            I => \CONTROL.bus_7_ns_1_15\
        );

    \I__10204\ : InMux
    port map (
            O => \N__49607\,
            I => \N__49601\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__49606\,
            I => \N__49597\
        );

    \I__10202\ : InMux
    port map (
            O => \N__49605\,
            I => \N__49589\
        );

    \I__10201\ : InMux
    port map (
            O => \N__49604\,
            I => \N__49584\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__49601\,
            I => \N__49569\
        );

    \I__10199\ : InMux
    port map (
            O => \N__49600\,
            I => \N__49564\
        );

    \I__10198\ : InMux
    port map (
            O => \N__49597\,
            I => \N__49564\
        );

    \I__10197\ : InMux
    port map (
            O => \N__49596\,
            I => \N__49554\
        );

    \I__10196\ : InMux
    port map (
            O => \N__49595\,
            I => \N__49554\
        );

    \I__10195\ : InMux
    port map (
            O => \N__49594\,
            I => \N__49554\
        );

    \I__10194\ : InMux
    port map (
            O => \N__49593\,
            I => \N__49547\
        );

    \I__10193\ : InMux
    port map (
            O => \N__49592\,
            I => \N__49547\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__49589\,
            I => \N__49541\
        );

    \I__10191\ : InMux
    port map (
            O => \N__49588\,
            I => \N__49538\
        );

    \I__10190\ : InMux
    port map (
            O => \N__49587\,
            I => \N__49535\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__49584\,
            I => \N__49529\
        );

    \I__10188\ : InMux
    port map (
            O => \N__49583\,
            I => \N__49525\
        );

    \I__10187\ : CascadeMux
    port map (
            O => \N__49582\,
            I => \N__49520\
        );

    \I__10186\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49516\
        );

    \I__10185\ : InMux
    port map (
            O => \N__49580\,
            I => \N__49513\
        );

    \I__10184\ : CascadeMux
    port map (
            O => \N__49579\,
            I => \N__49509\
        );

    \I__10183\ : CascadeMux
    port map (
            O => \N__49578\,
            I => \N__49506\
        );

    \I__10182\ : InMux
    port map (
            O => \N__49577\,
            I => \N__49502\
        );

    \I__10181\ : InMux
    port map (
            O => \N__49576\,
            I => \N__49496\
        );

    \I__10180\ : InMux
    port map (
            O => \N__49575\,
            I => \N__49496\
        );

    \I__10179\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49486\
        );

    \I__10178\ : InMux
    port map (
            O => \N__49573\,
            I => \N__49486\
        );

    \I__10177\ : InMux
    port map (
            O => \N__49572\,
            I => \N__49486\
        );

    \I__10176\ : Span4Mux_v
    port map (
            O => \N__49569\,
            I => \N__49481\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__49564\,
            I => \N__49481\
        );

    \I__10174\ : InMux
    port map (
            O => \N__49563\,
            I => \N__49478\
        );

    \I__10173\ : InMux
    port map (
            O => \N__49562\,
            I => \N__49475\
        );

    \I__10172\ : InMux
    port map (
            O => \N__49561\,
            I => \N__49472\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__49554\,
            I => \N__49469\
        );

    \I__10170\ : InMux
    port map (
            O => \N__49553\,
            I => \N__49464\
        );

    \I__10169\ : InMux
    port map (
            O => \N__49552\,
            I => \N__49464\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__49547\,
            I => \N__49461\
        );

    \I__10167\ : InMux
    port map (
            O => \N__49546\,
            I => \N__49456\
        );

    \I__10166\ : InMux
    port map (
            O => \N__49545\,
            I => \N__49456\
        );

    \I__10165\ : InMux
    port map (
            O => \N__49544\,
            I => \N__49453\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__49541\,
            I => \N__49450\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__49538\,
            I => \N__49445\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__49535\,
            I => \N__49445\
        );

    \I__10161\ : InMux
    port map (
            O => \N__49534\,
            I => \N__49438\
        );

    \I__10160\ : InMux
    port map (
            O => \N__49533\,
            I => \N__49438\
        );

    \I__10159\ : InMux
    port map (
            O => \N__49532\,
            I => \N__49438\
        );

    \I__10158\ : Span4Mux_h
    port map (
            O => \N__49529\,
            I => \N__49435\
        );

    \I__10157\ : CascadeMux
    port map (
            O => \N__49528\,
            I => \N__49432\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__49525\,
            I => \N__49428\
        );

    \I__10155\ : InMux
    port map (
            O => \N__49524\,
            I => \N__49423\
        );

    \I__10154\ : InMux
    port map (
            O => \N__49523\,
            I => \N__49423\
        );

    \I__10153\ : InMux
    port map (
            O => \N__49520\,
            I => \N__49418\
        );

    \I__10152\ : InMux
    port map (
            O => \N__49519\,
            I => \N__49418\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__49516\,
            I => \N__49413\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__49513\,
            I => \N__49413\
        );

    \I__10149\ : InMux
    port map (
            O => \N__49512\,
            I => \N__49408\
        );

    \I__10148\ : InMux
    port map (
            O => \N__49509\,
            I => \N__49408\
        );

    \I__10147\ : InMux
    port map (
            O => \N__49506\,
            I => \N__49405\
        );

    \I__10146\ : CascadeMux
    port map (
            O => \N__49505\,
            I => \N__49402\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__49502\,
            I => \N__49399\
        );

    \I__10144\ : InMux
    port map (
            O => \N__49501\,
            I => \N__49396\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__49496\,
            I => \N__49393\
        );

    \I__10142\ : InMux
    port map (
            O => \N__49495\,
            I => \N__49384\
        );

    \I__10141\ : InMux
    port map (
            O => \N__49494\,
            I => \N__49384\
        );

    \I__10140\ : InMux
    port map (
            O => \N__49493\,
            I => \N__49384\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__49486\,
            I => \N__49375\
        );

    \I__10138\ : Span4Mux_h
    port map (
            O => \N__49481\,
            I => \N__49375\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__49478\,
            I => \N__49375\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__49475\,
            I => \N__49375\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__49472\,
            I => \N__49370\
        );

    \I__10134\ : Span4Mux_v
    port map (
            O => \N__49469\,
            I => \N__49370\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__49464\,
            I => \N__49367\
        );

    \I__10132\ : Span4Mux_v
    port map (
            O => \N__49461\,
            I => \N__49364\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__49456\,
            I => \N__49361\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__49453\,
            I => \N__49354\
        );

    \I__10129\ : Span4Mux_v
    port map (
            O => \N__49450\,
            I => \N__49354\
        );

    \I__10128\ : Span4Mux_h
    port map (
            O => \N__49445\,
            I => \N__49354\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__49438\,
            I => \N__49351\
        );

    \I__10126\ : Span4Mux_v
    port map (
            O => \N__49435\,
            I => \N__49348\
        );

    \I__10125\ : InMux
    port map (
            O => \N__49432\,
            I => \N__49343\
        );

    \I__10124\ : InMux
    port map (
            O => \N__49431\,
            I => \N__49343\
        );

    \I__10123\ : Span4Mux_v
    port map (
            O => \N__49428\,
            I => \N__49334\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__49423\,
            I => \N__49334\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__49418\,
            I => \N__49331\
        );

    \I__10120\ : Span4Mux_h
    port map (
            O => \N__49413\,
            I => \N__49324\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__49408\,
            I => \N__49324\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__49405\,
            I => \N__49324\
        );

    \I__10117\ : InMux
    port map (
            O => \N__49402\,
            I => \N__49317\
        );

    \I__10116\ : Span4Mux_v
    port map (
            O => \N__49399\,
            I => \N__49312\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__49396\,
            I => \N__49312\
        );

    \I__10114\ : Span4Mux_v
    port map (
            O => \N__49393\,
            I => \N__49309\
        );

    \I__10113\ : InMux
    port map (
            O => \N__49392\,
            I => \N__49304\
        );

    \I__10112\ : InMux
    port map (
            O => \N__49391\,
            I => \N__49304\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__49384\,
            I => \N__49295\
        );

    \I__10110\ : Span4Mux_v
    port map (
            O => \N__49375\,
            I => \N__49295\
        );

    \I__10109\ : Span4Mux_h
    port map (
            O => \N__49370\,
            I => \N__49295\
        );

    \I__10108\ : Span4Mux_h
    port map (
            O => \N__49367\,
            I => \N__49295\
        );

    \I__10107\ : Span4Mux_h
    port map (
            O => \N__49364\,
            I => \N__49286\
        );

    \I__10106\ : Span4Mux_v
    port map (
            O => \N__49361\,
            I => \N__49286\
        );

    \I__10105\ : Span4Mux_v
    port map (
            O => \N__49354\,
            I => \N__49286\
        );

    \I__10104\ : Span4Mux_v
    port map (
            O => \N__49351\,
            I => \N__49286\
        );

    \I__10103\ : Span4Mux_v
    port map (
            O => \N__49348\,
            I => \N__49281\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__49343\,
            I => \N__49281\
        );

    \I__10101\ : InMux
    port map (
            O => \N__49342\,
            I => \N__49272\
        );

    \I__10100\ : InMux
    port map (
            O => \N__49341\,
            I => \N__49272\
        );

    \I__10099\ : InMux
    port map (
            O => \N__49340\,
            I => \N__49272\
        );

    \I__10098\ : InMux
    port map (
            O => \N__49339\,
            I => \N__49272\
        );

    \I__10097\ : Span4Mux_v
    port map (
            O => \N__49334\,
            I => \N__49269\
        );

    \I__10096\ : Span4Mux_v
    port map (
            O => \N__49331\,
            I => \N__49264\
        );

    \I__10095\ : Span4Mux_h
    port map (
            O => \N__49324\,
            I => \N__49264\
        );

    \I__10094\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49255\
        );

    \I__10093\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49255\
        );

    \I__10092\ : InMux
    port map (
            O => \N__49321\,
            I => \N__49255\
        );

    \I__10091\ : InMux
    port map (
            O => \N__49320\,
            I => \N__49255\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__49317\,
            I => \busState_2\
        );

    \I__10089\ : Odrv4
    port map (
            O => \N__49312\,
            I => \busState_2\
        );

    \I__10088\ : Odrv4
    port map (
            O => \N__49309\,
            I => \busState_2\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__49304\,
            I => \busState_2\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__49295\,
            I => \busState_2\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__49286\,
            I => \busState_2\
        );

    \I__10084\ : Odrv4
    port map (
            O => \N__49281\,
            I => \busState_2\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__49272\,
            I => \busState_2\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__49269\,
            I => \busState_2\
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__49264\,
            I => \busState_2\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__49255\,
            I => \busState_2\
        );

    \I__10079\ : IoInMux
    port map (
            O => \N__49232\,
            I => \N__49229\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__49229\,
            I => \N__49226\
        );

    \I__10077\ : IoSpan4Mux
    port map (
            O => \N__49226\,
            I => \N__49223\
        );

    \I__10076\ : Span4Mux_s3_h
    port map (
            O => \N__49223\,
            I => \N__49220\
        );

    \I__10075\ : Span4Mux_h
    port map (
            O => \N__49220\,
            I => \N__49216\
        );

    \I__10074\ : IoInMux
    port map (
            O => \N__49219\,
            I => \N__49213\
        );

    \I__10073\ : Span4Mux_h
    port map (
            O => \N__49216\,
            I => \N__49210\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__49213\,
            I => \N__49207\
        );

    \I__10071\ : Sp12to4
    port map (
            O => \N__49210\,
            I => \N__49204\
        );

    \I__10070\ : Span4Mux_s2_h
    port map (
            O => \N__49207\,
            I => \N__49201\
        );

    \I__10069\ : Span12Mux_h
    port map (
            O => \N__49204\,
            I => \N__49198\
        );

    \I__10068\ : Span4Mux_v
    port map (
            O => \N__49201\,
            I => \N__49195\
        );

    \I__10067\ : Span12Mux_v
    port map (
            O => \N__49198\,
            I => \N__49189\
        );

    \I__10066\ : Sp12to4
    port map (
            O => \N__49195\,
            I => \N__49189\
        );

    \I__10065\ : InMux
    port map (
            O => \N__49194\,
            I => \N__49186\
        );

    \I__10064\ : Odrv12
    port map (
            O => \N__49189\,
            I => bus_15
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__49186\,
            I => bus_15
        );

    \I__10062\ : CascadeMux
    port map (
            O => \N__49181\,
            I => \N__49178\
        );

    \I__10061\ : InMux
    port map (
            O => \N__49178\,
            I => \N__49174\
        );

    \I__10060\ : CascadeMux
    port map (
            O => \N__49177\,
            I => \N__49171\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__49174\,
            I => \N__49168\
        );

    \I__10058\ : InMux
    port map (
            O => \N__49171\,
            I => \N__49165\
        );

    \I__10057\ : Span4Mux_v
    port map (
            O => \N__49168\,
            I => \N__49159\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__49165\,
            I => \N__49159\
        );

    \I__10055\ : InMux
    port map (
            O => \N__49164\,
            I => \N__49156\
        );

    \I__10054\ : Span4Mux_h
    port map (
            O => \N__49159\,
            I => \N__49153\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__49156\,
            I => \N__49150\
        );

    \I__10052\ : Span4Mux_h
    port map (
            O => \N__49153\,
            I => \N__49147\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__49150\,
            I => \N__49144\
        );

    \I__10050\ : Span4Mux_v
    port map (
            O => \N__49147\,
            I => \N__49139\
        );

    \I__10049\ : Span4Mux_h
    port map (
            O => \N__49144\,
            I => \N__49139\
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__49139\,
            I => f_1
        );

    \I__10047\ : CascadeMux
    port map (
            O => \N__49136\,
            I => \N__49133\
        );

    \I__10046\ : InMux
    port map (
            O => \N__49133\,
            I => \N__49128\
        );

    \I__10045\ : CascadeMux
    port map (
            O => \N__49132\,
            I => \N__49125\
        );

    \I__10044\ : InMux
    port map (
            O => \N__49131\,
            I => \N__49122\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__49128\,
            I => \N__49119\
        );

    \I__10042\ : InMux
    port map (
            O => \N__49125\,
            I => \N__49116\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__49122\,
            I => \N__49113\
        );

    \I__10040\ : Span4Mux_v
    port map (
            O => \N__49119\,
            I => \N__49108\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__49116\,
            I => \N__49108\
        );

    \I__10038\ : Span4Mux_v
    port map (
            O => \N__49113\,
            I => \N__49105\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__49108\,
            I => \N__49102\
        );

    \I__10036\ : Span4Mux_v
    port map (
            O => \N__49105\,
            I => \N__49097\
        );

    \I__10035\ : Span4Mux_h
    port map (
            O => \N__49102\,
            I => \N__49097\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__49097\,
            I => \N__49094\
        );

    \I__10033\ : Odrv4
    port map (
            O => \N__49094\,
            I => f_0
        );

    \I__10032\ : CascadeMux
    port map (
            O => \N__49091\,
            I => \N__49088\
        );

    \I__10031\ : InMux
    port map (
            O => \N__49088\,
            I => \N__49085\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__49085\,
            I => \N__49082\
        );

    \I__10029\ : Span4Mux_v
    port map (
            O => \N__49082\,
            I => \N__49077\
        );

    \I__10028\ : CascadeMux
    port map (
            O => \N__49081\,
            I => \N__49074\
        );

    \I__10027\ : CascadeMux
    port map (
            O => \N__49080\,
            I => \N__49071\
        );

    \I__10026\ : Span4Mux_h
    port map (
            O => \N__49077\,
            I => \N__49068\
        );

    \I__10025\ : InMux
    port map (
            O => \N__49074\,
            I => \N__49063\
        );

    \I__10024\ : InMux
    port map (
            O => \N__49071\,
            I => \N__49063\
        );

    \I__10023\ : Span4Mux_h
    port map (
            O => \N__49068\,
            I => \N__49058\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__49063\,
            I => \N__49058\
        );

    \I__10021\ : Span4Mux_v
    port map (
            O => \N__49058\,
            I => \N__49055\
        );

    \I__10020\ : Odrv4
    port map (
            O => \N__49055\,
            I => f_7
        );

    \I__10019\ : InMux
    port map (
            O => \N__49052\,
            I => \N__49049\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__49049\,
            I => \N__49046\
        );

    \I__10017\ : Span4Mux_h
    port map (
            O => \N__49046\,
            I => \N__49041\
        );

    \I__10016\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49038\
        );

    \I__10015\ : CascadeMux
    port map (
            O => \N__49044\,
            I => \N__49035\
        );

    \I__10014\ : Span4Mux_v
    port map (
            O => \N__49041\,
            I => \N__49030\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__49038\,
            I => \N__49030\
        );

    \I__10012\ : InMux
    port map (
            O => \N__49035\,
            I => \N__49027\
        );

    \I__10011\ : Span4Mux_v
    port map (
            O => \N__49030\,
            I => \N__49024\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__49027\,
            I => \N__49021\
        );

    \I__10009\ : Span4Mux_h
    port map (
            O => \N__49024\,
            I => \N__49018\
        );

    \I__10008\ : Span4Mux_v
    port map (
            O => \N__49021\,
            I => \N__49015\
        );

    \I__10007\ : Sp12to4
    port map (
            O => \N__49018\,
            I => \N__49012\
        );

    \I__10006\ : Span4Mux_h
    port map (
            O => \N__49015\,
            I => \N__49009\
        );

    \I__10005\ : Span12Mux_h
    port map (
            O => \N__49012\,
            I => \N__49006\
        );

    \I__10004\ : Span4Mux_h
    port map (
            O => \N__49009\,
            I => \N__49003\
        );

    \I__10003\ : Odrv12
    port map (
            O => \N__49006\,
            I => f_8
        );

    \I__10002\ : Odrv4
    port map (
            O => \N__49003\,
            I => f_8
        );

    \I__10001\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48995\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__48995\,
            I => \N__48992\
        );

    \I__9999\ : Span4Mux_v
    port map (
            O => \N__48992\,
            I => \N__48988\
        );

    \I__9998\ : CascadeMux
    port map (
            O => \N__48991\,
            I => \N__48985\
        );

    \I__9997\ : Span4Mux_h
    port map (
            O => \N__48988\,
            I => \N__48982\
        );

    \I__9996\ : InMux
    port map (
            O => \N__48985\,
            I => \N__48978\
        );

    \I__9995\ : Span4Mux_h
    port map (
            O => \N__48982\,
            I => \N__48975\
        );

    \I__9994\ : InMux
    port map (
            O => \N__48981\,
            I => \N__48972\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__48978\,
            I => \N__48969\
        );

    \I__9992\ : Span4Mux_v
    port map (
            O => \N__48975\,
            I => \N__48966\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__48972\,
            I => \N__48963\
        );

    \I__9990\ : Span12Mux_h
    port map (
            O => \N__48969\,
            I => \N__48960\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__48966\,
            I => \N__48955\
        );

    \I__9988\ : Span4Mux_h
    port map (
            O => \N__48963\,
            I => \N__48955\
        );

    \I__9987\ : Odrv12
    port map (
            O => \N__48960\,
            I => f_9
        );

    \I__9986\ : Odrv4
    port map (
            O => \N__48955\,
            I => f_9
        );

    \I__9985\ : InMux
    port map (
            O => \N__48950\,
            I => \N__48947\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__48947\,
            I => \N__48944\
        );

    \I__9983\ : Span4Mux_v
    port map (
            O => \N__48944\,
            I => \N__48939\
        );

    \I__9982\ : InMux
    port map (
            O => \N__48943\,
            I => \N__48936\
        );

    \I__9981\ : InMux
    port map (
            O => \N__48942\,
            I => \N__48933\
        );

    \I__9980\ : Span4Mux_h
    port map (
            O => \N__48939\,
            I => \N__48928\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__48936\,
            I => \N__48928\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__48933\,
            I => \N__48925\
        );

    \I__9977\ : Span4Mux_v
    port map (
            O => \N__48928\,
            I => \N__48920\
        );

    \I__9976\ : Span4Mux_h
    port map (
            O => \N__48925\,
            I => \N__48920\
        );

    \I__9975\ : Span4Mux_h
    port map (
            O => \N__48920\,
            I => \N__48917\
        );

    \I__9974\ : Odrv4
    port map (
            O => \N__48917\,
            I => g_1
        );

    \I__9973\ : CascadeMux
    port map (
            O => \N__48914\,
            I => \N__48911\
        );

    \I__9972\ : InMux
    port map (
            O => \N__48911\,
            I => \N__48908\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__48908\,
            I => \N__48905\
        );

    \I__9970\ : Span4Mux_v
    port map (
            O => \N__48905\,
            I => \N__48902\
        );

    \I__9969\ : Span4Mux_h
    port map (
            O => \N__48902\,
            I => \N__48897\
        );

    \I__9968\ : InMux
    port map (
            O => \N__48901\,
            I => \N__48894\
        );

    \I__9967\ : InMux
    port map (
            O => \N__48900\,
            I => \N__48891\
        );

    \I__9966\ : Span4Mux_h
    port map (
            O => \N__48897\,
            I => \N__48886\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__48894\,
            I => \N__48886\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__48891\,
            I => \N__48883\
        );

    \I__9963\ : Span4Mux_v
    port map (
            O => \N__48886\,
            I => \N__48878\
        );

    \I__9962\ : Span4Mux_h
    port map (
            O => \N__48883\,
            I => \N__48878\
        );

    \I__9961\ : Span4Mux_h
    port map (
            O => \N__48878\,
            I => \N__48875\
        );

    \I__9960\ : Odrv4
    port map (
            O => \N__48875\,
            I => g_0
        );

    \I__9959\ : InMux
    port map (
            O => \N__48872\,
            I => \N__48868\
        );

    \I__9958\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48864\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__48868\,
            I => \N__48861\
        );

    \I__9956\ : CascadeMux
    port map (
            O => \N__48867\,
            I => \N__48858\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__48864\,
            I => \N__48855\
        );

    \I__9954\ : Span12Mux_v
    port map (
            O => \N__48861\,
            I => \N__48852\
        );

    \I__9953\ : InMux
    port map (
            O => \N__48858\,
            I => \N__48849\
        );

    \I__9952\ : Span4Mux_v
    port map (
            O => \N__48855\,
            I => \N__48846\
        );

    \I__9951\ : Span12Mux_h
    port map (
            O => \N__48852\,
            I => \N__48843\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__48849\,
            I => \N__48838\
        );

    \I__9949\ : Sp12to4
    port map (
            O => \N__48846\,
            I => \N__48838\
        );

    \I__9948\ : Odrv12
    port map (
            O => \N__48843\,
            I => g_7
        );

    \I__9947\ : Odrv12
    port map (
            O => \N__48838\,
            I => g_7
        );

    \I__9946\ : InMux
    port map (
            O => \N__48833\,
            I => \N__48829\
        );

    \I__9945\ : InMux
    port map (
            O => \N__48832\,
            I => \N__48826\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__48829\,
            I => \N__48823\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__48826\,
            I => \N__48820\
        );

    \I__9942\ : Span4Mux_v
    port map (
            O => \N__48823\,
            I => \N__48817\
        );

    \I__9941\ : Span12Mux_h
    port map (
            O => \N__48820\,
            I => \N__48814\
        );

    \I__9940\ : Sp12to4
    port map (
            O => \N__48817\,
            I => \N__48811\
        );

    \I__9939\ : Odrv12
    port map (
            O => \N__48814\,
            I => \ALU.bZ0Z_9\
        );

    \I__9938\ : Odrv12
    port map (
            O => \N__48811\,
            I => \ALU.bZ0Z_9\
        );

    \I__9937\ : CascadeMux
    port map (
            O => \N__48806\,
            I => \N__48803\
        );

    \I__9936\ : InMux
    port map (
            O => \N__48803\,
            I => \N__48800\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__48800\,
            I => \N__48797\
        );

    \I__9934\ : Span4Mux_v
    port map (
            O => \N__48797\,
            I => \N__48794\
        );

    \I__9933\ : Span4Mux_h
    port map (
            O => \N__48794\,
            I => \N__48791\
        );

    \I__9932\ : Span4Mux_h
    port map (
            O => \N__48791\,
            I => \N__48787\
        );

    \I__9931\ : InMux
    port map (
            O => \N__48790\,
            I => \N__48784\
        );

    \I__9930\ : Odrv4
    port map (
            O => \N__48787\,
            I => \ALU.mult_9_8\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__48784\,
            I => \ALU.mult_9_8\
        );

    \I__9928\ : InMux
    port map (
            O => \N__48779\,
            I => \N__48776\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__48776\,
            I => \N__48773\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__48773\,
            I => \N__48769\
        );

    \I__9925\ : CascadeMux
    port map (
            O => \N__48772\,
            I => \N__48766\
        );

    \I__9924\ : Span4Mux_h
    port map (
            O => \N__48769\,
            I => \N__48763\
        );

    \I__9923\ : InMux
    port map (
            O => \N__48766\,
            I => \N__48760\
        );

    \I__9922\ : Odrv4
    port map (
            O => \N__48763\,
            I => \ALU.mult_25_8\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__48760\,
            I => \ALU.mult_25_8\
        );

    \I__9920\ : CascadeMux
    port map (
            O => \N__48755\,
            I => \ALU.mult_495_c_RNIKOB51JZ0_cascade_\
        );

    \I__9919\ : InMux
    port map (
            O => \N__48752\,
            I => \N__48749\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__48749\,
            I => \N__48746\
        );

    \I__9917\ : Span4Mux_v
    port map (
            O => \N__48746\,
            I => \N__48742\
        );

    \I__9916\ : InMux
    port map (
            O => \N__48745\,
            I => \N__48739\
        );

    \I__9915\ : Span4Mux_h
    port map (
            O => \N__48742\,
            I => \N__48736\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__48739\,
            I => \N__48733\
        );

    \I__9913\ : Span4Mux_h
    port map (
            O => \N__48736\,
            I => \N__48730\
        );

    \I__9912\ : Span12Mux_h
    port map (
            O => \N__48733\,
            I => \N__48727\
        );

    \I__9911\ : Span4Mux_v
    port map (
            O => \N__48730\,
            I => \N__48724\
        );

    \I__9910\ : Odrv12
    port map (
            O => \N__48727\,
            I => \ALU.aZ0Z_8\
        );

    \I__9909\ : Odrv4
    port map (
            O => \N__48724\,
            I => \ALU.aZ0Z_8\
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__48719\,
            I => \N__48716\
        );

    \I__9907\ : InMux
    port map (
            O => \N__48716\,
            I => \N__48713\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__48713\,
            I => \ALU.lshift_15_ns_1_8\
        );

    \I__9905\ : InMux
    port map (
            O => \N__48710\,
            I => \N__48706\
        );

    \I__9904\ : InMux
    port map (
            O => \N__48709\,
            I => \N__48703\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__48706\,
            I => \N__48700\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__48703\,
            I => \N__48697\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__48700\,
            I => \N__48694\
        );

    \I__9900\ : Span4Mux_v
    port map (
            O => \N__48697\,
            I => \N__48691\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__48694\,
            I => \N__48688\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__48691\,
            I => \N__48685\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__48688\,
            I => \N__48680\
        );

    \I__9896\ : Span4Mux_h
    port map (
            O => \N__48685\,
            I => \N__48680\
        );

    \I__9895\ : Odrv4
    port map (
            O => \N__48680\,
            I => \ALU.N_610\
        );

    \I__9894\ : InMux
    port map (
            O => \N__48677\,
            I => \N__48674\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__48674\,
            I => \N__48669\
        );

    \I__9892\ : InMux
    port map (
            O => \N__48673\,
            I => \N__48666\
        );

    \I__9891\ : InMux
    port map (
            O => \N__48672\,
            I => \N__48663\
        );

    \I__9890\ : Span4Mux_v
    port map (
            O => \N__48669\,
            I => \N__48660\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__48666\,
            I => \N__48657\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__48663\,
            I => \N__48654\
        );

    \I__9887\ : Span4Mux_h
    port map (
            O => \N__48660\,
            I => \N__48651\
        );

    \I__9886\ : Span4Mux_h
    port map (
            O => \N__48657\,
            I => \N__48648\
        );

    \I__9885\ : Span4Mux_v
    port map (
            O => \N__48654\,
            I => \N__48645\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__48651\,
            I => \N__48640\
        );

    \I__9883\ : Span4Mux_v
    port map (
            O => \N__48648\,
            I => \N__48640\
        );

    \I__9882\ : Span4Mux_h
    port map (
            O => \N__48645\,
            I => \N__48637\
        );

    \I__9881\ : Sp12to4
    port map (
            O => \N__48640\,
            I => \N__48634\
        );

    \I__9880\ : Span4Mux_h
    port map (
            O => \N__48637\,
            I => \N__48631\
        );

    \I__9879\ : Odrv12
    port map (
            O => \N__48634\,
            I => \ALU.N_608\
        );

    \I__9878\ : Odrv4
    port map (
            O => \N__48631\,
            I => \ALU.N_608\
        );

    \I__9877\ : InMux
    port map (
            O => \N__48626\,
            I => \N__48623\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__48623\,
            I => \ALU.N_640\
        );

    \I__9875\ : CascadeMux
    port map (
            O => \N__48620\,
            I => \ALU.addsub_cry_7_c_RNIDLTNZ0Z71_cascade_\
        );

    \I__9874\ : InMux
    port map (
            O => \N__48617\,
            I => \N__48614\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__48614\,
            I => \ALU.lshift_8\
        );

    \I__9872\ : InMux
    port map (
            O => \N__48611\,
            I => \N__48607\
        );

    \I__9871\ : InMux
    port map (
            O => \N__48610\,
            I => \N__48604\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__48607\,
            I => \N__48599\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__48604\,
            I => \N__48599\
        );

    \I__9868\ : Odrv4
    port map (
            O => \N__48599\,
            I => \ALU.N_636\
        );

    \I__9867\ : CascadeMux
    port map (
            O => \N__48596\,
            I => \N__48592\
        );

    \I__9866\ : CascadeMux
    port map (
            O => \N__48595\,
            I => \N__48589\
        );

    \I__9865\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48584\
        );

    \I__9864\ : InMux
    port map (
            O => \N__48589\,
            I => \N__48584\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__48584\,
            I => \N__48580\
        );

    \I__9862\ : InMux
    port map (
            O => \N__48583\,
            I => \N__48577\
        );

    \I__9861\ : Span4Mux_v
    port map (
            O => \N__48580\,
            I => \N__48574\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__48577\,
            I => \N__48571\
        );

    \I__9859\ : Span4Mux_v
    port map (
            O => \N__48574\,
            I => \N__48568\
        );

    \I__9858\ : Span4Mux_v
    port map (
            O => \N__48571\,
            I => \N__48565\
        );

    \I__9857\ : Span4Mux_h
    port map (
            O => \N__48568\,
            I => \N__48562\
        );

    \I__9856\ : Span4Mux_v
    port map (
            O => \N__48565\,
            I => \N__48559\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__48562\,
            I => \ALU.N_794_1\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__48559\,
            I => \ALU.N_794_1\
        );

    \I__9853\ : InMux
    port map (
            O => \N__48554\,
            I => \N__48551\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__48551\,
            I => \N__48548\
        );

    \I__9851\ : Span4Mux_v
    port map (
            O => \N__48548\,
            I => \N__48545\
        );

    \I__9850\ : Span4Mux_h
    port map (
            O => \N__48545\,
            I => \N__48542\
        );

    \I__9849\ : Span4Mux_h
    port map (
            O => \N__48542\,
            I => \N__48539\
        );

    \I__9848\ : Span4Mux_h
    port map (
            O => \N__48539\,
            I => \N__48536\
        );

    \I__9847\ : Span4Mux_h
    port map (
            O => \N__48536\,
            I => \N__48532\
        );

    \I__9846\ : InMux
    port map (
            O => \N__48535\,
            I => \N__48529\
        );

    \I__9845\ : Span4Mux_h
    port map (
            O => \N__48532\,
            I => \N__48526\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__48529\,
            I => \N__48523\
        );

    \I__9843\ : Odrv4
    port map (
            O => \N__48526\,
            I => \ALU.N_809\
        );

    \I__9842\ : Odrv12
    port map (
            O => \N__48523\,
            I => \ALU.N_809\
        );

    \I__9841\ : InMux
    port map (
            O => \N__48518\,
            I => \N__48515\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__48515\,
            I => \N__48512\
        );

    \I__9839\ : Span4Mux_h
    port map (
            O => \N__48512\,
            I => \N__48509\
        );

    \I__9838\ : Odrv4
    port map (
            O => \N__48509\,
            I => \ALU.mult_12\
        );

    \I__9837\ : InMux
    port map (
            O => \N__48506\,
            I => \N__48503\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__48503\,
            I => \ALU.mult_555_c_RNI5VJUOIZ0\
        );

    \I__9835\ : InMux
    port map (
            O => \N__48500\,
            I => \N__48497\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__48497\,
            I => \N__48494\
        );

    \I__9833\ : Span4Mux_h
    port map (
            O => \N__48494\,
            I => \N__48491\
        );

    \I__9832\ : Odrv4
    port map (
            O => \N__48491\,
            I => \ALU.mult_546_c_RNIG1E6IZ0Z8\
        );

    \I__9831\ : CascadeMux
    port map (
            O => \N__48488\,
            I => \N__48484\
        );

    \I__9830\ : InMux
    port map (
            O => \N__48487\,
            I => \N__48481\
        );

    \I__9829\ : InMux
    port map (
            O => \N__48484\,
            I => \N__48478\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__48481\,
            I => \N__48475\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__48478\,
            I => \N__48472\
        );

    \I__9826\ : Span4Mux_v
    port map (
            O => \N__48475\,
            I => \N__48469\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__48472\,
            I => \N__48465\
        );

    \I__9824\ : Span4Mux_v
    port map (
            O => \N__48469\,
            I => \N__48460\
        );

    \I__9823\ : InMux
    port map (
            O => \N__48468\,
            I => \N__48457\
        );

    \I__9822\ : Span4Mux_h
    port map (
            O => \N__48465\,
            I => \N__48454\
        );

    \I__9821\ : CascadeMux
    port map (
            O => \N__48464\,
            I => \N__48450\
        );

    \I__9820\ : InMux
    port map (
            O => \N__48463\,
            I => \N__48447\
        );

    \I__9819\ : Span4Mux_h
    port map (
            O => \N__48460\,
            I => \N__48440\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__48457\,
            I => \N__48440\
        );

    \I__9817\ : Span4Mux_h
    port map (
            O => \N__48454\,
            I => \N__48440\
        );

    \I__9816\ : InMux
    port map (
            O => \N__48453\,
            I => \N__48435\
        );

    \I__9815\ : InMux
    port map (
            O => \N__48450\,
            I => \N__48435\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__48447\,
            I => \aluStatus_0\
        );

    \I__9813\ : Odrv4
    port map (
            O => \N__48440\,
            I => \aluStatus_0\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__48435\,
            I => \aluStatus_0\
        );

    \I__9811\ : CascadeMux
    port map (
            O => \N__48428\,
            I => \ALU.status_14_12_0_cascade_\
        );

    \I__9810\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48422\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__48422\,
            I => \N__48419\
        );

    \I__9808\ : Span4Mux_h
    port map (
            O => \N__48419\,
            I => \N__48416\
        );

    \I__9807\ : Span4Mux_v
    port map (
            O => \N__48416\,
            I => \N__48413\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__48413\,
            I => \ALU.status_RNO_1Z0Z_0\
        );

    \I__9805\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48406\
        );

    \I__9804\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48403\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__48406\,
            I => \N__48400\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__48403\,
            I => \N__48397\
        );

    \I__9801\ : Span4Mux_v
    port map (
            O => \N__48400\,
            I => \N__48392\
        );

    \I__9800\ : Span4Mux_v
    port map (
            O => \N__48397\,
            I => \N__48392\
        );

    \I__9799\ : Span4Mux_h
    port map (
            O => \N__48392\,
            I => \N__48389\
        );

    \I__9798\ : Span4Mux_h
    port map (
            O => \N__48389\,
            I => \N__48386\
        );

    \I__9797\ : Span4Mux_v
    port map (
            O => \N__48386\,
            I => \N__48383\
        );

    \I__9796\ : Odrv4
    port map (
            O => \N__48383\,
            I => \ALU.bZ0Z_1\
        );

    \I__9795\ : InMux
    port map (
            O => \N__48380\,
            I => \N__48377\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__48377\,
            I => \N__48373\
        );

    \I__9793\ : InMux
    port map (
            O => \N__48376\,
            I => \N__48370\
        );

    \I__9792\ : Span4Mux_v
    port map (
            O => \N__48373\,
            I => \N__48367\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__48370\,
            I => \N__48364\
        );

    \I__9790\ : Span4Mux_h
    port map (
            O => \N__48367\,
            I => \N__48361\
        );

    \I__9789\ : Span4Mux_h
    port map (
            O => \N__48364\,
            I => \N__48358\
        );

    \I__9788\ : Span4Mux_h
    port map (
            O => \N__48361\,
            I => \N__48353\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__48358\,
            I => \N__48353\
        );

    \I__9786\ : Span4Mux_v
    port map (
            O => \N__48353\,
            I => \N__48350\
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__48350\,
            I => \ALU.bZ0Z_0\
        );

    \I__9784\ : InMux
    port map (
            O => \N__48347\,
            I => \N__48343\
        );

    \I__9783\ : InMux
    port map (
            O => \N__48346\,
            I => \N__48340\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__48343\,
            I => \N__48335\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__48340\,
            I => \N__48335\
        );

    \I__9780\ : Span4Mux_h
    port map (
            O => \N__48335\,
            I => \N__48332\
        );

    \I__9779\ : Span4Mux_v
    port map (
            O => \N__48332\,
            I => \N__48329\
        );

    \I__9778\ : Odrv4
    port map (
            O => \N__48329\,
            I => \ALU.bZ0Z_7\
        );

    \I__9777\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48322\
        );

    \I__9776\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48319\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__48322\,
            I => \N__48316\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__48319\,
            I => \N__48313\
        );

    \I__9773\ : Span4Mux_h
    port map (
            O => \N__48316\,
            I => \N__48310\
        );

    \I__9772\ : Span4Mux_v
    port map (
            O => \N__48313\,
            I => \N__48307\
        );

    \I__9771\ : Span4Mux_h
    port map (
            O => \N__48310\,
            I => \N__48304\
        );

    \I__9770\ : Span4Mux_h
    port map (
            O => \N__48307\,
            I => \N__48301\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__48304\,
            I => \N__48298\
        );

    \I__9768\ : Span4Mux_h
    port map (
            O => \N__48301\,
            I => \N__48295\
        );

    \I__9767\ : Odrv4
    port map (
            O => \N__48298\,
            I => \ALU.bZ0Z_8\
        );

    \I__9766\ : Odrv4
    port map (
            O => \N__48295\,
            I => \ALU.bZ0Z_8\
        );

    \I__9765\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48287\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__48287\,
            I => \N__48284\
        );

    \I__9763\ : Span4Mux_v
    port map (
            O => \N__48284\,
            I => \N__48281\
        );

    \I__9762\ : Span4Mux_h
    port map (
            O => \N__48281\,
            I => \N__48278\
        );

    \I__9761\ : Span4Mux_h
    port map (
            O => \N__48278\,
            I => \N__48275\
        );

    \I__9760\ : Odrv4
    port map (
            O => \N__48275\,
            I => \ALU.d_RNILTVJG3Z0Z_3\
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__48272\,
            I => \ALU.mult_555_c_RNIJF56AMZ0_cascade_\
        );

    \I__9758\ : InMux
    port map (
            O => \N__48269\,
            I => \N__48266\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__48266\,
            I => \N__48262\
        );

    \I__9756\ : InMux
    port map (
            O => \N__48265\,
            I => \N__48259\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__48262\,
            I => \N__48256\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__48259\,
            I => \N__48253\
        );

    \I__9753\ : Span4Mux_h
    port map (
            O => \N__48256\,
            I => \N__48250\
        );

    \I__9752\ : Span4Mux_v
    port map (
            O => \N__48253\,
            I => \N__48247\
        );

    \I__9751\ : Span4Mux_v
    port map (
            O => \N__48250\,
            I => \N__48242\
        );

    \I__9750\ : Span4Mux_h
    port map (
            O => \N__48247\,
            I => \N__48242\
        );

    \I__9749\ : Span4Mux_h
    port map (
            O => \N__48242\,
            I => \N__48239\
        );

    \I__9748\ : Odrv4
    port map (
            O => \N__48239\,
            I => \ALU.aZ0Z_12\
        );

    \I__9747\ : InMux
    port map (
            O => \N__48236\,
            I => \N__48233\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__48233\,
            I => \N__48229\
        );

    \I__9745\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48226\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__48229\,
            I => \N__48223\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__48226\,
            I => \N__48220\
        );

    \I__9742\ : Span4Mux_h
    port map (
            O => \N__48223\,
            I => \N__48217\
        );

    \I__9741\ : Odrv4
    port map (
            O => \N__48220\,
            I => \ALU.N_612\
        );

    \I__9740\ : Odrv4
    port map (
            O => \N__48217\,
            I => \ALU.N_612\
        );

    \I__9739\ : CascadeMux
    port map (
            O => \N__48212\,
            I => \N__48209\
        );

    \I__9738\ : InMux
    port map (
            O => \N__48209\,
            I => \N__48206\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__48206\,
            I => \N__48203\
        );

    \I__9736\ : Span4Mux_v
    port map (
            O => \N__48203\,
            I => \N__48200\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__48200\,
            I => \N__48197\
        );

    \I__9734\ : Odrv4
    port map (
            O => \N__48197\,
            I => \ALU.N_614\
        );

    \I__9733\ : CascadeMux
    port map (
            O => \N__48194\,
            I => \ALU.lshift_7_ns_1_12_cascade_\
        );

    \I__9732\ : CascadeMux
    port map (
            O => \N__48191\,
            I => \ALU.N_704_cascade_\
        );

    \I__9731\ : CascadeMux
    port map (
            O => \N__48188\,
            I => \N__48185\
        );

    \I__9730\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48182\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__48182\,
            I => \ALU.d_RNIGNBT49Z0Z_8\
        );

    \I__9728\ : CascadeMux
    port map (
            O => \N__48179\,
            I => \ALU.d_RNIGNBT49Z0Z_8_cascade_\
        );

    \I__9727\ : InMux
    port map (
            O => \N__48176\,
            I => \N__48171\
        );

    \I__9726\ : InMux
    port map (
            O => \N__48175\,
            I => \N__48166\
        );

    \I__9725\ : InMux
    port map (
            O => \N__48174\,
            I => \N__48166\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__48171\,
            I => \N__48163\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__48166\,
            I => \N__48158\
        );

    \I__9722\ : Span4Mux_h
    port map (
            O => \N__48163\,
            I => \N__48158\
        );

    \I__9721\ : Span4Mux_v
    port map (
            O => \N__48158\,
            I => \N__48155\
        );

    \I__9720\ : Span4Mux_h
    port map (
            O => \N__48155\,
            I => \N__48152\
        );

    \I__9719\ : Span4Mux_v
    port map (
            O => \N__48152\,
            I => \N__48149\
        );

    \I__9718\ : Odrv4
    port map (
            O => \N__48149\,
            I => \ALU.N_18_0\
        );

    \I__9717\ : CascadeMux
    port map (
            O => \N__48146\,
            I => \N__48143\
        );

    \I__9716\ : InMux
    port map (
            O => \N__48143\,
            I => \N__48138\
        );

    \I__9715\ : InMux
    port map (
            O => \N__48142\,
            I => \N__48135\
        );

    \I__9714\ : InMux
    port map (
            O => \N__48141\,
            I => \N__48132\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__48138\,
            I => \N__48129\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__48135\,
            I => \N__48126\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__48132\,
            I => \N__48123\
        );

    \I__9710\ : Span4Mux_v
    port map (
            O => \N__48129\,
            I => \N__48118\
        );

    \I__9709\ : Span4Mux_h
    port map (
            O => \N__48126\,
            I => \N__48118\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__48123\,
            I => \N__48115\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__48118\,
            I => \N__48112\
        );

    \I__9706\ : Span4Mux_v
    port map (
            O => \N__48115\,
            I => \N__48109\
        );

    \I__9705\ : Span4Mux_h
    port map (
            O => \N__48112\,
            I => \N__48106\
        );

    \I__9704\ : Span4Mux_h
    port map (
            O => \N__48109\,
            I => \N__48103\
        );

    \I__9703\ : Span4Mux_v
    port map (
            O => \N__48106\,
            I => \N__48100\
        );

    \I__9702\ : Sp12to4
    port map (
            O => \N__48103\,
            I => \N__48097\
        );

    \I__9701\ : Odrv4
    port map (
            O => \N__48100\,
            I => h_8
        );

    \I__9700\ : Odrv12
    port map (
            O => \N__48097\,
            I => h_8
        );

    \I__9699\ : CascadeMux
    port map (
            O => \N__48092\,
            I => \ALU.lshift_3_ns_1_13_cascade_\
        );

    \I__9698\ : CascadeMux
    port map (
            O => \N__48089\,
            I => \ALU.N_645_cascade_\
        );

    \I__9697\ : InMux
    port map (
            O => \N__48086\,
            I => \N__48083\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__48083\,
            I => \N__48079\
        );

    \I__9695\ : InMux
    port map (
            O => \N__48082\,
            I => \N__48076\
        );

    \I__9694\ : Span4Mux_v
    port map (
            O => \N__48079\,
            I => \N__48073\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__48076\,
            I => \N__48068\
        );

    \I__9692\ : Span4Mux_h
    port map (
            O => \N__48073\,
            I => \N__48068\
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__48068\,
            I => \ALU.N_806_1\
        );

    \I__9690\ : CascadeMux
    port map (
            O => \N__48065\,
            I => \ALU.a_15_m1_am_1_13_cascade_\
        );

    \I__9689\ : CascadeMux
    port map (
            O => \N__48062\,
            I => \ALU.N_611_cascade_\
        );

    \I__9688\ : InMux
    port map (
            O => \N__48059\,
            I => \N__48055\
        );

    \I__9687\ : InMux
    port map (
            O => \N__48058\,
            I => \N__48052\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__48055\,
            I => \N__48049\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__48052\,
            I => \N__48046\
        );

    \I__9684\ : Span4Mux_h
    port map (
            O => \N__48049\,
            I => \N__48043\
        );

    \I__9683\ : Span12Mux_h
    port map (
            O => \N__48046\,
            I => \N__48040\
        );

    \I__9682\ : Span4Mux_h
    port map (
            O => \N__48043\,
            I => \N__48037\
        );

    \I__9681\ : Odrv12
    port map (
            O => \N__48040\,
            I => \ALU.N_609\
        );

    \I__9680\ : Odrv4
    port map (
            O => \N__48037\,
            I => \ALU.N_609\
        );

    \I__9679\ : InMux
    port map (
            O => \N__48032\,
            I => \N__48029\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__48029\,
            I => \ALU.N_641\
        );

    \I__9677\ : CascadeMux
    port map (
            O => \N__48026\,
            I => \ALU.N_641_cascade_\
        );

    \I__9676\ : InMux
    port map (
            O => \N__48023\,
            I => \N__48020\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__48020\,
            I => \N__48017\
        );

    \I__9674\ : Span4Mux_v
    port map (
            O => \N__48017\,
            I => \N__48012\
        );

    \I__9673\ : InMux
    port map (
            O => \N__48016\,
            I => \N__48007\
        );

    \I__9672\ : InMux
    port map (
            O => \N__48015\,
            I => \N__48007\
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__48012\,
            I => \ALU.N_637\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__48007\,
            I => \ALU.N_637\
        );

    \I__9669\ : InMux
    port map (
            O => \N__48002\,
            I => \N__47999\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__47999\,
            I => \N__47996\
        );

    \I__9667\ : Span12Mux_v
    port map (
            O => \N__47996\,
            I => \N__47993\
        );

    \I__9666\ : Odrv12
    port map (
            O => \N__47993\,
            I => \ALU.d_RNITG2137Z0Z_0\
        );

    \I__9665\ : CascadeMux
    port map (
            O => \N__47990\,
            I => \N__47987\
        );

    \I__9664\ : InMux
    port map (
            O => \N__47987\,
            I => \N__47982\
        );

    \I__9663\ : InMux
    port map (
            O => \N__47986\,
            I => \N__47979\
        );

    \I__9662\ : InMux
    port map (
            O => \N__47985\,
            I => \N__47975\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__47982\,
            I => \N__47972\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__47979\,
            I => \N__47969\
        );

    \I__9659\ : InMux
    port map (
            O => \N__47978\,
            I => \N__47966\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__47975\,
            I => \N__47963\
        );

    \I__9657\ : Span4Mux_h
    port map (
            O => \N__47972\,
            I => \N__47960\
        );

    \I__9656\ : Span4Mux_v
    port map (
            O => \N__47969\,
            I => \N__47957\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__47966\,
            I => \N__47954\
        );

    \I__9654\ : Span4Mux_h
    port map (
            O => \N__47963\,
            I => \N__47949\
        );

    \I__9653\ : Span4Mux_h
    port map (
            O => \N__47960\,
            I => \N__47949\
        );

    \I__9652\ : Odrv4
    port map (
            O => \N__47957\,
            I => \ALU.N_765\
        );

    \I__9651\ : Odrv12
    port map (
            O => \N__47954\,
            I => \ALU.N_765\
        );

    \I__9650\ : Odrv4
    port map (
            O => \N__47949\,
            I => \ALU.N_765\
        );

    \I__9649\ : InMux
    port map (
            O => \N__47942\,
            I => \N__47939\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__47939\,
            I => \ALU.a_15_m1_am_1_9\
        );

    \I__9647\ : InMux
    port map (
            O => \N__47936\,
            I => \N__47933\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__47933\,
            I => \N__47930\
        );

    \I__9645\ : Span4Mux_h
    port map (
            O => \N__47930\,
            I => \N__47927\
        );

    \I__9644\ : Span4Mux_h
    port map (
            O => \N__47927\,
            I => \N__47924\
        );

    \I__9643\ : Span4Mux_h
    port map (
            O => \N__47924\,
            I => \N__47921\
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__47921\,
            I => \ALU.a_15_m3_d_d_0_ns_1_3\
        );

    \I__9641\ : CascadeMux
    port map (
            O => \N__47918\,
            I => \PROM.ROMDATA.m451_bm_cascade_\
        );

    \I__9640\ : InMux
    port map (
            O => \N__47915\,
            I => \N__47912\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__47912\,
            I => \N__47909\
        );

    \I__9638\ : Odrv12
    port map (
            O => \N__47909\,
            I => \PROM.ROMDATA.m451_am\
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__47906\,
            I => \N__47903\
        );

    \I__9636\ : InMux
    port map (
            O => \N__47903\,
            I => \N__47900\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__47900\,
            I => \PROM.ROMDATA.m451_ns\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__47897\,
            I => \N__47894\
        );

    \I__9633\ : InMux
    port map (
            O => \N__47894\,
            I => \N__47891\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__47891\,
            I => \N__47888\
        );

    \I__9631\ : Odrv12
    port map (
            O => \N__47888\,
            I => \PROM.ROMDATA.m375_bm\
        );

    \I__9630\ : CascadeMux
    port map (
            O => \N__47885\,
            I => \N__47882\
        );

    \I__9629\ : InMux
    port map (
            O => \N__47882\,
            I => \N__47879\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__47879\,
            I => \N__47876\
        );

    \I__9627\ : Odrv4
    port map (
            O => \N__47876\,
            I => \PROM.ROMDATA.m376\
        );

    \I__9626\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47870\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__47870\,
            I => \PROM.ROMDATA.N_256_i\
        );

    \I__9624\ : InMux
    port map (
            O => \N__47867\,
            I => \N__47864\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__47864\,
            I => \N__47861\
        );

    \I__9622\ : Odrv4
    port map (
            O => \N__47861\,
            I => \PROM.ROMDATA.m389_bm\
        );

    \I__9621\ : CascadeMux
    port map (
            O => \N__47858\,
            I => \PROM.ROMDATA.m389_am_cascade_\
        );

    \I__9620\ : InMux
    port map (
            O => \N__47855\,
            I => \N__47852\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__47852\,
            I => \N__47849\
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__47849\,
            I => \PROM.ROMDATA.m389_ns\
        );

    \I__9617\ : InMux
    port map (
            O => \N__47846\,
            I => \N__47843\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__47843\,
            I => \N__47840\
        );

    \I__9615\ : Span4Mux_v
    port map (
            O => \N__47840\,
            I => \N__47836\
        );

    \I__9614\ : InMux
    port map (
            O => \N__47839\,
            I => \N__47833\
        );

    \I__9613\ : Span4Mux_h
    port map (
            O => \N__47836\,
            I => \N__47830\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__47833\,
            I => \N__47827\
        );

    \I__9611\ : Span4Mux_h
    port map (
            O => \N__47830\,
            I => \N__47824\
        );

    \I__9610\ : Span4Mux_h
    port map (
            O => \N__47827\,
            I => \N__47821\
        );

    \I__9609\ : Odrv4
    port map (
            O => \N__47824\,
            I => \CONTROL.programCounter_1_6\
        );

    \I__9608\ : Odrv4
    port map (
            O => \N__47821\,
            I => \CONTROL.programCounter_1_6\
        );

    \I__9607\ : CascadeMux
    port map (
            O => \N__47816\,
            I => \N__47813\
        );

    \I__9606\ : InMux
    port map (
            O => \N__47813\,
            I => \N__47810\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__47810\,
            I => \N__47807\
        );

    \I__9604\ : Odrv4
    port map (
            O => \N__47807\,
            I => \CONTROL.programCounter_1_reto_6\
        );

    \I__9603\ : InMux
    port map (
            O => \N__47804\,
            I => \N__47801\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__47801\,
            I => \PROM.ROMDATA.m51\
        );

    \I__9601\ : InMux
    port map (
            O => \N__47798\,
            I => \N__47795\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__47795\,
            I => \N__47792\
        );

    \I__9599\ : Span4Mux_h
    port map (
            O => \N__47792\,
            I => \N__47789\
        );

    \I__9598\ : Odrv4
    port map (
            O => \N__47789\,
            I => \PROM.ROMDATA.m433_am\
        );

    \I__9597\ : CascadeMux
    port map (
            O => \N__47786\,
            I => \PROM.ROMDATA.m399_am_cascade_\
        );

    \I__9596\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47780\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__47780\,
            I => \N__47777\
        );

    \I__9594\ : Span12Mux_v
    port map (
            O => \N__47777\,
            I => \N__47774\
        );

    \I__9593\ : Odrv12
    port map (
            O => \N__47774\,
            I => \PROM.ROMDATA.m399_bm\
        );

    \I__9592\ : InMux
    port map (
            O => \N__47771\,
            I => \N__47768\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__47768\,
            I => \N__47765\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__47765\,
            I => \PROM.ROMDATA.m399_ns\
        );

    \I__9589\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47759\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47756\
        );

    \I__9587\ : Span4Mux_h
    port map (
            O => \N__47756\,
            I => \N__47753\
        );

    \I__9586\ : Span4Mux_h
    port map (
            O => \N__47753\,
            I => \N__47750\
        );

    \I__9585\ : Span4Mux_h
    port map (
            O => \N__47750\,
            I => \N__47747\
        );

    \I__9584\ : Odrv4
    port map (
            O => \N__47747\,
            I => \PROM.ROMDATA.m461_ns_1\
        );

    \I__9583\ : InMux
    port map (
            O => \N__47744\,
            I => \N__47741\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__47741\,
            I => \N__47738\
        );

    \I__9581\ : Span4Mux_v
    port map (
            O => \N__47738\,
            I => \N__47735\
        );

    \I__9580\ : Span4Mux_h
    port map (
            O => \N__47735\,
            I => \N__47732\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__47732\,
            I => \N__47729\
        );

    \I__9578\ : Odrv4
    port map (
            O => \N__47729\,
            I => \CONTROL.addrstack_4\
        );

    \I__9577\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47723\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__47723\,
            I => \N__47720\
        );

    \I__9575\ : Odrv12
    port map (
            O => \N__47720\,
            I => \PROM.ROMDATA.m22\
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__47717\,
            I => \PROM.ROMDATA.m215_ns_1_1_1_cascade_\
        );

    \I__9573\ : InMux
    port map (
            O => \N__47714\,
            I => \N__47711\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__47711\,
            I => \PROM.ROMDATA.m215_ns_1_1\
        );

    \I__9571\ : InMux
    port map (
            O => \N__47708\,
            I => \N__47705\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__47705\,
            I => \PROM.ROMDATA.m256\
        );

    \I__9569\ : InMux
    port map (
            O => \N__47702\,
            I => \N__47699\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__47699\,
            I => \N__47696\
        );

    \I__9567\ : Odrv12
    port map (
            O => \N__47696\,
            I => \PROM.ROMDATA.m38\
        );

    \I__9566\ : InMux
    port map (
            O => \N__47693\,
            I => \N__47690\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__47690\,
            I => \PROM.ROMDATA.m251\
        );

    \I__9564\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47684\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__47684\,
            I => \PROM.ROMDATA.m253\
        );

    \I__9562\ : CascadeMux
    port map (
            O => \N__47681\,
            I => \N__47677\
        );

    \I__9561\ : CascadeMux
    port map (
            O => \N__47680\,
            I => \N__47674\
        );

    \I__9560\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47669\
        );

    \I__9559\ : InMux
    port map (
            O => \N__47674\,
            I => \N__47669\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__47669\,
            I => \N__47666\
        );

    \I__9557\ : Span4Mux_v
    port map (
            O => \N__47666\,
            I => \N__47663\
        );

    \I__9556\ : Odrv4
    port map (
            O => \N__47663\,
            I => \N_419\
        );

    \I__9555\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47657\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__47657\,
            I => \N__47654\
        );

    \I__9553\ : Span4Mux_v
    port map (
            O => \N__47654\,
            I => \N__47651\
        );

    \I__9552\ : Span4Mux_h
    port map (
            O => \N__47651\,
            I => \N__47648\
        );

    \I__9551\ : Span4Mux_h
    port map (
            O => \N__47648\,
            I => \N__47645\
        );

    \I__9550\ : Span4Mux_h
    port map (
            O => \N__47645\,
            I => \N__47642\
        );

    \I__9549\ : Odrv4
    port map (
            O => \N__47642\,
            I => \CONTROL.addrstackZ0Z_1\
        );

    \I__9548\ : InMux
    port map (
            O => \N__47639\,
            I => \N__47636\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__47636\,
            I => \N__47632\
        );

    \I__9546\ : InMux
    port map (
            O => \N__47635\,
            I => \N__47629\
        );

    \I__9545\ : Odrv4
    port map (
            O => \N__47632\,
            I => \CONTROL.dout_reto_3\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__47629\,
            I => \CONTROL.dout_reto_3\
        );

    \I__9543\ : CascadeMux
    port map (
            O => \N__47624\,
            I => \CONTROL.programCounter_ret_1_RNILA8IZ0Z_3_cascade_\
        );

    \I__9542\ : InMux
    port map (
            O => \N__47621\,
            I => \N__47618\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__47618\,
            I => \CONTROL.programCounter_ret_19_RNIEO8JZ0Z_3\
        );

    \I__9540\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47612\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__47612\,
            I => \N__47608\
        );

    \I__9538\ : InMux
    port map (
            O => \N__47611\,
            I => \N__47605\
        );

    \I__9537\ : Odrv4
    port map (
            O => \N__47608\,
            I => \CONTROL.programCounter_1_reto_0\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__47605\,
            I => \CONTROL.programCounter_1_reto_0\
        );

    \I__9535\ : InMux
    port map (
            O => \N__47600\,
            I => \N__47597\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__47597\,
            I => \N__47594\
        );

    \I__9533\ : Span12Mux_v
    port map (
            O => \N__47594\,
            I => \N__47591\
        );

    \I__9532\ : Odrv12
    port map (
            O => \N__47591\,
            I => \CONTROL.addrstack_3\
        );

    \I__9531\ : InMux
    port map (
            O => \N__47588\,
            I => \N__47585\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__47585\,
            I => \PROM.ROMDATA.m30\
        );

    \I__9529\ : InMux
    port map (
            O => \N__47582\,
            I => \N__47579\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__47579\,
            I => \N__47576\
        );

    \I__9527\ : Span4Mux_h
    port map (
            O => \N__47576\,
            I => \N__47573\
        );

    \I__9526\ : Odrv4
    port map (
            O => \N__47573\,
            I => \PROM.ROMDATA.m35_1\
        );

    \I__9525\ : InMux
    port map (
            O => \N__47570\,
            I => \N__47567\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__47567\,
            I => \PROM.ROMDATA.m35\
        );

    \I__9523\ : InMux
    port map (
            O => \N__47564\,
            I => \N__47560\
        );

    \I__9522\ : InMux
    port map (
            O => \N__47563\,
            I => \N__47557\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__47560\,
            I => \CONTROL.programCounter_1_reto_2\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__47557\,
            I => \CONTROL.programCounter_1_reto_2\
        );

    \I__9519\ : InMux
    port map (
            O => \N__47552\,
            I => \N__47549\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__47549\,
            I => \N__47546\
        );

    \I__9517\ : Span4Mux_v
    port map (
            O => \N__47546\,
            I => \N__47543\
        );

    \I__9516\ : Odrv4
    port map (
            O => \N__47543\,
            I => \PROM.ROMDATA.m392_am\
        );

    \I__9515\ : CascadeMux
    port map (
            O => \N__47540\,
            I => \PROM.ROMDATA.m163_cascade_\
        );

    \I__9514\ : InMux
    port map (
            O => \N__47537\,
            I => \N__47534\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__47534\,
            I => \N__47531\
        );

    \I__9512\ : Odrv4
    port map (
            O => \N__47531\,
            I => \PROM.ROMDATA.m176_x\
        );

    \I__9511\ : CascadeMux
    port map (
            O => \N__47528\,
            I => \N__47525\
        );

    \I__9510\ : InMux
    port map (
            O => \N__47525\,
            I => \N__47518\
        );

    \I__9509\ : InMux
    port map (
            O => \N__47524\,
            I => \N__47518\
        );

    \I__9508\ : CascadeMux
    port map (
            O => \N__47523\,
            I => \N__47515\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__47518\,
            I => \N__47511\
        );

    \I__9506\ : InMux
    port map (
            O => \N__47515\,
            I => \N__47508\
        );

    \I__9505\ : InMux
    port map (
            O => \N__47514\,
            I => \N__47505\
        );

    \I__9504\ : Span4Mux_v
    port map (
            O => \N__47511\,
            I => \N__47502\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__47508\,
            I => \PROM.ROMDATA.N_543_mux_2\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__47505\,
            I => \PROM.ROMDATA.N_543_mux_2\
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__47502\,
            I => \PROM.ROMDATA.N_543_mux_2\
        );

    \I__9500\ : CascadeMux
    port map (
            O => \N__47495\,
            I => \N__47491\
        );

    \I__9499\ : InMux
    port map (
            O => \N__47494\,
            I => \N__47485\
        );

    \I__9498\ : InMux
    port map (
            O => \N__47491\,
            I => \N__47478\
        );

    \I__9497\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47478\
        );

    \I__9496\ : InMux
    port map (
            O => \N__47489\,
            I => \N__47478\
        );

    \I__9495\ : CascadeMux
    port map (
            O => \N__47488\,
            I => \N__47472\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__47485\,
            I => \N__47469\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__47478\,
            I => \N__47466\
        );

    \I__9492\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47463\
        );

    \I__9491\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47456\
        );

    \I__9490\ : InMux
    port map (
            O => \N__47475\,
            I => \N__47456\
        );

    \I__9489\ : InMux
    port map (
            O => \N__47472\,
            I => \N__47456\
        );

    \I__9488\ : Span4Mux_v
    port map (
            O => \N__47469\,
            I => \N__47453\
        );

    \I__9487\ : Sp12to4
    port map (
            O => \N__47466\,
            I => \N__47450\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__47463\,
            I => \N__47447\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__47456\,
            I => \N__47442\
        );

    \I__9484\ : Sp12to4
    port map (
            O => \N__47453\,
            I => \N__47442\
        );

    \I__9483\ : Span12Mux_v
    port map (
            O => \N__47450\,
            I => \N__47437\
        );

    \I__9482\ : Span12Mux_h
    port map (
            O => \N__47447\,
            I => \N__47437\
        );

    \I__9481\ : Span12Mux_h
    port map (
            O => \N__47442\,
            I => \N__47434\
        );

    \I__9480\ : Odrv12
    port map (
            O => \N__47437\,
            I => \PROM.ROMDATA.N_569_mux\
        );

    \I__9479\ : Odrv12
    port map (
            O => \N__47434\,
            I => \PROM.ROMDATA.N_569_mux\
        );

    \I__9478\ : CascadeMux
    port map (
            O => \N__47429\,
            I => \PROM.ROMDATA.m109_am_1_cascade_\
        );

    \I__9477\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47423\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__47423\,
            I => \N__47420\
        );

    \I__9475\ : Sp12to4
    port map (
            O => \N__47420\,
            I => \N__47417\
        );

    \I__9474\ : Span12Mux_v
    port map (
            O => \N__47417\,
            I => \N__47414\
        );

    \I__9473\ : Span12Mux_h
    port map (
            O => \N__47414\,
            I => \N__47411\
        );

    \I__9472\ : Odrv12
    port map (
            O => \N__47411\,
            I => \CONTROL.addrstack_0\
        );

    \I__9471\ : InMux
    port map (
            O => \N__47408\,
            I => \N__47404\
        );

    \I__9470\ : InMux
    port map (
            O => \N__47407\,
            I => \N__47400\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__47404\,
            I => \N__47397\
        );

    \I__9468\ : InMux
    port map (
            O => \N__47403\,
            I => \N__47394\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__47400\,
            I => \N__47391\
        );

    \I__9466\ : Sp12to4
    port map (
            O => \N__47397\,
            I => \N__47388\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__47394\,
            I => \N__47383\
        );

    \I__9464\ : Span4Mux_h
    port map (
            O => \N__47391\,
            I => \N__47383\
        );

    \I__9463\ : Span12Mux_v
    port map (
            O => \N__47388\,
            I => \N__47380\
        );

    \I__9462\ : Span4Mux_v
    port map (
            O => \N__47383\,
            I => \N__47377\
        );

    \I__9461\ : Odrv12
    port map (
            O => \N__47380\,
            I => \N_415\
        );

    \I__9460\ : Odrv4
    port map (
            O => \N__47377\,
            I => \N_415\
        );

    \I__9459\ : InMux
    port map (
            O => \N__47372\,
            I => \N__47369\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__47369\,
            I => \PROM.ROMDATA.m422_am\
        );

    \I__9457\ : CascadeMux
    port map (
            O => \N__47366\,
            I => \PROM.ROMDATA.m422_bm_cascade_\
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__47363\,
            I => \N__47360\
        );

    \I__9455\ : InMux
    port map (
            O => \N__47360\,
            I => \N__47357\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__47357\,
            I => \N__47354\
        );

    \I__9453\ : Span4Mux_h
    port map (
            O => \N__47354\,
            I => \N__47351\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__47351\,
            I => \N__47348\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__47348\,
            I => \PROM.ROMDATA.m381_bm\
        );

    \I__9450\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47342\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__47342\,
            I => \N__47339\
        );

    \I__9448\ : Span4Mux_v
    port map (
            O => \N__47339\,
            I => \N__47336\
        );

    \I__9447\ : Span4Mux_h
    port map (
            O => \N__47336\,
            I => \N__47333\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__47333\,
            I => \PROM.ROMDATA.m298_am\
        );

    \I__9445\ : InMux
    port map (
            O => \N__47330\,
            I => \N__47327\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__47327\,
            I => \N__47324\
        );

    \I__9443\ : Span4Mux_v
    port map (
            O => \N__47324\,
            I => \N__47321\
        );

    \I__9442\ : Span4Mux_h
    port map (
            O => \N__47321\,
            I => \N__47318\
        );

    \I__9441\ : Span4Mux_h
    port map (
            O => \N__47318\,
            I => \N__47315\
        );

    \I__9440\ : Odrv4
    port map (
            O => \N__47315\,
            I => \CONTROL.programCounter_1_axb_4\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__47312\,
            I => \PROM.ROMDATA.N_543_mux_2_cascade_\
        );

    \I__9438\ : InMux
    port map (
            O => \N__47309\,
            I => \N__47306\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__47306\,
            I => \N__47302\
        );

    \I__9436\ : InMux
    port map (
            O => \N__47305\,
            I => \N__47299\
        );

    \I__9435\ : Span4Mux_v
    port map (
            O => \N__47302\,
            I => \N__47296\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__47299\,
            I => \N__47293\
        );

    \I__9433\ : Span4Mux_h
    port map (
            O => \N__47296\,
            I => \N__47288\
        );

    \I__9432\ : Span4Mux_h
    port map (
            O => \N__47293\,
            I => \N__47288\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__47288\,
            I => \PROM.ROMDATA.N_559_mux\
        );

    \I__9430\ : InMux
    port map (
            O => \N__47285\,
            I => \N__47281\
        );

    \I__9429\ : InMux
    port map (
            O => \N__47284\,
            I => \N__47278\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__47281\,
            I => \N__47268\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__47278\,
            I => \N__47265\
        );

    \I__9426\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47260\
        );

    \I__9425\ : InMux
    port map (
            O => \N__47276\,
            I => \N__47260\
        );

    \I__9424\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47255\
        );

    \I__9423\ : InMux
    port map (
            O => \N__47274\,
            I => \N__47255\
        );

    \I__9422\ : InMux
    port map (
            O => \N__47273\,
            I => \N__47250\
        );

    \I__9421\ : InMux
    port map (
            O => \N__47272\,
            I => \N__47250\
        );

    \I__9420\ : CascadeMux
    port map (
            O => \N__47271\,
            I => \N__47247\
        );

    \I__9419\ : Span4Mux_h
    port map (
            O => \N__47268\,
            I => \N__47243\
        );

    \I__9418\ : Span4Mux_h
    port map (
            O => \N__47265\,
            I => \N__47240\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__47260\,
            I => \N__47237\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__47255\,
            I => \N__47232\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__47250\,
            I => \N__47232\
        );

    \I__9414\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47227\
        );

    \I__9413\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47227\
        );

    \I__9412\ : Odrv4
    port map (
            O => \N__47243\,
            I => \aluOperand1_2\
        );

    \I__9411\ : Odrv4
    port map (
            O => \N__47240\,
            I => \aluOperand1_2\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__47237\,
            I => \aluOperand1_2\
        );

    \I__9409\ : Odrv12
    port map (
            O => \N__47232\,
            I => \aluOperand1_2\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__47227\,
            I => \aluOperand1_2\
        );

    \I__9407\ : CascadeMux
    port map (
            O => \N__47216\,
            I => \ALU.dout_6_ns_1_14_cascade_\
        );

    \I__9406\ : InMux
    port map (
            O => \N__47213\,
            I => \N__47205\
        );

    \I__9405\ : InMux
    port map (
            O => \N__47212\,
            I => \N__47205\
        );

    \I__9404\ : InMux
    port map (
            O => \N__47211\,
            I => \N__47196\
        );

    \I__9403\ : InMux
    port map (
            O => \N__47210\,
            I => \N__47196\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__47205\,
            I => \N__47185\
        );

    \I__9401\ : InMux
    port map (
            O => \N__47204\,
            I => \N__47180\
        );

    \I__9400\ : InMux
    port map (
            O => \N__47203\,
            I => \N__47180\
        );

    \I__9399\ : InMux
    port map (
            O => \N__47202\,
            I => \N__47175\
        );

    \I__9398\ : InMux
    port map (
            O => \N__47201\,
            I => \N__47175\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__47196\,
            I => \N__47172\
        );

    \I__9396\ : InMux
    port map (
            O => \N__47195\,
            I => \N__47167\
        );

    \I__9395\ : InMux
    port map (
            O => \N__47194\,
            I => \N__47167\
        );

    \I__9394\ : InMux
    port map (
            O => \N__47193\,
            I => \N__47162\
        );

    \I__9393\ : InMux
    port map (
            O => \N__47192\,
            I => \N__47162\
        );

    \I__9392\ : InMux
    port map (
            O => \N__47191\,
            I => \N__47157\
        );

    \I__9391\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47157\
        );

    \I__9390\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47152\
        );

    \I__9389\ : InMux
    port map (
            O => \N__47188\,
            I => \N__47152\
        );

    \I__9388\ : Span4Mux_h
    port map (
            O => \N__47185\,
            I => \N__47149\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__47180\,
            I => \N__47146\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__47175\,
            I => \N__47139\
        );

    \I__9385\ : Span4Mux_h
    port map (
            O => \N__47172\,
            I => \N__47136\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__47167\,
            I => \N__47133\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__47162\,
            I => \N__47128\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__47157\,
            I => \N__47128\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__47152\,
            I => \N__47121\
        );

    \I__9380\ : Span4Mux_v
    port map (
            O => \N__47149\,
            I => \N__47121\
        );

    \I__9379\ : Span4Mux_h
    port map (
            O => \N__47146\,
            I => \N__47121\
        );

    \I__9378\ : InMux
    port map (
            O => \N__47145\,
            I => \N__47112\
        );

    \I__9377\ : InMux
    port map (
            O => \N__47144\,
            I => \N__47112\
        );

    \I__9376\ : InMux
    port map (
            O => \N__47143\,
            I => \N__47112\
        );

    \I__9375\ : InMux
    port map (
            O => \N__47142\,
            I => \N__47112\
        );

    \I__9374\ : Odrv4
    port map (
            O => \N__47139\,
            I => \aluOperand1_1\
        );

    \I__9373\ : Odrv4
    port map (
            O => \N__47136\,
            I => \aluOperand1_1\
        );

    \I__9372\ : Odrv4
    port map (
            O => \N__47133\,
            I => \aluOperand1_1\
        );

    \I__9371\ : Odrv12
    port map (
            O => \N__47128\,
            I => \aluOperand1_1\
        );

    \I__9370\ : Odrv4
    port map (
            O => \N__47121\,
            I => \aluOperand1_1\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__47112\,
            I => \aluOperand1_1\
        );

    \I__9368\ : InMux
    port map (
            O => \N__47099\,
            I => \N__47096\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__47096\,
            I => \ALU.N_1099\
        );

    \I__9366\ : CascadeMux
    port map (
            O => \N__47093\,
            I => \ALU.N_1147_cascade_\
        );

    \I__9365\ : InMux
    port map (
            O => \N__47090\,
            I => \N__47087\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__47087\,
            I => \N__47084\
        );

    \I__9363\ : Span4Mux_v
    port map (
            O => \N__47084\,
            I => \N__47081\
        );

    \I__9362\ : Sp12to4
    port map (
            O => \N__47081\,
            I => \N__47078\
        );

    \I__9361\ : Odrv12
    port map (
            O => \N__47078\,
            I => \DROM_ROMDATA_dintern_14ro\
        );

    \I__9360\ : CascadeMux
    port map (
            O => \N__47075\,
            I => \aluOut_14_cascade_\
        );

    \I__9359\ : InMux
    port map (
            O => \N__47072\,
            I => \N__47069\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__47069\,
            I => \N__47066\
        );

    \I__9357\ : Span4Mux_h
    port map (
            O => \N__47066\,
            I => \N__47063\
        );

    \I__9356\ : Span4Mux_h
    port map (
            O => \N__47063\,
            I => \N__47059\
        );

    \I__9355\ : InMux
    port map (
            O => \N__47062\,
            I => \N__47056\
        );

    \I__9354\ : Odrv4
    port map (
            O => \N__47059\,
            I => \N_207\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__47056\,
            I => \N_207\
        );

    \I__9352\ : InMux
    port map (
            O => \N__47051\,
            I => \N__47047\
        );

    \I__9351\ : InMux
    port map (
            O => \N__47050\,
            I => \N__47044\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__47047\,
            I => \N__47040\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__47044\,
            I => \N__47037\
        );

    \I__9348\ : InMux
    port map (
            O => \N__47043\,
            I => \N__47034\
        );

    \I__9347\ : Span4Mux_h
    port map (
            O => \N__47040\,
            I => \N__47030\
        );

    \I__9346\ : Span4Mux_h
    port map (
            O => \N__47037\,
            I => \N__47025\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__47034\,
            I => \N__47025\
        );

    \I__9344\ : InMux
    port map (
            O => \N__47033\,
            I => \N__47022\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__47030\,
            I => \CONTROL.un1_busState114_2_0_o2_0_0\
        );

    \I__9342\ : Odrv4
    port map (
            O => \N__47025\,
            I => \CONTROL.un1_busState114_2_0_o2_0_0\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__47022\,
            I => \CONTROL.un1_busState114_2_0_o2_0_0\
        );

    \I__9340\ : InMux
    port map (
            O => \N__47015\,
            I => \N__47012\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__47012\,
            I => \N__47006\
        );

    \I__9338\ : InMux
    port map (
            O => \N__47011\,
            I => \N__47003\
        );

    \I__9337\ : InMux
    port map (
            O => \N__47010\,
            I => \N__46997\
        );

    \I__9336\ : InMux
    port map (
            O => \N__47009\,
            I => \N__46997\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__47006\,
            I => \N__46994\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__47003\,
            I => \N__46991\
        );

    \I__9333\ : InMux
    port map (
            O => \N__47002\,
            I => \N__46988\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__46997\,
            I => \N__46985\
        );

    \I__9331\ : Span4Mux_v
    port map (
            O => \N__46994\,
            I => \N__46981\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__46991\,
            I => \N__46974\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__46988\,
            I => \N__46974\
        );

    \I__9328\ : Span4Mux_v
    port map (
            O => \N__46985\,
            I => \N__46974\
        );

    \I__9327\ : InMux
    port map (
            O => \N__46984\,
            I => \N__46971\
        );

    \I__9326\ : Odrv4
    port map (
            O => \N__46981\,
            I => \CONTROL.N_361_1\
        );

    \I__9325\ : Odrv4
    port map (
            O => \N__46974\,
            I => \CONTROL.N_361_1\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__46971\,
            I => \CONTROL.N_361_1\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__46964\,
            I => \N__46961\
        );

    \I__9322\ : InMux
    port map (
            O => \N__46961\,
            I => \N__46958\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__46958\,
            I => \N__46955\
        );

    \I__9320\ : Span4Mux_h
    port map (
            O => \N__46955\,
            I => \N__46952\
        );

    \I__9319\ : Span4Mux_h
    port map (
            O => \N__46952\,
            I => \N__46949\
        );

    \I__9318\ : Odrv4
    port map (
            O => \N__46949\,
            I => \CONTROL.un1_busState114_2_0_0_0\
        );

    \I__9317\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46939\
        );

    \I__9316\ : CascadeMux
    port map (
            O => \N__46945\,
            I => \N__46936\
        );

    \I__9315\ : InMux
    port map (
            O => \N__46944\,
            I => \N__46932\
        );

    \I__9314\ : InMux
    port map (
            O => \N__46943\,
            I => \N__46927\
        );

    \I__9313\ : InMux
    port map (
            O => \N__46942\,
            I => \N__46927\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__46939\,
            I => \N__46919\
        );

    \I__9311\ : InMux
    port map (
            O => \N__46936\,
            I => \N__46914\
        );

    \I__9310\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46914\
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__46932\,
            I => \N__46909\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__46927\,
            I => \N__46909\
        );

    \I__9307\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46904\
        );

    \I__9306\ : InMux
    port map (
            O => \N__46925\,
            I => \N__46904\
        );

    \I__9305\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46899\
        );

    \I__9304\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46899\
        );

    \I__9303\ : CascadeMux
    port map (
            O => \N__46922\,
            I => \N__46893\
        );

    \I__9302\ : Span4Mux_v
    port map (
            O => \N__46919\,
            I => \N__46889\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__46914\,
            I => \N__46884\
        );

    \I__9300\ : Span4Mux_h
    port map (
            O => \N__46909\,
            I => \N__46884\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__46904\,
            I => \N__46881\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__46899\,
            I => \N__46878\
        );

    \I__9297\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46871\
        );

    \I__9296\ : InMux
    port map (
            O => \N__46897\,
            I => \N__46871\
        );

    \I__9295\ : InMux
    port map (
            O => \N__46896\,
            I => \N__46871\
        );

    \I__9294\ : InMux
    port map (
            O => \N__46893\,
            I => \N__46866\
        );

    \I__9293\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46866\
        );

    \I__9292\ : Span4Mux_h
    port map (
            O => \N__46889\,
            I => \N__46859\
        );

    \I__9291\ : Span4Mux_h
    port map (
            O => \N__46884\,
            I => \N__46859\
        );

    \I__9290\ : Span4Mux_v
    port map (
            O => \N__46881\,
            I => \N__46859\
        );

    \I__9289\ : Odrv4
    port map (
            O => \N__46878\,
            I => \aluOperand2_2_rep2\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__46871\,
            I => \aluOperand2_2_rep2\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__46866\,
            I => \aluOperand2_2_rep2\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__46859\,
            I => \aluOperand2_2_rep2\
        );

    \I__9285\ : InMux
    port map (
            O => \N__46850\,
            I => \N__46847\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__46847\,
            I => \ALU.c_RNI9SHFZ0Z_14\
        );

    \I__9283\ : CascadeMux
    port map (
            O => \N__46844\,
            I => \ALU.a_RNI5CPUZ0Z_14_cascade_\
        );

    \I__9282\ : InMux
    port map (
            O => \N__46841\,
            I => \N__46837\
        );

    \I__9281\ : InMux
    port map (
            O => \N__46840\,
            I => \N__46833\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__46837\,
            I => \N__46828\
        );

    \I__9279\ : InMux
    port map (
            O => \N__46836\,
            I => \N__46824\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__46833\,
            I => \N__46821\
        );

    \I__9277\ : InMux
    port map (
            O => \N__46832\,
            I => \N__46816\
        );

    \I__9276\ : InMux
    port map (
            O => \N__46831\,
            I => \N__46816\
        );

    \I__9275\ : Span4Mux_h
    port map (
            O => \N__46828\,
            I => \N__46808\
        );

    \I__9274\ : InMux
    port map (
            O => \N__46827\,
            I => \N__46805\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__46824\,
            I => \N__46798\
        );

    \I__9272\ : Span4Mux_h
    port map (
            O => \N__46821\,
            I => \N__46798\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__46816\,
            I => \N__46798\
        );

    \I__9270\ : InMux
    port map (
            O => \N__46815\,
            I => \N__46789\
        );

    \I__9269\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46789\
        );

    \I__9268\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46789\
        );

    \I__9267\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46789\
        );

    \I__9266\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46786\
        );

    \I__9265\ : Span4Mux_h
    port map (
            O => \N__46808\,
            I => \N__46783\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__46805\,
            I => \N__46776\
        );

    \I__9263\ : Span4Mux_h
    port map (
            O => \N__46798\,
            I => \N__46773\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__46789\,
            I => \N__46770\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__46786\,
            I => \N__46767\
        );

    \I__9260\ : Span4Mux_h
    port map (
            O => \N__46783\,
            I => \N__46764\
        );

    \I__9259\ : InMux
    port map (
            O => \N__46782\,
            I => \N__46761\
        );

    \I__9258\ : InMux
    port map (
            O => \N__46781\,
            I => \N__46756\
        );

    \I__9257\ : InMux
    port map (
            O => \N__46780\,
            I => \N__46756\
        );

    \I__9256\ : InMux
    port map (
            O => \N__46779\,
            I => \N__46753\
        );

    \I__9255\ : Span4Mux_h
    port map (
            O => \N__46776\,
            I => \N__46746\
        );

    \I__9254\ : Span4Mux_h
    port map (
            O => \N__46773\,
            I => \N__46746\
        );

    \I__9253\ : Span4Mux_h
    port map (
            O => \N__46770\,
            I => \N__46746\
        );

    \I__9252\ : Odrv12
    port map (
            O => \N__46767\,
            I => \aluOperand2_1\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__46764\,
            I => \aluOperand2_1\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__46761\,
            I => \aluOperand2_1\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__46756\,
            I => \aluOperand2_1\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__46753\,
            I => \aluOperand2_1\
        );

    \I__9247\ : Odrv4
    port map (
            O => \N__46746\,
            I => \aluOperand2_1\
        );

    \I__9246\ : InMux
    port map (
            O => \N__46733\,
            I => \N__46730\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__46730\,
            I => \N__46727\
        );

    \I__9244\ : Odrv12
    port map (
            O => \N__46727\,
            I => \ALU.d_RNICJCTZ0Z_14\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__46724\,
            I => \ALU.operand2_7_ns_1_14_cascade_\
        );

    \I__9242\ : InMux
    port map (
            O => \N__46721\,
            I => \N__46718\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__46718\,
            I => \N__46715\
        );

    \I__9240\ : Odrv4
    port map (
            O => \N__46715\,
            I => \ALU.b_RNI83KC1Z0Z_14\
        );

    \I__9239\ : InMux
    port map (
            O => \N__46712\,
            I => \N__46709\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__46709\,
            I => \N__46706\
        );

    \I__9237\ : Span4Mux_h
    port map (
            O => \N__46706\,
            I => \N__46703\
        );

    \I__9236\ : Odrv4
    port map (
            O => \N__46703\,
            I => \N_191\
        );

    \I__9235\ : CascadeMux
    port map (
            O => \N__46700\,
            I => \ALU.operand2_14_cascade_\
        );

    \I__9234\ : CascadeMux
    port map (
            O => \N__46697\,
            I => \N__46694\
        );

    \I__9233\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46691\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__46691\,
            I => \ALU.d_RNINISC7Z0Z_14\
        );

    \I__9231\ : CascadeMux
    port map (
            O => \N__46688\,
            I => \ALU.dout_3_ns_1_14_cascade_\
        );

    \I__9230\ : InMux
    port map (
            O => \N__46685\,
            I => \N__46679\
        );

    \I__9229\ : InMux
    port map (
            O => \N__46684\,
            I => \N__46679\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__46679\,
            I => \N__46676\
        );

    \I__9227\ : Span4Mux_h
    port map (
            O => \N__46676\,
            I => \N__46673\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__46673\,
            I => \N__46670\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__46670\,
            I => \ALU.cZ0Z_15\
        );

    \I__9224\ : InMux
    port map (
            O => \N__46667\,
            I => \N__46664\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__46664\,
            I => \N__46661\
        );

    \I__9222\ : Span4Mux_v
    port map (
            O => \N__46661\,
            I => \N__46658\
        );

    \I__9221\ : Span4Mux_h
    port map (
            O => \N__46658\,
            I => \N__46655\
        );

    \I__9220\ : Span4Mux_h
    port map (
            O => \N__46655\,
            I => \N__46651\
        );

    \I__9219\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46648\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__46651\,
            I => \ALU.cZ0Z_9\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__46648\,
            I => \ALU.cZ0Z_9\
        );

    \I__9216\ : CascadeMux
    port map (
            O => \N__46643\,
            I => \ALU.log_1_7_cascade_\
        );

    \I__9215\ : InMux
    port map (
            O => \N__46640\,
            I => \N__46637\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__46637\,
            I => \N__46634\
        );

    \I__9213\ : Span4Mux_v
    port map (
            O => \N__46634\,
            I => \N__46631\
        );

    \I__9212\ : Span4Mux_h
    port map (
            O => \N__46631\,
            I => \N__46628\
        );

    \I__9211\ : Odrv4
    port map (
            O => \N__46628\,
            I => \ALU.mult_7\
        );

    \I__9210\ : CascadeMux
    port map (
            O => \N__46625\,
            I => \ALU.mult_492_c_RNIQ5BZ0Z457_cascade_\
        );

    \I__9209\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46619\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__46619\,
            I => \N__46616\
        );

    \I__9207\ : Odrv12
    port map (
            O => \N__46616\,
            I => \ALU.lshift_7\
        );

    \I__9206\ : CascadeMux
    port map (
            O => \N__46613\,
            I => \ALU.mult_492_c_RNIGN2JECZ0_cascade_\
        );

    \I__9205\ : InMux
    port map (
            O => \N__46610\,
            I => \N__46606\
        );

    \I__9204\ : CascadeMux
    port map (
            O => \N__46609\,
            I => \N__46603\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__46606\,
            I => \N__46600\
        );

    \I__9202\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46597\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__46600\,
            I => \N__46594\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__46597\,
            I => \N__46591\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__46594\,
            I => \ALU.aZ0Z_7\
        );

    \I__9198\ : Odrv4
    port map (
            O => \N__46591\,
            I => \ALU.aZ0Z_7\
        );

    \I__9197\ : CascadeMux
    port map (
            O => \N__46586\,
            I => \N__46583\
        );

    \I__9196\ : InMux
    port map (
            O => \N__46583\,
            I => \N__46580\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__46580\,
            I => \N__46577\
        );

    \I__9194\ : Span4Mux_h
    port map (
            O => \N__46577\,
            I => \N__46574\
        );

    \I__9193\ : Span4Mux_v
    port map (
            O => \N__46574\,
            I => \N__46571\
        );

    \I__9192\ : Span4Mux_h
    port map (
            O => \N__46571\,
            I => \N__46568\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__46568\,
            I => \ALU.d_RNIO75BGZ0Z_7\
        );

    \I__9190\ : InMux
    port map (
            O => \N__46565\,
            I => \N__46562\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__46562\,
            I => \N__46559\
        );

    \I__9188\ : Span4Mux_h
    port map (
            O => \N__46559\,
            I => \N__46556\
        );

    \I__9187\ : Odrv4
    port map (
            O => \N__46556\,
            I => \ALU.c_RNIE4B6N4Z0Z_15\
        );

    \I__9186\ : CascadeMux
    port map (
            O => \N__46553\,
            I => \ALU.a_15_1_15_cascade_\
        );

    \I__9185\ : InMux
    port map (
            O => \N__46550\,
            I => \N__46546\
        );

    \I__9184\ : InMux
    port map (
            O => \N__46549\,
            I => \N__46543\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__46546\,
            I => \N__46538\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__46543\,
            I => \N__46538\
        );

    \I__9181\ : Span4Mux_v
    port map (
            O => \N__46538\,
            I => \N__46535\
        );

    \I__9180\ : Span4Mux_h
    port map (
            O => \N__46535\,
            I => \N__46532\
        );

    \I__9179\ : Sp12to4
    port map (
            O => \N__46532\,
            I => \N__46529\
        );

    \I__9178\ : Span12Mux_v
    port map (
            O => \N__46529\,
            I => \N__46526\
        );

    \I__9177\ : Odrv12
    port map (
            O => \N__46526\,
            I => \ALU.aZ0Z_15\
        );

    \I__9176\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46520\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__46520\,
            I => \ALU.N_812\
        );

    \I__9174\ : CascadeMux
    port map (
            O => \N__46517\,
            I => \ALU.N_812_cascade_\
        );

    \I__9173\ : InMux
    port map (
            O => \N__46514\,
            I => \N__46511\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__46511\,
            I => \ALU.addsub_cry_14_c_RNI134CVZ0Z5\
        );

    \I__9171\ : CascadeMux
    port map (
            O => \N__46508\,
            I => \N__46505\
        );

    \I__9170\ : InMux
    port map (
            O => \N__46505\,
            I => \N__46502\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__46502\,
            I => \N__46497\
        );

    \I__9168\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46494\
        );

    \I__9167\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46491\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__46497\,
            I => \N__46488\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__46494\,
            I => \ALU.N_635\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__46491\,
            I => \ALU.N_635\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__46488\,
            I => \ALU.N_635\
        );

    \I__9162\ : CascadeMux
    port map (
            O => \N__46481\,
            I => \N__46478\
        );

    \I__9161\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46472\
        );

    \I__9160\ : InMux
    port map (
            O => \N__46477\,
            I => \N__46472\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__46472\,
            I => \N__46469\
        );

    \I__9158\ : Span4Mux_v
    port map (
            O => \N__46469\,
            I => \N__46466\
        );

    \I__9157\ : Odrv4
    port map (
            O => \N__46466\,
            I => \ALU.N_639\
        );

    \I__9156\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46459\
        );

    \I__9155\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46456\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__46459\,
            I => \N__46453\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__46456\,
            I => \N__46450\
        );

    \I__9152\ : Span4Mux_v
    port map (
            O => \N__46453\,
            I => \N__46447\
        );

    \I__9151\ : Span4Mux_h
    port map (
            O => \N__46450\,
            I => \N__46444\
        );

    \I__9150\ : Span4Mux_h
    port map (
            O => \N__46447\,
            I => \N__46441\
        );

    \I__9149\ : Span4Mux_h
    port map (
            O => \N__46444\,
            I => \N__46438\
        );

    \I__9148\ : Odrv4
    port map (
            O => \N__46441\,
            I => \ALU.cZ0Z_1\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__46438\,
            I => \ALU.cZ0Z_1\
        );

    \I__9146\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46430\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__46430\,
            I => \N__46426\
        );

    \I__9144\ : InMux
    port map (
            O => \N__46429\,
            I => \N__46423\
        );

    \I__9143\ : Span4Mux_h
    port map (
            O => \N__46426\,
            I => \N__46420\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__46423\,
            I => \N__46417\
        );

    \I__9141\ : Span4Mux_h
    port map (
            O => \N__46420\,
            I => \N__46414\
        );

    \I__9140\ : Span4Mux_h
    port map (
            O => \N__46417\,
            I => \N__46411\
        );

    \I__9139\ : Span4Mux_v
    port map (
            O => \N__46414\,
            I => \N__46408\
        );

    \I__9138\ : Odrv4
    port map (
            O => \N__46411\,
            I => \ALU.cZ0Z_0\
        );

    \I__9137\ : Odrv4
    port map (
            O => \N__46408\,
            I => \ALU.cZ0Z_0\
        );

    \I__9136\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46399\
        );

    \I__9135\ : InMux
    port map (
            O => \N__46402\,
            I => \N__46396\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__46399\,
            I => \N__46393\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__46396\,
            I => \N__46390\
        );

    \I__9132\ : Span4Mux_v
    port map (
            O => \N__46393\,
            I => \N__46387\
        );

    \I__9131\ : Span4Mux_v
    port map (
            O => \N__46390\,
            I => \N__46382\
        );

    \I__9130\ : Span4Mux_h
    port map (
            O => \N__46387\,
            I => \N__46382\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__46382\,
            I => \ALU.cZ0Z_7\
        );

    \I__9128\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46373\
        );

    \I__9127\ : InMux
    port map (
            O => \N__46378\,
            I => \N__46373\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__46373\,
            I => \N__46370\
        );

    \I__9125\ : Span4Mux_h
    port map (
            O => \N__46370\,
            I => \N__46367\
        );

    \I__9124\ : Span4Mux_h
    port map (
            O => \N__46367\,
            I => \N__46364\
        );

    \I__9123\ : Span4Mux_h
    port map (
            O => \N__46364\,
            I => \N__46361\
        );

    \I__9122\ : Odrv4
    port map (
            O => \N__46361\,
            I => \ALU.cZ0Z_8\
        );

    \I__9121\ : CascadeMux
    port map (
            O => \N__46358\,
            I => \N__46355\
        );

    \I__9120\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46352\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__46352\,
            I => \N__46348\
        );

    \I__9118\ : CascadeMux
    port map (
            O => \N__46351\,
            I => \N__46345\
        );

    \I__9117\ : Span4Mux_h
    port map (
            O => \N__46348\,
            I => \N__46342\
        );

    \I__9116\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46339\
        );

    \I__9115\ : Span4Mux_v
    port map (
            O => \N__46342\,
            I => \N__46334\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__46339\,
            I => \N__46334\
        );

    \I__9113\ : Span4Mux_v
    port map (
            O => \N__46334\,
            I => \N__46331\
        );

    \I__9112\ : Span4Mux_h
    port map (
            O => \N__46331\,
            I => \N__46328\
        );

    \I__9111\ : Odrv4
    port map (
            O => \N__46328\,
            I => \ALU.eZ0Z_1\
        );

    \I__9110\ : InMux
    port map (
            O => \N__46325\,
            I => \N__46321\
        );

    \I__9109\ : InMux
    port map (
            O => \N__46324\,
            I => \N__46318\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__46321\,
            I => \N__46315\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__46318\,
            I => \N__46312\
        );

    \I__9106\ : Span4Mux_v
    port map (
            O => \N__46315\,
            I => \N__46307\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__46312\,
            I => \N__46307\
        );

    \I__9104\ : Span4Mux_h
    port map (
            O => \N__46307\,
            I => \N__46304\
        );

    \I__9103\ : Span4Mux_v
    port map (
            O => \N__46304\,
            I => \N__46301\
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__46301\,
            I => \ALU.eZ0Z_0\
        );

    \I__9101\ : CascadeMux
    port map (
            O => \N__46298\,
            I => \N__46295\
        );

    \I__9100\ : InMux
    port map (
            O => \N__46295\,
            I => \N__46289\
        );

    \I__9099\ : InMux
    port map (
            O => \N__46294\,
            I => \N__46289\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__46289\,
            I => \N__46286\
        );

    \I__9097\ : Sp12to4
    port map (
            O => \N__46286\,
            I => \N__46283\
        );

    \I__9096\ : Odrv12
    port map (
            O => \N__46283\,
            I => \ALU.eZ0Z_7\
        );

    \I__9095\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46276\
        );

    \I__9094\ : CascadeMux
    port map (
            O => \N__46279\,
            I => \N__46273\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__46276\,
            I => \N__46270\
        );

    \I__9092\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46267\
        );

    \I__9091\ : Span4Mux_h
    port map (
            O => \N__46270\,
            I => \N__46264\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__46267\,
            I => \N__46261\
        );

    \I__9089\ : Span4Mux_v
    port map (
            O => \N__46264\,
            I => \N__46258\
        );

    \I__9088\ : Span4Mux_v
    port map (
            O => \N__46261\,
            I => \N__46255\
        );

    \I__9087\ : Span4Mux_h
    port map (
            O => \N__46258\,
            I => \N__46252\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__46255\,
            I => \N__46249\
        );

    \I__9085\ : Sp12to4
    port map (
            O => \N__46252\,
            I => \N__46246\
        );

    \I__9084\ : Span4Mux_h
    port map (
            O => \N__46249\,
            I => \N__46243\
        );

    \I__9083\ : Odrv12
    port map (
            O => \N__46246\,
            I => \ALU.eZ0Z_8\
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__46243\,
            I => \ALU.eZ0Z_8\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__46238\,
            I => \N__46234\
        );

    \I__9080\ : CascadeMux
    port map (
            O => \N__46237\,
            I => \N__46231\
        );

    \I__9079\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46228\
        );

    \I__9078\ : InMux
    port map (
            O => \N__46231\,
            I => \N__46225\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__46228\,
            I => \N__46220\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__46225\,
            I => \N__46220\
        );

    \I__9075\ : Span4Mux_v
    port map (
            O => \N__46220\,
            I => \N__46217\
        );

    \I__9074\ : Span4Mux_h
    port map (
            O => \N__46217\,
            I => \N__46214\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__46214\,
            I => \ALU.eZ0Z_15\
        );

    \I__9072\ : CascadeMux
    port map (
            O => \N__46211\,
            I => \N__46208\
        );

    \I__9071\ : InMux
    port map (
            O => \N__46208\,
            I => \N__46204\
        );

    \I__9070\ : InMux
    port map (
            O => \N__46207\,
            I => \N__46201\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__46204\,
            I => \N__46198\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__46201\,
            I => \N__46195\
        );

    \I__9067\ : Span4Mux_v
    port map (
            O => \N__46198\,
            I => \N__46192\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__46195\,
            I => \N__46189\
        );

    \I__9065\ : Span4Mux_h
    port map (
            O => \N__46192\,
            I => \N__46186\
        );

    \I__9064\ : Span4Mux_h
    port map (
            O => \N__46189\,
            I => \N__46183\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__46186\,
            I => \ALU.eZ0Z_9\
        );

    \I__9062\ : Odrv4
    port map (
            O => \N__46183\,
            I => \ALU.eZ0Z_9\
        );

    \I__9061\ : InMux
    port map (
            O => \N__46178\,
            I => \N__46175\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__46175\,
            I => \N__46172\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__46172\,
            I => \N__46169\
        );

    \I__9058\ : Span4Mux_v
    port map (
            O => \N__46169\,
            I => \N__46166\
        );

    \I__9057\ : Odrv4
    port map (
            O => \N__46166\,
            I => \ALU.N_647\
        );

    \I__9056\ : InMux
    port map (
            O => \N__46163\,
            I => \N__46160\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__46160\,
            I => \N__46156\
        );

    \I__9054\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46153\
        );

    \I__9053\ : Span4Mux_h
    port map (
            O => \N__46156\,
            I => \N__46150\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__46153\,
            I => \N__46147\
        );

    \I__9051\ : Span4Mux_h
    port map (
            O => \N__46150\,
            I => \N__46144\
        );

    \I__9050\ : Odrv12
    port map (
            O => \N__46147\,
            I => \ALU.N_643\
        );

    \I__9049\ : Odrv4
    port map (
            O => \N__46144\,
            I => \ALU.N_643\
        );

    \I__9048\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46136\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__46136\,
            I => \ALU.N_707\
        );

    \I__9046\ : CascadeMux
    port map (
            O => \N__46133\,
            I => \ALU.addsub_cry_14_c_RNI134CV5Z0Z_0_cascade_\
        );

    \I__9045\ : CascadeMux
    port map (
            O => \N__46130\,
            I => \ALU.addsub_cry_14_c_RNIKS9S5HZ0_cascade_\
        );

    \I__9044\ : InMux
    port map (
            O => \N__46127\,
            I => \N__46124\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__46124\,
            I => \ALU.mult_335_c_RNOZ0Z_0\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__46121\,
            I => \ALU.N_835_cascade_\
        );

    \I__9041\ : InMux
    port map (
            O => \N__46118\,
            I => \N__46114\
        );

    \I__9040\ : CascadeMux
    port map (
            O => \N__46117\,
            I => \N__46111\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__46114\,
            I => \N__46108\
        );

    \I__9038\ : InMux
    port map (
            O => \N__46111\,
            I => \N__46105\
        );

    \I__9037\ : Odrv4
    port map (
            O => \N__46108\,
            I => \ALU.N_852\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__46105\,
            I => \ALU.N_852\
        );

    \I__9035\ : CascadeMux
    port map (
            O => \N__46100\,
            I => \ALU.rshift_7_ns_1_7_cascade_\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__46097\,
            I => \ALU.N_925_cascade_\
        );

    \I__9033\ : CascadeMux
    port map (
            O => \N__46094\,
            I => \N__46091\
        );

    \I__9032\ : InMux
    port map (
            O => \N__46091\,
            I => \N__46088\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__46088\,
            I => \N__46085\
        );

    \I__9030\ : Span4Mux_v
    port map (
            O => \N__46085\,
            I => \N__46082\
        );

    \I__9029\ : Sp12to4
    port map (
            O => \N__46082\,
            I => \N__46079\
        );

    \I__9028\ : Odrv12
    port map (
            O => \N__46079\,
            I => \ALU.N_833\
        );

    \I__9027\ : InMux
    port map (
            O => \N__46076\,
            I => \N__46070\
        );

    \I__9026\ : InMux
    port map (
            O => \N__46075\,
            I => \N__46070\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__46070\,
            I => \N__46067\
        );

    \I__9024\ : Span4Mux_h
    port map (
            O => \N__46067\,
            I => \N__46063\
        );

    \I__9023\ : InMux
    port map (
            O => \N__46066\,
            I => \N__46060\
        );

    \I__9022\ : Odrv4
    port map (
            O => \N__46063\,
            I => \ALU.N_837\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__46060\,
            I => \ALU.N_837\
        );

    \I__9020\ : CascadeMux
    port map (
            O => \N__46055\,
            I => \ALU.rshift_7_ns_1_3_cascade_\
        );

    \I__9019\ : InMux
    port map (
            O => \N__46052\,
            I => \N__46049\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__46049\,
            I => \N__46046\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__46046\,
            I => \ALU.N_921\
        );

    \I__9016\ : IoInMux
    port map (
            O => \N__46043\,
            I => \N__46040\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__46040\,
            I => \N__46036\
        );

    \I__9014\ : IoInMux
    port map (
            O => \N__46039\,
            I => \N__46033\
        );

    \I__9013\ : Span4Mux_s0_h
    port map (
            O => \N__46036\,
            I => \N__46029\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__46033\,
            I => \N__46026\
        );

    \I__9011\ : InMux
    port map (
            O => \N__46032\,
            I => \N__46023\
        );

    \I__9010\ : Span4Mux_h
    port map (
            O => \N__46029\,
            I => \N__46020\
        );

    \I__9009\ : IoSpan4Mux
    port map (
            O => \N__46026\,
            I => \N__46017\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__46023\,
            I => \N__46014\
        );

    \I__9007\ : Sp12to4
    port map (
            O => \N__46020\,
            I => \N__46011\
        );

    \I__9006\ : Span4Mux_s3_h
    port map (
            O => \N__46017\,
            I => \N__46008\
        );

    \I__9005\ : Span4Mux_v
    port map (
            O => \N__46014\,
            I => \N__46005\
        );

    \I__9004\ : Span12Mux_v
    port map (
            O => \N__46011\,
            I => \N__46002\
        );

    \I__9003\ : Sp12to4
    port map (
            O => \N__46008\,
            I => \N__45999\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__46005\,
            I => \N__45996\
        );

    \I__9001\ : Span12Mux_h
    port map (
            O => \N__46002\,
            I => \N__45991\
        );

    \I__9000\ : Span12Mux_v
    port map (
            O => \N__45999\,
            I => \N__45991\
        );

    \I__8999\ : Span4Mux_h
    port map (
            O => \N__45996\,
            I => \N__45988\
        );

    \I__8998\ : Odrv12
    port map (
            O => \N__45991\,
            I => bus_7
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__45988\,
            I => bus_7
        );

    \I__8996\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45980\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__45980\,
            I => \N__45977\
        );

    \I__8994\ : Span4Mux_v
    port map (
            O => \N__45977\,
            I => \N__45974\
        );

    \I__8993\ : Span4Mux_h
    port map (
            O => \N__45974\,
            I => \N__45971\
        );

    \I__8992\ : Odrv4
    port map (
            O => \N__45971\,
            I => \ALU.N_1030\
        );

    \I__8991\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45965\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__45965\,
            I => \ALU.c_RNI08R632Z0Z_15\
        );

    \I__8989\ : InMux
    port map (
            O => \N__45962\,
            I => \N__45959\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__45959\,
            I => \N__45956\
        );

    \I__8987\ : Span4Mux_v
    port map (
            O => \N__45956\,
            I => \N__45953\
        );

    \I__8986\ : Span4Mux_h
    port map (
            O => \N__45953\,
            I => \N__45950\
        );

    \I__8985\ : Odrv4
    port map (
            O => \N__45950\,
            I => \ALU.lshift_3_ns_1_11\
        );

    \I__8984\ : InMux
    port map (
            O => \N__45947\,
            I => \N__45944\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__45944\,
            I => \N__45941\
        );

    \I__8982\ : Odrv4
    port map (
            O => \N__45941\,
            I => \ALU.d_RNI4N3K21Z0Z_8\
        );

    \I__8981\ : CascadeMux
    port map (
            O => \N__45938\,
            I => \N__45935\
        );

    \I__8980\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45932\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__45932\,
            I => \ALU.d_RNIH8D821Z0Z_8\
        );

    \I__8978\ : CascadeMux
    port map (
            O => \N__45929\,
            I => \N__45926\
        );

    \I__8977\ : InMux
    port map (
            O => \N__45926\,
            I => \N__45923\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__45923\,
            I => \N__45920\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__45920\,
            I => \ALU.mult_335_c_RNOZ0\
        );

    \I__8974\ : InMux
    port map (
            O => \N__45917\,
            I => \N__45914\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__45914\,
            I => \ALU.c_RNIBQSTOZ0Z_11\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__45911\,
            I => \N__45908\
        );

    \I__8971\ : InMux
    port map (
            O => \N__45908\,
            I => \N__45905\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__45905\,
            I => \ALU.c_RNIG5G6F1Z0Z_10\
        );

    \I__8969\ : CascadeMux
    port map (
            O => \N__45902\,
            I => \N__45899\
        );

    \I__8968\ : InMux
    port map (
            O => \N__45899\,
            I => \N__45896\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__45896\,
            I => \ALU.mult_11_12\
        );

    \I__8966\ : InMux
    port map (
            O => \N__45893\,
            I => \ALU.mult_11_c11\
        );

    \I__8965\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45887\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__45887\,
            I => \N__45884\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__45884\,
            I => \N__45881\
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__45881\,
            I => \ALU.c_RNIN266MZ0Z_11\
        );

    \I__8961\ : CascadeMux
    port map (
            O => \N__45878\,
            I => \N__45875\
        );

    \I__8960\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45872\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__45872\,
            I => \ALU.c_RNIT73F71Z0Z_10\
        );

    \I__8958\ : CascadeMux
    port map (
            O => \N__45869\,
            I => \N__45866\
        );

    \I__8957\ : InMux
    port map (
            O => \N__45866\,
            I => \N__45863\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__45863\,
            I => \ALU.mult_11_13\
        );

    \I__8955\ : InMux
    port map (
            O => \N__45860\,
            I => \ALU.mult_11_c12\
        );

    \I__8954\ : CascadeMux
    port map (
            O => \N__45857\,
            I => \N__45854\
        );

    \I__8953\ : InMux
    port map (
            O => \N__45854\,
            I => \N__45851\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__45851\,
            I => \N__45848\
        );

    \I__8951\ : Span4Mux_v
    port map (
            O => \N__45848\,
            I => \N__45845\
        );

    \I__8950\ : Span4Mux_h
    port map (
            O => \N__45845\,
            I => \N__45842\
        );

    \I__8949\ : Span4Mux_h
    port map (
            O => \N__45842\,
            I => \N__45839\
        );

    \I__8948\ : Odrv4
    port map (
            O => \N__45839\,
            I => \ALU.c_RNIK31N31Z0Z_10\
        );

    \I__8947\ : CascadeMux
    port map (
            O => \N__45836\,
            I => \N__45833\
        );

    \I__8946\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45830\
        );

    \I__8945\ : LocalMux
    port map (
            O => \N__45830\,
            I => \ALU.mult_11_14\
        );

    \I__8944\ : InMux
    port map (
            O => \N__45827\,
            I => \ALU.mult_11_c13\
        );

    \I__8943\ : InMux
    port map (
            O => \N__45824\,
            I => \ALU.mult_11_c14\
        );

    \I__8942\ : InMux
    port map (
            O => \N__45821\,
            I => \N__45818\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__45818\,
            I => \ALU.mult_11_c14_THRU_CO\
        );

    \I__8940\ : InMux
    port map (
            O => \N__45815\,
            I => \N__45812\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__45812\,
            I => \ALU.c_RNIOSF6HZ0Z_11\
        );

    \I__8938\ : InMux
    port map (
            O => \N__45809\,
            I => \N__45806\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__45806\,
            I => \N__45802\
        );

    \I__8936\ : CascadeMux
    port map (
            O => \N__45805\,
            I => \N__45799\
        );

    \I__8935\ : Span4Mux_v
    port map (
            O => \N__45802\,
            I => \N__45796\
        );

    \I__8934\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45793\
        );

    \I__8933\ : Span4Mux_v
    port map (
            O => \N__45796\,
            I => \N__45790\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__45793\,
            I => \PROM.ROMDATA.m134\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__45790\,
            I => \PROM.ROMDATA.m134\
        );

    \I__8930\ : InMux
    port map (
            O => \N__45785\,
            I => \N__45782\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__45782\,
            I => \PROM.ROMDATA.m396_bm\
        );

    \I__8928\ : CascadeMux
    port map (
            O => \N__45779\,
            I => \PROM.ROMDATA.m396_am_cascade_\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__45776\,
            I => \PROM.ROMDATA.m396_ns_cascade_\
        );

    \I__8926\ : InMux
    port map (
            O => \N__45773\,
            I => \N__45770\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__45770\,
            I => \PROM.ROMDATA.m401_ns_1\
        );

    \I__8924\ : InMux
    port map (
            O => \N__45767\,
            I => \N__45763\
        );

    \I__8923\ : InMux
    port map (
            O => \N__45766\,
            I => \N__45760\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__45763\,
            I => \N__45757\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__45760\,
            I => \N__45754\
        );

    \I__8920\ : Span4Mux_h
    port map (
            O => \N__45757\,
            I => \N__45751\
        );

    \I__8919\ : Span4Mux_h
    port map (
            O => \N__45754\,
            I => \N__45748\
        );

    \I__8918\ : Span4Mux_v
    port map (
            O => \N__45751\,
            I => \N__45745\
        );

    \I__8917\ : Odrv4
    port map (
            O => \N__45748\,
            I => \PROM.ROMDATA.m401_ns\
        );

    \I__8916\ : Odrv4
    port map (
            O => \N__45745\,
            I => \PROM.ROMDATA.m401_ns\
        );

    \I__8915\ : CascadeMux
    port map (
            O => \N__45740\,
            I => \N__45737\
        );

    \I__8914\ : InMux
    port map (
            O => \N__45737\,
            I => \N__45734\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__45734\,
            I => \N__45731\
        );

    \I__8912\ : Odrv4
    port map (
            O => \N__45731\,
            I => \ALU.N_607\
        );

    \I__8911\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45725\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__45725\,
            I => \N__45720\
        );

    \I__8909\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45717\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__45723\,
            I => \N__45714\
        );

    \I__8907\ : Span4Mux_h
    port map (
            O => \N__45720\,
            I => \N__45711\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__45717\,
            I => \N__45708\
        );

    \I__8905\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45705\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__45711\,
            I => \N__45702\
        );

    \I__8903\ : Span4Mux_v
    port map (
            O => \N__45708\,
            I => \N__45699\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__45705\,
            I => \N__45696\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__45702\,
            I => \N__45693\
        );

    \I__8900\ : Span4Mux_h
    port map (
            O => \N__45699\,
            I => \N__45690\
        );

    \I__8899\ : Odrv12
    port map (
            O => \N__45696\,
            I => \ALU.N_767\
        );

    \I__8898\ : Odrv4
    port map (
            O => \N__45693\,
            I => \ALU.N_767\
        );

    \I__8897\ : Odrv4
    port map (
            O => \N__45690\,
            I => \ALU.N_767\
        );

    \I__8896\ : CascadeMux
    port map (
            O => \N__45683\,
            I => \ALU.N_607_cascade_\
        );

    \I__8895\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45677\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__45677\,
            I => \N__45674\
        );

    \I__8893\ : Span12Mux_v
    port map (
            O => \N__45674\,
            I => \N__45670\
        );

    \I__8892\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45667\
        );

    \I__8891\ : Odrv12
    port map (
            O => \N__45670\,
            I => \CONTROL.ctrlOut_5\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__45667\,
            I => \CONTROL.ctrlOut_5\
        );

    \I__8889\ : InMux
    port map (
            O => \N__45662\,
            I => \N__45659\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__45659\,
            I => \N__45655\
        );

    \I__8887\ : InMux
    port map (
            O => \N__45658\,
            I => \N__45652\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__45655\,
            I => \N__45649\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__45652\,
            I => \N__45646\
        );

    \I__8884\ : Odrv4
    port map (
            O => \N__45649\,
            I => \CONTROL.dout_reto_5\
        );

    \I__8883\ : Odrv4
    port map (
            O => \N__45646\,
            I => \CONTROL.dout_reto_5\
        );

    \I__8882\ : InMux
    port map (
            O => \N__45641\,
            I => \N__45638\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__45638\,
            I => \N__45635\
        );

    \I__8880\ : Odrv12
    port map (
            O => \N__45635\,
            I => \CONTROL.programCounter_ret_19_RNIV5IGZ0Z_6\
        );

    \I__8879\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45629\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__45629\,
            I => \N__45626\
        );

    \I__8877\ : Span4Mux_h
    port map (
            O => \N__45626\,
            I => \N__45623\
        );

    \I__8876\ : Span4Mux_h
    port map (
            O => \N__45623\,
            I => \N__45620\
        );

    \I__8875\ : Span4Mux_h
    port map (
            O => \N__45620\,
            I => \N__45617\
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__45617\,
            I => \CONTROL.addrstack_6\
        );

    \I__8873\ : InMux
    port map (
            O => \N__45614\,
            I => \N__45610\
        );

    \I__8872\ : InMux
    port map (
            O => \N__45613\,
            I => \N__45607\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__45610\,
            I => \N__45604\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__45607\,
            I => \CONTROL.addrstack_reto_6\
        );

    \I__8869\ : Odrv12
    port map (
            O => \N__45604\,
            I => \CONTROL.addrstack_reto_6\
        );

    \I__8868\ : InMux
    port map (
            O => \N__45599\,
            I => \N__45596\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__45596\,
            I => \PROM.ROMDATA.m48\
        );

    \I__8866\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45590\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__45590\,
            I => \N__45587\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__45587\,
            I => \N__45584\
        );

    \I__8863\ : Sp12to4
    port map (
            O => \N__45584\,
            I => \N__45580\
        );

    \I__8862\ : InMux
    port map (
            O => \N__45583\,
            I => \N__45577\
        );

    \I__8861\ : Odrv12
    port map (
            O => \N__45580\,
            I => \CONTROL.ctrlOut_6\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__45577\,
            I => \CONTROL.ctrlOut_6\
        );

    \I__8859\ : InMux
    port map (
            O => \N__45572\,
            I => \N__45569\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__45569\,
            I => \CONTROL.dout_reto_6\
        );

    \I__8857\ : InMux
    port map (
            O => \N__45566\,
            I => \N__45563\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__45563\,
            I => \PROM.ROMDATA.m7\
        );

    \I__8855\ : CascadeMux
    port map (
            O => \N__45560\,
            I => \PROM.ROMDATA.m392_bm_cascade_\
        );

    \I__8854\ : CascadeMux
    port map (
            O => \N__45557\,
            I => \PROM.ROMDATA.m392_ns_cascade_\
        );

    \I__8853\ : CascadeMux
    port map (
            O => \N__45554\,
            I => \N__45551\
        );

    \I__8852\ : InMux
    port map (
            O => \N__45551\,
            I => \N__45548\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__45548\,
            I => \N__45545\
        );

    \I__8850\ : Odrv12
    port map (
            O => \N__45545\,
            I => \PROM.ROMDATA.m36\
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__45542\,
            I => \PROM.ROMDATA.N_526_mux_cascade_\
        );

    \I__8848\ : InMux
    port map (
            O => \N__45539\,
            I => \N__45536\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__45536\,
            I => \N__45533\
        );

    \I__8846\ : Span4Mux_h
    port map (
            O => \N__45533\,
            I => \N__45530\
        );

    \I__8845\ : Span4Mux_v
    port map (
            O => \N__45530\,
            I => \N__45527\
        );

    \I__8844\ : Odrv4
    port map (
            O => \N__45527\,
            I => \PROM.ROMDATA.m238_bm\
        );

    \I__8843\ : CascadeMux
    port map (
            O => \N__45524\,
            I => \N__45520\
        );

    \I__8842\ : CascadeMux
    port map (
            O => \N__45523\,
            I => \N__45517\
        );

    \I__8841\ : InMux
    port map (
            O => \N__45520\,
            I => \N__45510\
        );

    \I__8840\ : InMux
    port map (
            O => \N__45517\,
            I => \N__45510\
        );

    \I__8839\ : CascadeMux
    port map (
            O => \N__45516\,
            I => \N__45506\
        );

    \I__8838\ : CascadeMux
    port map (
            O => \N__45515\,
            I => \N__45502\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__45510\,
            I => \N__45499\
        );

    \I__8836\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45492\
        );

    \I__8835\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45492\
        );

    \I__8834\ : InMux
    port map (
            O => \N__45505\,
            I => \N__45492\
        );

    \I__8833\ : InMux
    port map (
            O => \N__45502\,
            I => \N__45489\
        );

    \I__8832\ : Span4Mux_h
    port map (
            O => \N__45499\,
            I => \N__45486\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__45492\,
            I => \N__45483\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__45489\,
            I => \N__45480\
        );

    \I__8829\ : Span4Mux_h
    port map (
            O => \N__45486\,
            I => \N__45476\
        );

    \I__8828\ : Span4Mux_h
    port map (
            O => \N__45483\,
            I => \N__45473\
        );

    \I__8827\ : Span4Mux_v
    port map (
            O => \N__45480\,
            I => \N__45470\
        );

    \I__8826\ : CascadeMux
    port map (
            O => \N__45479\,
            I => \N__45467\
        );

    \I__8825\ : Span4Mux_h
    port map (
            O => \N__45476\,
            I => \N__45464\
        );

    \I__8824\ : Span4Mux_v
    port map (
            O => \N__45473\,
            I => \N__45461\
        );

    \I__8823\ : Span4Mux_v
    port map (
            O => \N__45470\,
            I => \N__45458\
        );

    \I__8822\ : InMux
    port map (
            O => \N__45467\,
            I => \N__45455\
        );

    \I__8821\ : Span4Mux_v
    port map (
            O => \N__45464\,
            I => \N__45452\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__45461\,
            I => \N__45449\
        );

    \I__8819\ : Span4Mux_h
    port map (
            O => \N__45458\,
            I => \N__45445\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__45455\,
            I => \N__45442\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__45452\,
            I => \N__45439\
        );

    \I__8816\ : Span4Mux_h
    port map (
            O => \N__45449\,
            I => \N__45436\
        );

    \I__8815\ : InMux
    port map (
            O => \N__45448\,
            I => \N__45433\
        );

    \I__8814\ : Span4Mux_v
    port map (
            O => \N__45445\,
            I => \N__45430\
        );

    \I__8813\ : Span12Mux_v
    port map (
            O => \N__45442\,
            I => \N__45427\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__45439\,
            I => \N__45424\
        );

    \I__8811\ : Span4Mux_v
    port map (
            O => \N__45436\,
            I => \N__45421\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__45433\,
            I => \aluStatus_i_3\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__45430\,
            I => \aluStatus_i_3\
        );

    \I__8808\ : Odrv12
    port map (
            O => \N__45427\,
            I => \aluStatus_i_3\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__45424\,
            I => \aluStatus_i_3\
        );

    \I__8806\ : Odrv4
    port map (
            O => \N__45421\,
            I => \aluStatus_i_3\
        );

    \I__8805\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45407\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__45407\,
            I => \N__45404\
        );

    \I__8803\ : Span4Mux_v
    port map (
            O => \N__45404\,
            I => \N__45398\
        );

    \I__8802\ : InMux
    port map (
            O => \N__45403\,
            I => \N__45393\
        );

    \I__8801\ : InMux
    port map (
            O => \N__45402\,
            I => \N__45393\
        );

    \I__8800\ : InMux
    port map (
            O => \N__45401\,
            I => \N__45387\
        );

    \I__8799\ : Span4Mux_h
    port map (
            O => \N__45398\,
            I => \N__45382\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__45393\,
            I => \N__45382\
        );

    \I__8797\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45375\
        );

    \I__8796\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45375\
        );

    \I__8795\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45375\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__45387\,
            I => \PROM_ROMDATA_dintern_10ro\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__45382\,
            I => \PROM_ROMDATA_dintern_10ro\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__45375\,
            I => \PROM_ROMDATA_dintern_10ro\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__45368\,
            I => \N__45365\
        );

    \I__8790\ : InMux
    port map (
            O => \N__45365\,
            I => \N__45362\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__45362\,
            I => \N__45359\
        );

    \I__8788\ : Odrv12
    port map (
            O => \N__45359\,
            I => \CONTROL.g0_5Z0Z_0\
        );

    \I__8787\ : InMux
    port map (
            O => \N__45356\,
            I => \N__45353\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__45353\,
            I => \N__45350\
        );

    \I__8785\ : Span4Mux_h
    port map (
            O => \N__45350\,
            I => \N__45347\
        );

    \I__8784\ : Odrv4
    port map (
            O => \N__45347\,
            I => \PROM.ROMDATA.m258_am\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__45344\,
            I => \N__45340\
        );

    \I__8782\ : InMux
    port map (
            O => \N__45343\,
            I => \N__45335\
        );

    \I__8781\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45335\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__45335\,
            I => \N__45332\
        );

    \I__8779\ : Span4Mux_h
    port map (
            O => \N__45332\,
            I => \N__45329\
        );

    \I__8778\ : Odrv4
    port map (
            O => \N__45329\,
            I => \PROM_ROMDATA_dintern_31_0__N_555_mux\
        );

    \I__8777\ : CascadeMux
    port map (
            O => \N__45326\,
            I => \N_417_cascade_\
        );

    \I__8776\ : InMux
    port map (
            O => \N__45323\,
            I => \N__45320\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__45320\,
            I => \N__45317\
        );

    \I__8774\ : Span4Mux_v
    port map (
            O => \N__45317\,
            I => \N__45313\
        );

    \I__8773\ : InMux
    port map (
            O => \N__45316\,
            I => \N__45310\
        );

    \I__8772\ : Span4Mux_h
    port map (
            O => \N__45313\,
            I => \N__45305\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__45310\,
            I => \N__45305\
        );

    \I__8770\ : Span4Mux_h
    port map (
            O => \N__45305\,
            I => \N__45302\
        );

    \I__8769\ : Span4Mux_v
    port map (
            O => \N__45302\,
            I => \N__45299\
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__45299\,
            I => \CONTROL.programCounter_1_2\
        );

    \I__8767\ : InMux
    port map (
            O => \N__45296\,
            I => \N__45293\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__45293\,
            I => \CONTROL.programCounter_ret_1_RNI6OHFZ0Z_6\
        );

    \I__8765\ : InMux
    port map (
            O => \N__45290\,
            I => \N__45287\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__45287\,
            I => \N__45284\
        );

    \I__8763\ : Span4Mux_v
    port map (
            O => \N__45284\,
            I => \N__45281\
        );

    \I__8762\ : Span4Mux_h
    port map (
            O => \N__45281\,
            I => \N__45277\
        );

    \I__8761\ : InMux
    port map (
            O => \N__45280\,
            I => \N__45274\
        );

    \I__8760\ : Sp12to4
    port map (
            O => \N__45277\,
            I => \N__45269\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__45274\,
            I => \N__45269\
        );

    \I__8758\ : Odrv12
    port map (
            O => \N__45269\,
            I => \CONTROL.ctrlOut_3\
        );

    \I__8757\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45263\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__45263\,
            I => \N__45259\
        );

    \I__8755\ : InMux
    port map (
            O => \N__45262\,
            I => \N__45256\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__45259\,
            I => \N__45253\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__45256\,
            I => \N__45250\
        );

    \I__8752\ : Span4Mux_h
    port map (
            O => \N__45253\,
            I => \N__45245\
        );

    \I__8751\ : Span4Mux_v
    port map (
            O => \N__45250\,
            I => \N__45245\
        );

    \I__8750\ : Odrv4
    port map (
            O => \N__45245\,
            I => \CONTROL.programCounter_1_4\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__45242\,
            I => \PROM.ROMDATA.m215_ns_1_N_2L1_cascade_\
        );

    \I__8748\ : InMux
    port map (
            O => \N__45239\,
            I => \N__45233\
        );

    \I__8747\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45233\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__45233\,
            I => \N__45230\
        );

    \I__8745\ : Span4Mux_h
    port map (
            O => \N__45230\,
            I => \N__45227\
        );

    \I__8744\ : Span4Mux_v
    port map (
            O => \N__45227\,
            I => \N__45224\
        );

    \I__8743\ : Odrv4
    port map (
            O => \N__45224\,
            I => \PROM.ROMDATA.m215_ns_1\
        );

    \I__8742\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45218\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__45218\,
            I => \N__45215\
        );

    \I__8740\ : Span4Mux_v
    port map (
            O => \N__45215\,
            I => \N__45212\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__45212\,
            I => \N__45209\
        );

    \I__8738\ : Odrv4
    port map (
            O => \N__45209\,
            I => \CONTROL.g0_3_i_a7_0_0\
        );

    \I__8737\ : InMux
    port map (
            O => \N__45206\,
            I => \N__45203\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__45203\,
            I => \N__45200\
        );

    \I__8735\ : Span12Mux_v
    port map (
            O => \N__45200\,
            I => \N__45197\
        );

    \I__8734\ : Odrv12
    port map (
            O => \N__45197\,
            I => \CONTROL.addrstack_2\
        );

    \I__8733\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45191\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__45191\,
            I => \PROM.ROMDATA.m258_bm\
        );

    \I__8731\ : InMux
    port map (
            O => \N__45188\,
            I => \N__45184\
        );

    \I__8730\ : InMux
    port map (
            O => \N__45187\,
            I => \N__45181\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__45184\,
            I => \N__45178\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__45181\,
            I => \N__45175\
        );

    \I__8727\ : Span4Mux_h
    port map (
            O => \N__45178\,
            I => \N__45172\
        );

    \I__8726\ : Span12Mux_h
    port map (
            O => \N__45175\,
            I => \N__45169\
        );

    \I__8725\ : Span4Mux_v
    port map (
            O => \N__45172\,
            I => \N__45166\
        );

    \I__8724\ : Odrv12
    port map (
            O => \N__45169\,
            I => \CONTROL.programCounter_1_1\
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__45166\,
            I => \CONTROL.programCounter_1_1\
        );

    \I__8722\ : InMux
    port map (
            O => \N__45161\,
            I => \N__45158\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__45158\,
            I => \CONTROL.programCounter_ret_19_RNIT3IGZ0Z_5\
        );

    \I__8720\ : InMux
    port map (
            O => \N__45155\,
            I => \N__45152\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__45152\,
            I => \N__45149\
        );

    \I__8718\ : Odrv4
    port map (
            O => \N__45149\,
            I => \CONTROL.programCounter_ret_1_RNI4MHFZ0Z_5\
        );

    \I__8717\ : InMux
    port map (
            O => \N__45146\,
            I => \N__45138\
        );

    \I__8716\ : InMux
    port map (
            O => \N__45145\,
            I => \N__45138\
        );

    \I__8715\ : InMux
    port map (
            O => \N__45144\,
            I => \N__45133\
        );

    \I__8714\ : InMux
    port map (
            O => \N__45143\,
            I => \N__45133\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__45138\,
            I => \N__45130\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__45133\,
            I => \N__45127\
        );

    \I__8711\ : Span4Mux_v
    port map (
            O => \N__45130\,
            I => \N__45122\
        );

    \I__8710\ : Span4Mux_h
    port map (
            O => \N__45127\,
            I => \N__45122\
        );

    \I__8709\ : Span4Mux_h
    port map (
            O => \N__45122\,
            I => \N__45116\
        );

    \I__8708\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45113\
        );

    \I__8707\ : InMux
    port map (
            O => \N__45120\,
            I => \N__45110\
        );

    \I__8706\ : InMux
    port map (
            O => \N__45119\,
            I => \N__45107\
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__45116\,
            I => \CONTROL.un1_programCounter9_reto\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__45113\,
            I => \CONTROL.un1_programCounter9_reto\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__45110\,
            I => \CONTROL.un1_programCounter9_reto\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__45107\,
            I => \CONTROL.un1_programCounter9_reto\
        );

    \I__8701\ : CascadeMux
    port map (
            O => \N__45098\,
            I => \progRomAddress_5_cascade_\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__45095\,
            I => \PROM.ROMDATA.m243_1_cascade_\
        );

    \I__8699\ : InMux
    port map (
            O => \N__45092\,
            I => \N__45089\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__45089\,
            I => \N__45086\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__45086\,
            I => \N__45083\
        );

    \I__8696\ : Odrv4
    port map (
            O => \N__45083\,
            I => \PROM.ROMDATA.m244_ns_1_1\
        );

    \I__8695\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45077\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__45077\,
            I => \N__45073\
        );

    \I__8693\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45070\
        );

    \I__8692\ : Odrv12
    port map (
            O => \N__45073\,
            I => \CONTROL.ctrlOut_0\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__45070\,
            I => \CONTROL.ctrlOut_0\
        );

    \I__8690\ : InMux
    port map (
            O => \N__45065\,
            I => \N__45062\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__45062\,
            I => \PROM.ROMDATA.m243_1\
        );

    \I__8688\ : CascadeMux
    port map (
            O => \N__45059\,
            I => \N__45055\
        );

    \I__8687\ : CascadeMux
    port map (
            O => \N__45058\,
            I => \N__45052\
        );

    \I__8686\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45045\
        );

    \I__8685\ : InMux
    port map (
            O => \N__45052\,
            I => \N__45045\
        );

    \I__8684\ : InMux
    port map (
            O => \N__45051\,
            I => \N__45040\
        );

    \I__8683\ : InMux
    port map (
            O => \N__45050\,
            I => \N__45040\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__45045\,
            I => \N__45035\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__45040\,
            I => \N__45035\
        );

    \I__8680\ : Span4Mux_h
    port map (
            O => \N__45035\,
            I => \N__45032\
        );

    \I__8679\ : Span4Mux_v
    port map (
            O => \N__45032\,
            I => \N__45028\
        );

    \I__8678\ : InMux
    port map (
            O => \N__45031\,
            I => \N__45025\
        );

    \I__8677\ : Odrv4
    port map (
            O => \N__45028\,
            I => \PROM.ROMDATA.m260_1\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__45025\,
            I => \PROM.ROMDATA.m260_1\
        );

    \I__8675\ : InMux
    port map (
            O => \N__45020\,
            I => \N__45017\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__45017\,
            I => \N__45014\
        );

    \I__8673\ : Span4Mux_h
    port map (
            O => \N__45014\,
            I => \N__45011\
        );

    \I__8672\ : Span4Mux_h
    port map (
            O => \N__45011\,
            I => \N__45006\
        );

    \I__8671\ : InMux
    port map (
            O => \N__45010\,
            I => \N__45003\
        );

    \I__8670\ : InMux
    port map (
            O => \N__45009\,
            I => \N__45000\
        );

    \I__8669\ : Span4Mux_h
    port map (
            O => \N__45006\,
            I => \N__44995\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__45003\,
            I => \N__44995\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__45000\,
            I => \N__44992\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__44995\,
            I => \N__44989\
        );

    \I__8665\ : Span4Mux_h
    port map (
            O => \N__44992\,
            I => \N__44986\
        );

    \I__8664\ : Span4Mux_h
    port map (
            O => \N__44989\,
            I => \N__44983\
        );

    \I__8663\ : Odrv4
    port map (
            O => \N__44986\,
            I => \controlWord_31\
        );

    \I__8662\ : Odrv4
    port map (
            O => \N__44983\,
            I => \controlWord_31\
        );

    \I__8661\ : IoInMux
    port map (
            O => \N__44978\,
            I => \N__44975\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__44975\,
            I => \N__44972\
        );

    \I__8659\ : IoSpan4Mux
    port map (
            O => \N__44972\,
            I => \N__44969\
        );

    \I__8658\ : Span4Mux_s1_v
    port map (
            O => \N__44969\,
            I => \N__44966\
        );

    \I__8657\ : Sp12to4
    port map (
            O => \N__44966\,
            I => \N__44963\
        );

    \I__8656\ : Span12Mux_h
    port map (
            O => \N__44963\,
            I => \N__44959\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__44962\,
            I => \N__44956\
        );

    \I__8654\ : Span12Mux_v
    port map (
            O => \N__44959\,
            I => \N__44953\
        );

    \I__8653\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44950\
        );

    \I__8652\ : Odrv12
    port map (
            O => \N__44953\,
            I => \A15_c\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__44950\,
            I => \A15_c\
        );

    \I__8650\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44942\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__44942\,
            I => \PROM.ROMDATA.m266\
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__44939\,
            I => \PROM.ROMDATA.m157_cascade_\
        );

    \I__8647\ : CascadeMux
    port map (
            O => \N__44936\,
            I => \PROM.ROMDATA.m265_cascade_\
        );

    \I__8646\ : InMux
    port map (
            O => \N__44933\,
            I => \N__44930\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__44930\,
            I => \PROM.ROMDATA.m268\
        );

    \I__8644\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44924\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__44924\,
            I => \N__44921\
        );

    \I__8642\ : Span4Mux_h
    port map (
            O => \N__44921\,
            I => \N__44917\
        );

    \I__8641\ : InMux
    port map (
            O => \N__44920\,
            I => \N__44914\
        );

    \I__8640\ : Odrv4
    port map (
            O => \N__44917\,
            I => \PROM.ROMDATA.m270_bm\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__44914\,
            I => \PROM.ROMDATA.m270_bm\
        );

    \I__8638\ : InMux
    port map (
            O => \N__44909\,
            I => \N__44906\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__44906\,
            I => \CONTROL.aluOperation_12_i_0_6\
        );

    \I__8636\ : InMux
    port map (
            O => \N__44903\,
            I => \N__44891\
        );

    \I__8635\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44891\
        );

    \I__8634\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44888\
        );

    \I__8633\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44885\
        );

    \I__8632\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44879\
        );

    \I__8631\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44872\
        );

    \I__8630\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44872\
        );

    \I__8629\ : InMux
    port map (
            O => \N__44896\,
            I => \N__44872\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__44891\,
            I => \N__44859\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__44888\,
            I => \N__44854\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__44885\,
            I => \N__44854\
        );

    \I__8625\ : InMux
    port map (
            O => \N__44884\,
            I => \N__44849\
        );

    \I__8624\ : InMux
    port map (
            O => \N__44883\,
            I => \N__44849\
        );

    \I__8623\ : InMux
    port map (
            O => \N__44882\,
            I => \N__44846\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__44879\,
            I => \N__44841\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__44872\,
            I => \N__44841\
        );

    \I__8620\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44836\
        );

    \I__8619\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44827\
        );

    \I__8618\ : InMux
    port map (
            O => \N__44869\,
            I => \N__44827\
        );

    \I__8617\ : InMux
    port map (
            O => \N__44868\,
            I => \N__44827\
        );

    \I__8616\ : InMux
    port map (
            O => \N__44867\,
            I => \N__44827\
        );

    \I__8615\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44824\
        );

    \I__8614\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44819\
        );

    \I__8613\ : InMux
    port map (
            O => \N__44864\,
            I => \N__44819\
        );

    \I__8612\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44816\
        );

    \I__8611\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44813\
        );

    \I__8610\ : Span4Mux_h
    port map (
            O => \N__44859\,
            I => \N__44810\
        );

    \I__8609\ : Span4Mux_h
    port map (
            O => \N__44854\,
            I => \N__44801\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__44849\,
            I => \N__44801\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__44846\,
            I => \N__44801\
        );

    \I__8606\ : Span4Mux_h
    port map (
            O => \N__44841\,
            I => \N__44801\
        );

    \I__8605\ : InMux
    port map (
            O => \N__44840\,
            I => \N__44796\
        );

    \I__8604\ : InMux
    port map (
            O => \N__44839\,
            I => \N__44796\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__44836\,
            I => \N__44791\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__44827\,
            I => \N__44791\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__44824\,
            I => \controlWord_3\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__44819\,
            I => \controlWord_3\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__44816\,
            I => \controlWord_3\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__44813\,
            I => \controlWord_3\
        );

    \I__8597\ : Odrv4
    port map (
            O => \N__44810\,
            I => \controlWord_3\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__44801\,
            I => \controlWord_3\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__44796\,
            I => \controlWord_3\
        );

    \I__8594\ : Odrv4
    port map (
            O => \N__44791\,
            I => \controlWord_3\
        );

    \I__8593\ : CascadeMux
    port map (
            O => \N__44774\,
            I => \N__44770\
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__44773\,
            I => \N__44766\
        );

    \I__8591\ : InMux
    port map (
            O => \N__44770\,
            I => \N__44763\
        );

    \I__8590\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44760\
        );

    \I__8589\ : InMux
    port map (
            O => \N__44766\,
            I => \N__44756\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__44763\,
            I => \N__44753\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__44760\,
            I => \N__44750\
        );

    \I__8586\ : CascadeMux
    port map (
            O => \N__44759\,
            I => \N__44745\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__44756\,
            I => \N__44742\
        );

    \I__8584\ : Span4Mux_h
    port map (
            O => \N__44753\,
            I => \N__44739\
        );

    \I__8583\ : Span4Mux_h
    port map (
            O => \N__44750\,
            I => \N__44736\
        );

    \I__8582\ : InMux
    port map (
            O => \N__44749\,
            I => \N__44731\
        );

    \I__8581\ : InMux
    port map (
            O => \N__44748\,
            I => \N__44731\
        );

    \I__8580\ : InMux
    port map (
            O => \N__44745\,
            I => \N__44728\
        );

    \I__8579\ : Span4Mux_h
    port map (
            O => \N__44742\,
            I => \N__44725\
        );

    \I__8578\ : Odrv4
    port map (
            O => \N__44739\,
            I => \CONTROL.N_219\
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__44736\,
            I => \CONTROL.N_219\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__44731\,
            I => \CONTROL.N_219\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__44728\,
            I => \CONTROL.N_219\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__44725\,
            I => \CONTROL.N_219\
        );

    \I__8573\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44709\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__44713\,
            I => \N__44697\
        );

    \I__8571\ : InMux
    port map (
            O => \N__44712\,
            I => \N__44693\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__44709\,
            I => \N__44690\
        );

    \I__8569\ : InMux
    port map (
            O => \N__44708\,
            I => \N__44687\
        );

    \I__8568\ : InMux
    port map (
            O => \N__44707\,
            I => \N__44680\
        );

    \I__8567\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44680\
        );

    \I__8566\ : InMux
    port map (
            O => \N__44705\,
            I => \N__44680\
        );

    \I__8565\ : InMux
    port map (
            O => \N__44704\,
            I => \N__44676\
        );

    \I__8564\ : InMux
    port map (
            O => \N__44703\,
            I => \N__44673\
        );

    \I__8563\ : InMux
    port map (
            O => \N__44702\,
            I => \N__44670\
        );

    \I__8562\ : InMux
    port map (
            O => \N__44701\,
            I => \N__44667\
        );

    \I__8561\ : InMux
    port map (
            O => \N__44700\,
            I => \N__44664\
        );

    \I__8560\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44651\
        );

    \I__8559\ : InMux
    port map (
            O => \N__44696\,
            I => \N__44646\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__44693\,
            I => \N__44641\
        );

    \I__8557\ : Span4Mux_v
    port map (
            O => \N__44690\,
            I => \N__44641\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__44687\,
            I => \N__44626\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__44680\,
            I => \N__44626\
        );

    \I__8554\ : InMux
    port map (
            O => \N__44679\,
            I => \N__44623\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__44676\,
            I => \N__44620\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__44673\,
            I => \N__44615\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__44670\,
            I => \N__44615\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__44667\,
            I => \N__44612\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__44664\,
            I => \N__44609\
        );

    \I__8548\ : InMux
    port map (
            O => \N__44663\,
            I => \N__44604\
        );

    \I__8547\ : InMux
    port map (
            O => \N__44662\,
            I => \N__44604\
        );

    \I__8546\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44601\
        );

    \I__8545\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44594\
        );

    \I__8544\ : InMux
    port map (
            O => \N__44659\,
            I => \N__44594\
        );

    \I__8543\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44594\
        );

    \I__8542\ : InMux
    port map (
            O => \N__44657\,
            I => \N__44585\
        );

    \I__8541\ : InMux
    port map (
            O => \N__44656\,
            I => \N__44585\
        );

    \I__8540\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44585\
        );

    \I__8539\ : InMux
    port map (
            O => \N__44654\,
            I => \N__44585\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__44651\,
            I => \N__44582\
        );

    \I__8537\ : InMux
    port map (
            O => \N__44650\,
            I => \N__44579\
        );

    \I__8536\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44576\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__44646\,
            I => \N__44573\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__44641\,
            I => \N__44570\
        );

    \I__8533\ : InMux
    port map (
            O => \N__44640\,
            I => \N__44565\
        );

    \I__8532\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44565\
        );

    \I__8531\ : InMux
    port map (
            O => \N__44638\,
            I => \N__44560\
        );

    \I__8530\ : InMux
    port map (
            O => \N__44637\,
            I => \N__44560\
        );

    \I__8529\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44549\
        );

    \I__8528\ : InMux
    port map (
            O => \N__44635\,
            I => \N__44549\
        );

    \I__8527\ : InMux
    port map (
            O => \N__44634\,
            I => \N__44549\
        );

    \I__8526\ : InMux
    port map (
            O => \N__44633\,
            I => \N__44549\
        );

    \I__8525\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44549\
        );

    \I__8524\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44546\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__44626\,
            I => \N__44541\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__44623\,
            I => \N__44541\
        );

    \I__8521\ : Span4Mux_v
    port map (
            O => \N__44620\,
            I => \N__44530\
        );

    \I__8520\ : Span4Mux_v
    port map (
            O => \N__44615\,
            I => \N__44530\
        );

    \I__8519\ : Span4Mux_h
    port map (
            O => \N__44612\,
            I => \N__44530\
        );

    \I__8518\ : Span4Mux_v
    port map (
            O => \N__44609\,
            I => \N__44530\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__44604\,
            I => \N__44530\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__44601\,
            I => \N__44523\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__44594\,
            I => \N__44523\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__44585\,
            I => \N__44523\
        );

    \I__8513\ : Odrv4
    port map (
            O => \N__44582\,
            I => \controlWord_2\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__44579\,
            I => \controlWord_2\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__44576\,
            I => \controlWord_2\
        );

    \I__8510\ : Odrv12
    port map (
            O => \N__44573\,
            I => \controlWord_2\
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__44570\,
            I => \controlWord_2\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__44565\,
            I => \controlWord_2\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__44560\,
            I => \controlWord_2\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__44549\,
            I => \controlWord_2\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__44546\,
            I => \controlWord_2\
        );

    \I__8504\ : Odrv4
    port map (
            O => \N__44541\,
            I => \controlWord_2\
        );

    \I__8503\ : Odrv4
    port map (
            O => \N__44530\,
            I => \controlWord_2\
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__44523\,
            I => \controlWord_2\
        );

    \I__8501\ : InMux
    port map (
            O => \N__44498\,
            I => \N__44490\
        );

    \I__8500\ : InMux
    port map (
            O => \N__44497\,
            I => \N__44490\
        );

    \I__8499\ : InMux
    port map (
            O => \N__44496\,
            I => \N__44485\
        );

    \I__8498\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44485\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__44490\,
            I => \N__44482\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__44485\,
            I => \N__44479\
        );

    \I__8495\ : Span12Mux_v
    port map (
            O => \N__44482\,
            I => \N__44475\
        );

    \I__8494\ : Span4Mux_v
    port map (
            O => \N__44479\,
            I => \N__44472\
        );

    \I__8493\ : InMux
    port map (
            O => \N__44478\,
            I => \N__44469\
        );

    \I__8492\ : Odrv12
    port map (
            O => \N__44475\,
            I => \PROM.ROMDATA.N_544_mux\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__44472\,
            I => \PROM.ROMDATA.N_544_mux\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__44469\,
            I => \PROM.ROMDATA.N_544_mux\
        );

    \I__8489\ : CEMux
    port map (
            O => \N__44462\,
            I => \N__44458\
        );

    \I__8488\ : CEMux
    port map (
            O => \N__44461\,
            I => \N__44454\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__44458\,
            I => \N__44449\
        );

    \I__8486\ : CEMux
    port map (
            O => \N__44457\,
            I => \N__44446\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__44454\,
            I => \N__44442\
        );

    \I__8484\ : CEMux
    port map (
            O => \N__44453\,
            I => \N__44439\
        );

    \I__8483\ : CEMux
    port map (
            O => \N__44452\,
            I => \N__44436\
        );

    \I__8482\ : Span4Mux_h
    port map (
            O => \N__44449\,
            I => \N__44429\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__44446\,
            I => \N__44429\
        );

    \I__8480\ : CEMux
    port map (
            O => \N__44445\,
            I => \N__44426\
        );

    \I__8479\ : Span4Mux_h
    port map (
            O => \N__44442\,
            I => \N__44419\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__44439\,
            I => \N__44419\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__44436\,
            I => \N__44419\
        );

    \I__8476\ : CEMux
    port map (
            O => \N__44435\,
            I => \N__44416\
        );

    \I__8475\ : CEMux
    port map (
            O => \N__44434\,
            I => \N__44412\
        );

    \I__8474\ : Span4Mux_h
    port map (
            O => \N__44429\,
            I => \N__44407\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__44426\,
            I => \N__44407\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__44419\,
            I => \N__44402\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__44416\,
            I => \N__44402\
        );

    \I__8470\ : CEMux
    port map (
            O => \N__44415\,
            I => \N__44399\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__44412\,
            I => \N__44393\
        );

    \I__8468\ : Span4Mux_v
    port map (
            O => \N__44407\,
            I => \N__44390\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__44402\,
            I => \N__44385\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__44399\,
            I => \N__44385\
        );

    \I__8465\ : CEMux
    port map (
            O => \N__44398\,
            I => \N__44382\
        );

    \I__8464\ : CEMux
    port map (
            O => \N__44397\,
            I => \N__44379\
        );

    \I__8463\ : CEMux
    port map (
            O => \N__44396\,
            I => \N__44376\
        );

    \I__8462\ : Span4Mux_h
    port map (
            O => \N__44393\,
            I => \N__44373\
        );

    \I__8461\ : Span4Mux_h
    port map (
            O => \N__44390\,
            I => \N__44370\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__44385\,
            I => \N__44365\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__44382\,
            I => \N__44365\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__44379\,
            I => \N__44362\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__44376\,
            I => \N__44359\
        );

    \I__8456\ : Span4Mux_h
    port map (
            O => \N__44373\,
            I => \N__44356\
        );

    \I__8455\ : Span4Mux_h
    port map (
            O => \N__44370\,
            I => \N__44353\
        );

    \I__8454\ : Span4Mux_h
    port map (
            O => \N__44365\,
            I => \N__44350\
        );

    \I__8453\ : Span4Mux_v
    port map (
            O => \N__44362\,
            I => \N__44345\
        );

    \I__8452\ : Span4Mux_v
    port map (
            O => \N__44359\,
            I => \N__44345\
        );

    \I__8451\ : Odrv4
    port map (
            O => \N__44356\,
            I => \CONTROL.N_35\
        );

    \I__8450\ : Odrv4
    port map (
            O => \N__44353\,
            I => \CONTROL.N_35\
        );

    \I__8449\ : Odrv4
    port map (
            O => \N__44350\,
            I => \CONTROL.N_35\
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__44345\,
            I => \CONTROL.N_35\
        );

    \I__8447\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44333\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__44333\,
            I => \N__44330\
        );

    \I__8445\ : Odrv4
    port map (
            O => \N__44330\,
            I => \PROM.ROMDATA.m444_am\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__44327\,
            I => \PROM.ROMDATA.m444_bm_cascade_\
        );

    \I__8443\ : CascadeMux
    port map (
            O => \N__44324\,
            I => \N__44321\
        );

    \I__8442\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44315\
        );

    \I__8441\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44315\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__44315\,
            I => \N__44312\
        );

    \I__8439\ : Span4Mux_h
    port map (
            O => \N__44312\,
            I => \N__44309\
        );

    \I__8438\ : Span4Mux_h
    port map (
            O => \N__44309\,
            I => \N__44304\
        );

    \I__8437\ : InMux
    port map (
            O => \N__44308\,
            I => \N__44299\
        );

    \I__8436\ : InMux
    port map (
            O => \N__44307\,
            I => \N__44299\
        );

    \I__8435\ : Odrv4
    port map (
            O => \N__44304\,
            I => \PROM.ROMDATA.m289\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__44299\,
            I => \PROM.ROMDATA.m289\
        );

    \I__8433\ : CascadeMux
    port map (
            O => \N__44294\,
            I => \N__44291\
        );

    \I__8432\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44288\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44285\
        );

    \I__8430\ : Span4Mux_v
    port map (
            O => \N__44285\,
            I => \N__44282\
        );

    \I__8429\ : Odrv4
    port map (
            O => \N__44282\,
            I => \PROM.ROMDATA.m418_ns_1\
        );

    \I__8428\ : InMux
    port map (
            O => \N__44279\,
            I => \N__44273\
        );

    \I__8427\ : InMux
    port map (
            O => \N__44278\,
            I => \N__44273\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__44273\,
            I => \N__44270\
        );

    \I__8425\ : Span4Mux_h
    port map (
            O => \N__44270\,
            I => \N__44267\
        );

    \I__8424\ : Span4Mux_h
    port map (
            O => \N__44267\,
            I => \N__44264\
        );

    \I__8423\ : Span4Mux_h
    port map (
            O => \N__44264\,
            I => \N__44261\
        );

    \I__8422\ : Odrv4
    port map (
            O => \N__44261\,
            I => \PROM_ROMDATA_dintern_19ro\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__44258\,
            I => \PROM_ROMDATA_dintern_19ro_cascade_\
        );

    \I__8420\ : InMux
    port map (
            O => \N__44255\,
            I => \N__44252\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__44252\,
            I => \N__44249\
        );

    \I__8418\ : Span12Mux_h
    port map (
            O => \N__44249\,
            I => \N__44246\
        );

    \I__8417\ : Odrv12
    port map (
            O => \N__44246\,
            I => \controlWord_19\
        );

    \I__8416\ : InMux
    port map (
            O => \N__44243\,
            I => \N__44239\
        );

    \I__8415\ : CascadeMux
    port map (
            O => \N__44242\,
            I => \N__44236\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__44239\,
            I => \N__44232\
        );

    \I__8413\ : InMux
    port map (
            O => \N__44236\,
            I => \N__44229\
        );

    \I__8412\ : CascadeMux
    port map (
            O => \N__44235\,
            I => \N__44226\
        );

    \I__8411\ : Span4Mux_v
    port map (
            O => \N__44232\,
            I => \N__44223\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__44229\,
            I => \N__44220\
        );

    \I__8409\ : InMux
    port map (
            O => \N__44226\,
            I => \N__44217\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__44223\,
            I => \N__44212\
        );

    \I__8407\ : Span4Mux_v
    port map (
            O => \N__44220\,
            I => \N__44212\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__44217\,
            I => \N__44209\
        );

    \I__8405\ : Span4Mux_v
    port map (
            O => \N__44212\,
            I => \N__44206\
        );

    \I__8404\ : Span4Mux_v
    port map (
            O => \N__44209\,
            I => \N__44203\
        );

    \I__8403\ : Sp12to4
    port map (
            O => \N__44206\,
            I => \N__44200\
        );

    \I__8402\ : Odrv4
    port map (
            O => \N__44203\,
            I => f_3
        );

    \I__8401\ : Odrv12
    port map (
            O => \N__44200\,
            I => f_3
        );

    \I__8400\ : CascadeMux
    port map (
            O => \N__44195\,
            I => \controlWord_19_cascade_\
        );

    \I__8399\ : InMux
    port map (
            O => \N__44192\,
            I => \N__44189\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__44189\,
            I => \N__44185\
        );

    \I__8397\ : InMux
    port map (
            O => \N__44188\,
            I => \N__44182\
        );

    \I__8396\ : Span4Mux_h
    port map (
            O => \N__44185\,
            I => \N__44179\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__44182\,
            I => \N__44173\
        );

    \I__8394\ : Span4Mux_h
    port map (
            O => \N__44179\,
            I => \N__44173\
        );

    \I__8393\ : InMux
    port map (
            O => \N__44178\,
            I => \N__44170\
        );

    \I__8392\ : Span4Mux_h
    port map (
            O => \N__44173\,
            I => \N__44167\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__44170\,
            I => \controlWord_20\
        );

    \I__8390\ : Odrv4
    port map (
            O => \N__44167\,
            I => \controlWord_20\
        );

    \I__8389\ : CascadeMux
    port map (
            O => \N__44162\,
            I => \N__44159\
        );

    \I__8388\ : InMux
    port map (
            O => \N__44159\,
            I => \N__44156\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__44156\,
            I => \N__44152\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__44155\,
            I => \N__44149\
        );

    \I__8385\ : Span4Mux_h
    port map (
            O => \N__44152\,
            I => \N__44146\
        );

    \I__8384\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44143\
        );

    \I__8383\ : Span4Mux_h
    port map (
            O => \N__44146\,
            I => \N__44140\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__44143\,
            I => \N__44136\
        );

    \I__8381\ : Span4Mux_v
    port map (
            O => \N__44140\,
            I => \N__44133\
        );

    \I__8380\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44130\
        );

    \I__8379\ : Span4Mux_h
    port map (
            O => \N__44136\,
            I => \N__44127\
        );

    \I__8378\ : Span4Mux_h
    port map (
            O => \N__44133\,
            I => \N__44122\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__44130\,
            I => \N__44122\
        );

    \I__8376\ : Span4Mux_h
    port map (
            O => \N__44127\,
            I => \N__44119\
        );

    \I__8375\ : Span4Mux_h
    port map (
            O => \N__44122\,
            I => \N__44116\
        );

    \I__8374\ : Odrv4
    port map (
            O => \N__44119\,
            I => f_4
        );

    \I__8373\ : Odrv4
    port map (
            O => \N__44116\,
            I => f_4
        );

    \I__8372\ : IoInMux
    port map (
            O => \N__44111\,
            I => \N__44108\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__44108\,
            I => \N__44105\
        );

    \I__8370\ : Span4Mux_s2_v
    port map (
            O => \N__44105\,
            I => \N__44102\
        );

    \I__8369\ : Span4Mux_h
    port map (
            O => \N__44102\,
            I => \N__44098\
        );

    \I__8368\ : InMux
    port map (
            O => \N__44101\,
            I => \N__44095\
        );

    \I__8367\ : Span4Mux_h
    port map (
            O => \N__44098\,
            I => \N__44092\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__44095\,
            I => \N__44089\
        );

    \I__8365\ : Span4Mux_h
    port map (
            O => \N__44092\,
            I => \N__44086\
        );

    \I__8364\ : Span4Mux_v
    port map (
            O => \N__44089\,
            I => \N__44083\
        );

    \I__8363\ : Span4Mux_v
    port map (
            O => \N__44086\,
            I => \N__44078\
        );

    \I__8362\ : Span4Mux_v
    port map (
            O => \N__44083\,
            I => \N__44078\
        );

    \I__8361\ : Span4Mux_h
    port map (
            O => \N__44078\,
            I => \N__44075\
        );

    \I__8360\ : Odrv4
    port map (
            O => \N__44075\,
            I => \A14_c\
        );

    \I__8359\ : IoInMux
    port map (
            O => \N__44072\,
            I => \N__44069\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__44069\,
            I => \N__44066\
        );

    \I__8357\ : Span4Mux_s2_h
    port map (
            O => \N__44066\,
            I => \N__44063\
        );

    \I__8356\ : Span4Mux_v
    port map (
            O => \N__44063\,
            I => \N__44060\
        );

    \I__8355\ : Sp12to4
    port map (
            O => \N__44060\,
            I => \N__44056\
        );

    \I__8354\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44053\
        );

    \I__8353\ : Odrv12
    port map (
            O => \N__44056\,
            I => \A4_c\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__44053\,
            I => \A4_c\
        );

    \I__8351\ : IoInMux
    port map (
            O => \N__44048\,
            I => \N__44045\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__44045\,
            I => \N__44042\
        );

    \I__8349\ : Span4Mux_s1_h
    port map (
            O => \N__44042\,
            I => \N__44039\
        );

    \I__8348\ : Sp12to4
    port map (
            O => \N__44039\,
            I => \N__44036\
        );

    \I__8347\ : Span12Mux_v
    port map (
            O => \N__44036\,
            I => \N__44033\
        );

    \I__8346\ : Span12Mux_h
    port map (
            O => \N__44033\,
            I => \N__44029\
        );

    \I__8345\ : InMux
    port map (
            O => \N__44032\,
            I => \N__44026\
        );

    \I__8344\ : Odrv12
    port map (
            O => \N__44029\,
            I => \A3_c\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__44026\,
            I => \A3_c\
        );

    \I__8342\ : InMux
    port map (
            O => \N__44021\,
            I => \N__44018\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__44018\,
            I => \N__44015\
        );

    \I__8340\ : Span4Mux_h
    port map (
            O => \N__44015\,
            I => \N__44012\
        );

    \I__8339\ : Span4Mux_v
    port map (
            O => \N__44012\,
            I => \N__44009\
        );

    \I__8338\ : Sp12to4
    port map (
            O => \N__44009\,
            I => \N__44006\
        );

    \I__8337\ : Span12Mux_h
    port map (
            O => \N__44006\,
            I => \N__44003\
        );

    \I__8336\ : Odrv12
    port map (
            O => \N__44003\,
            I => \RAM.un1_WR_105_0Z0Z_7\
        );

    \I__8335\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43992\
        );

    \I__8334\ : InMux
    port map (
            O => \N__43999\,
            I => \N__43992\
        );

    \I__8333\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43987\
        );

    \I__8332\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43987\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__43992\,
            I => \N__43984\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__43987\,
            I => \N__43976\
        );

    \I__8329\ : Span4Mux_h
    port map (
            O => \N__43984\,
            I => \N__43971\
        );

    \I__8328\ : InMux
    port map (
            O => \N__43983\,
            I => \N__43964\
        );

    \I__8327\ : InMux
    port map (
            O => \N__43982\,
            I => \N__43964\
        );

    \I__8326\ : InMux
    port map (
            O => \N__43981\,
            I => \N__43964\
        );

    \I__8325\ : InMux
    port map (
            O => \N__43980\,
            I => \N__43959\
        );

    \I__8324\ : InMux
    port map (
            O => \N__43979\,
            I => \N__43959\
        );

    \I__8323\ : Span4Mux_h
    port map (
            O => \N__43976\,
            I => \N__43956\
        );

    \I__8322\ : InMux
    port map (
            O => \N__43975\,
            I => \N__43951\
        );

    \I__8321\ : InMux
    port map (
            O => \N__43974\,
            I => \N__43951\
        );

    \I__8320\ : Span4Mux_h
    port map (
            O => \N__43971\,
            I => \N__43948\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__43964\,
            I => \aluOperand2_2_rep1\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__43959\,
            I => \aluOperand2_2_rep1\
        );

    \I__8317\ : Odrv4
    port map (
            O => \N__43956\,
            I => \aluOperand2_2_rep1\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__43951\,
            I => \aluOperand2_2_rep1\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__43948\,
            I => \aluOperand2_2_rep1\
        );

    \I__8314\ : InMux
    port map (
            O => \N__43937\,
            I => \N__43934\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__43934\,
            I => \ALU.operand2_3_ns_1_7\
        );

    \I__8312\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43925\
        );

    \I__8311\ : InMux
    port map (
            O => \N__43930\,
            I => \N__43925\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__43925\,
            I => \N__43922\
        );

    \I__8309\ : Span4Mux_h
    port map (
            O => \N__43922\,
            I => \N__43909\
        );

    \I__8308\ : InMux
    port map (
            O => \N__43921\,
            I => \N__43904\
        );

    \I__8307\ : InMux
    port map (
            O => \N__43920\,
            I => \N__43904\
        );

    \I__8306\ : InMux
    port map (
            O => \N__43919\,
            I => \N__43898\
        );

    \I__8305\ : InMux
    port map (
            O => \N__43918\,
            I => \N__43898\
        );

    \I__8304\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43891\
        );

    \I__8303\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43891\
        );

    \I__8302\ : InMux
    port map (
            O => \N__43915\,
            I => \N__43886\
        );

    \I__8301\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43886\
        );

    \I__8300\ : InMux
    port map (
            O => \N__43913\,
            I => \N__43881\
        );

    \I__8299\ : InMux
    port map (
            O => \N__43912\,
            I => \N__43881\
        );

    \I__8298\ : Span4Mux_h
    port map (
            O => \N__43909\,
            I => \N__43878\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__43904\,
            I => \N__43875\
        );

    \I__8296\ : InMux
    port map (
            O => \N__43903\,
            I => \N__43872\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__43898\,
            I => \N__43869\
        );

    \I__8294\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43866\
        );

    \I__8293\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43863\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__43891\,
            I => \N__43858\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__43886\,
            I => \N__43858\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__43881\,
            I => \N__43853\
        );

    \I__8289\ : Span4Mux_v
    port map (
            O => \N__43878\,
            I => \N__43853\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__43875\,
            I => \N__43850\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__43872\,
            I => \aluOperand1_1_rep1\
        );

    \I__8286\ : Odrv4
    port map (
            O => \N__43869\,
            I => \aluOperand1_1_rep1\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__43866\,
            I => \aluOperand1_1_rep1\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__43863\,
            I => \aluOperand1_1_rep1\
        );

    \I__8283\ : Odrv12
    port map (
            O => \N__43858\,
            I => \aluOperand1_1_rep1\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__43853\,
            I => \aluOperand1_1_rep1\
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__43850\,
            I => \aluOperand1_1_rep1\
        );

    \I__8280\ : InMux
    port map (
            O => \N__43835\,
            I => \N__43832\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__43832\,
            I => \N__43829\
        );

    \I__8278\ : Span4Mux_v
    port map (
            O => \N__43829\,
            I => \N__43826\
        );

    \I__8277\ : Span4Mux_v
    port map (
            O => \N__43826\,
            I => \N__43823\
        );

    \I__8276\ : Sp12to4
    port map (
            O => \N__43823\,
            I => \N__43819\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__43822\,
            I => \N__43816\
        );

    \I__8274\ : Span12Mux_h
    port map (
            O => \N__43819\,
            I => \N__43812\
        );

    \I__8273\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43809\
        );

    \I__8272\ : InMux
    port map (
            O => \N__43815\,
            I => \N__43806\
        );

    \I__8271\ : Odrv12
    port map (
            O => \N__43812\,
            I => h_7
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__43809\,
            I => h_7
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__43806\,
            I => h_7
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__43799\,
            I => \ALU.dout_6_ns_1_7_cascade_\
        );

    \I__8267\ : CascadeMux
    port map (
            O => \N__43796\,
            I => \ALU.N_1140_cascade_\
        );

    \I__8266\ : InMux
    port map (
            O => \N__43793\,
            I => \N__43790\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__43790\,
            I => \ALU.N_1092\
        );

    \I__8264\ : InMux
    port map (
            O => \N__43787\,
            I => \N__43784\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__43784\,
            I => \N__43781\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__43781\,
            I => \N__43778\
        );

    \I__8261\ : Span4Mux_h
    port map (
            O => \N__43778\,
            I => \N__43775\
        );

    \I__8260\ : Odrv4
    port map (
            O => \N__43775\,
            I => \DROM_ROMDATA_dintern_7ro\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__43772\,
            I => \aluOut_7_cascade_\
        );

    \I__8258\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43766\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__43766\,
            I => \N__43763\
        );

    \I__8256\ : Span4Mux_h
    port map (
            O => \N__43763\,
            I => \N__43760\
        );

    \I__8255\ : Span4Mux_h
    port map (
            O => \N__43760\,
            I => \N__43756\
        );

    \I__8254\ : InMux
    port map (
            O => \N__43759\,
            I => \N__43753\
        );

    \I__8253\ : Odrv4
    port map (
            O => \N__43756\,
            I => \N_200\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__43753\,
            I => \N_200\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__43748\,
            I => \PROM.ROMDATA.m267_cascade_\
        );

    \I__8250\ : CascadeMux
    port map (
            O => \N__43745\,
            I => \N__43741\
        );

    \I__8249\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43736\
        );

    \I__8248\ : InMux
    port map (
            O => \N__43741\,
            I => \N__43736\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__43736\,
            I => \N__43733\
        );

    \I__8246\ : Span4Mux_v
    port map (
            O => \N__43733\,
            I => \N__43730\
        );

    \I__8245\ : Sp12to4
    port map (
            O => \N__43730\,
            I => \N__43727\
        );

    \I__8244\ : Span12Mux_h
    port map (
            O => \N__43727\,
            I => \N__43724\
        );

    \I__8243\ : Odrv12
    port map (
            O => \N__43724\,
            I => \PROM.ROMDATA.m442\
        );

    \I__8242\ : InMux
    port map (
            O => \N__43721\,
            I => \N__43718\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__43718\,
            I => \N__43715\
        );

    \I__8240\ : Span12Mux_h
    port map (
            O => \N__43715\,
            I => \N__43711\
        );

    \I__8239\ : InMux
    port map (
            O => \N__43714\,
            I => \N__43708\
        );

    \I__8238\ : Odrv12
    port map (
            O => \N__43711\,
            I => \PROM.ROMDATA.m282\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__43708\,
            I => \PROM.ROMDATA.m282\
        );

    \I__8236\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43700\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__43700\,
            I => \N__43697\
        );

    \I__8234\ : Span4Mux_h
    port map (
            O => \N__43697\,
            I => \N__43694\
        );

    \I__8233\ : Span4Mux_h
    port map (
            O => \N__43694\,
            I => \N__43691\
        );

    \I__8232\ : Span4Mux_h
    port map (
            O => \N__43691\,
            I => \N__43687\
        );

    \I__8231\ : InMux
    port map (
            O => \N__43690\,
            I => \N__43684\
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__43687\,
            I => \PROM.ROMDATA.dintern_29dfltZ0Z_1\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__43684\,
            I => \PROM.ROMDATA.dintern_29dfltZ0Z_1\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__43679\,
            I => \PROM.ROMDATA.m282_cascade_\
        );

    \I__8227\ : InMux
    port map (
            O => \N__43676\,
            I => \N__43673\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__43673\,
            I => \N__43670\
        );

    \I__8225\ : Span4Mux_v
    port map (
            O => \N__43670\,
            I => \N__43666\
        );

    \I__8224\ : InMux
    port map (
            O => \N__43669\,
            I => \N__43663\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__43666\,
            I => \N__43658\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__43663\,
            I => \N__43658\
        );

    \I__8221\ : Span4Mux_v
    port map (
            O => \N__43658\,
            I => \N__43655\
        );

    \I__8220\ : Span4Mux_h
    port map (
            O => \N__43655\,
            I => \N__43652\
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__43652\,
            I => \CONTROL.ctrlOut_13\
        );

    \I__8218\ : CascadeMux
    port map (
            O => \N__43649\,
            I => \ALU.N_1252_cascade_\
        );

    \I__8217\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43643\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__43643\,
            I => \ALU.N_1204\
        );

    \I__8215\ : CascadeMux
    port map (
            O => \N__43640\,
            I => \ALU.d_RNIO5IF4Z0Z_7_cascade_\
        );

    \I__8214\ : InMux
    port map (
            O => \N__43637\,
            I => \N__43634\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__43634\,
            I => \N__43631\
        );

    \I__8212\ : Span4Mux_h
    port map (
            O => \N__43631\,
            I => \N__43628\
        );

    \I__8211\ : Span4Mux_h
    port map (
            O => \N__43628\,
            I => \N__43625\
        );

    \I__8210\ : Odrv4
    port map (
            O => \N__43625\,
            I => \ALU.combOperand2_d_bmZ0Z_7\
        );

    \I__8209\ : CascadeMux
    port map (
            O => \N__43622\,
            I => \ALU.d_RNIM3JB6Z0Z_7_cascade_\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__43619\,
            I => \ALU.dout_3_ns_1_7_cascade_\
        );

    \I__8207\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__43613\,
            I => \ALU.operand2_6_ns_1_7\
        );

    \I__8205\ : InMux
    port map (
            O => \N__43610\,
            I => \N__43607\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__43607\,
            I => \ALU.N_606\
        );

    \I__8203\ : CascadeMux
    port map (
            O => \N__43604\,
            I => \N__43600\
        );

    \I__8202\ : InMux
    port map (
            O => \N__43603\,
            I => \N__43596\
        );

    \I__8201\ : InMux
    port map (
            O => \N__43600\,
            I => \N__43591\
        );

    \I__8200\ : InMux
    port map (
            O => \N__43599\,
            I => \N__43591\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__43596\,
            I => \N__43585\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__43591\,
            I => \N__43585\
        );

    \I__8197\ : InMux
    port map (
            O => \N__43590\,
            I => \N__43582\
        );

    \I__8196\ : Span4Mux_h
    port map (
            O => \N__43585\,
            I => \N__43579\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__43582\,
            I => \ALU.N_638\
        );

    \I__8194\ : Odrv4
    port map (
            O => \N__43579\,
            I => \ALU.N_638\
        );

    \I__8193\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43568\
        );

    \I__8192\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43568\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__43568\,
            I => \N__43565\
        );

    \I__8190\ : Span4Mux_v
    port map (
            O => \N__43565\,
            I => \N__43562\
        );

    \I__8189\ : Span4Mux_h
    port map (
            O => \N__43562\,
            I => \N__43559\
        );

    \I__8188\ : Odrv4
    port map (
            O => \N__43559\,
            I => \ALU.a_15_m0_amZ0Z_2\
        );

    \I__8187\ : CascadeMux
    port map (
            O => \N__43556\,
            I => \ALU.a_15_m1_9_cascade_\
        );

    \I__8186\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43549\
        );

    \I__8185\ : InMux
    port map (
            O => \N__43552\,
            I => \N__43546\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__43549\,
            I => \N__43543\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__43546\,
            I => \N__43540\
        );

    \I__8182\ : Span4Mux_h
    port map (
            O => \N__43543\,
            I => \N__43535\
        );

    \I__8181\ : Span4Mux_v
    port map (
            O => \N__43540\,
            I => \N__43535\
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__43535\,
            I => \ALU.aZ0Z_9\
        );

    \I__8179\ : InMux
    port map (
            O => \N__43532\,
            I => \N__43526\
        );

    \I__8178\ : InMux
    port map (
            O => \N__43531\,
            I => \N__43526\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__43526\,
            I => \N__43523\
        );

    \I__8176\ : Span4Mux_h
    port map (
            O => \N__43523\,
            I => \N__43520\
        );

    \I__8175\ : Span4Mux_h
    port map (
            O => \N__43520\,
            I => \N__43517\
        );

    \I__8174\ : Span4Mux_h
    port map (
            O => \N__43517\,
            I => \N__43514\
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__43514\,
            I => \N_227_0\
        );

    \I__8172\ : CascadeMux
    port map (
            O => \N__43511\,
            I => \N__43508\
        );

    \I__8171\ : InMux
    port map (
            O => \N__43508\,
            I => \N__43502\
        );

    \I__8170\ : InMux
    port map (
            O => \N__43507\,
            I => \N__43502\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__43502\,
            I => \N__43499\
        );

    \I__8168\ : Span4Mux_v
    port map (
            O => \N__43499\,
            I => \N__43496\
        );

    \I__8167\ : Span4Mux_h
    port map (
            O => \N__43496\,
            I => \N__43491\
        );

    \I__8166\ : InMux
    port map (
            O => \N__43495\,
            I => \N__43486\
        );

    \I__8165\ : InMux
    port map (
            O => \N__43494\,
            I => \N__43486\
        );

    \I__8164\ : Odrv4
    port map (
            O => \N__43491\,
            I => \N_179\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__43486\,
            I => \N_179\
        );

    \I__8162\ : IoInMux
    port map (
            O => \N__43481\,
            I => \N__43478\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__43478\,
            I => \N__43475\
        );

    \I__8160\ : IoSpan4Mux
    port map (
            O => \N__43475\,
            I => \N__43471\
        );

    \I__8159\ : IoInMux
    port map (
            O => \N__43474\,
            I => \N__43468\
        );

    \I__8158\ : Span4Mux_s3_h
    port map (
            O => \N__43471\,
            I => \N__43465\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__43468\,
            I => \N__43462\
        );

    \I__8156\ : Sp12to4
    port map (
            O => \N__43465\,
            I => \N__43459\
        );

    \I__8155\ : Span12Mux_s6_h
    port map (
            O => \N__43462\,
            I => \N__43456\
        );

    \I__8154\ : Span12Mux_h
    port map (
            O => \N__43459\,
            I => \N__43451\
        );

    \I__8153\ : Span12Mux_h
    port map (
            O => \N__43456\,
            I => \N__43451\
        );

    \I__8152\ : Odrv12
    port map (
            O => \N__43451\,
            I => bus_2
        );

    \I__8151\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43445\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__43445\,
            I => \N__43441\
        );

    \I__8149\ : InMux
    port map (
            O => \N__43444\,
            I => \N__43438\
        );

    \I__8148\ : Span12Mux_h
    port map (
            O => \N__43441\,
            I => \N__43435\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__43438\,
            I => \ALU.bZ0Z_4\
        );

    \I__8146\ : Odrv12
    port map (
            O => \N__43435\,
            I => \ALU.bZ0Z_4\
        );

    \I__8145\ : InMux
    port map (
            O => \N__43430\,
            I => \N__43427\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__43427\,
            I => \N__43424\
        );

    \I__8143\ : Span4Mux_h
    port map (
            O => \N__43424\,
            I => \N__43421\
        );

    \I__8142\ : Span4Mux_h
    port map (
            O => \N__43421\,
            I => \N__43418\
        );

    \I__8141\ : Odrv4
    port map (
            O => \N__43418\,
            I => \ALU.b_RNI5FSPZ0Z_4\
        );

    \I__8140\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43412\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__43412\,
            I => \N__43409\
        );

    \I__8138\ : Span4Mux_h
    port map (
            O => \N__43409\,
            I => \N__43406\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__43406\,
            I => \ALU.c_RNIHV2SZ0Z_9\
        );

    \I__8136\ : CascadeMux
    port map (
            O => \N__43403\,
            I => \N__43399\
        );

    \I__8135\ : InMux
    port map (
            O => \N__43402\,
            I => \N__43396\
        );

    \I__8134\ : InMux
    port map (
            O => \N__43399\,
            I => \N__43393\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__43396\,
            I => \N__43390\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__43393\,
            I => \N__43387\
        );

    \I__8131\ : Span4Mux_v
    port map (
            O => \N__43390\,
            I => \N__43383\
        );

    \I__8130\ : Span4Mux_v
    port map (
            O => \N__43387\,
            I => \N__43380\
        );

    \I__8129\ : InMux
    port map (
            O => \N__43386\,
            I => \N__43377\
        );

    \I__8128\ : Span4Mux_v
    port map (
            O => \N__43383\,
            I => \N__43374\
        );

    \I__8127\ : Span4Mux_v
    port map (
            O => \N__43380\,
            I => \N__43371\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__43377\,
            I => \N__43368\
        );

    \I__8125\ : Span4Mux_h
    port map (
            O => \N__43374\,
            I => \N__43365\
        );

    \I__8124\ : Span4Mux_h
    port map (
            O => \N__43371\,
            I => \N__43362\
        );

    \I__8123\ : Span4Mux_v
    port map (
            O => \N__43368\,
            I => \N__43359\
        );

    \I__8122\ : Sp12to4
    port map (
            O => \N__43365\,
            I => \N__43356\
        );

    \I__8121\ : Odrv4
    port map (
            O => \N__43362\,
            I => h_4
        );

    \I__8120\ : Odrv4
    port map (
            O => \N__43359\,
            I => h_4
        );

    \I__8119\ : Odrv12
    port map (
            O => \N__43356\,
            I => h_4
        );

    \I__8118\ : InMux
    port map (
            O => \N__43349\,
            I => \N__43345\
        );

    \I__8117\ : InMux
    port map (
            O => \N__43348\,
            I => \N__43342\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__43345\,
            I => \N__43339\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__43342\,
            I => \N__43336\
        );

    \I__8114\ : Span4Mux_h
    port map (
            O => \N__43339\,
            I => \N__43331\
        );

    \I__8113\ : Span4Mux_v
    port map (
            O => \N__43336\,
            I => \N__43331\
        );

    \I__8112\ : Span4Mux_h
    port map (
            O => \N__43331\,
            I => \N__43328\
        );

    \I__8111\ : Odrv4
    port map (
            O => \N__43328\,
            I => \ALU.dZ0Z_4\
        );

    \I__8110\ : InMux
    port map (
            O => \N__43325\,
            I => \N__43322\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__43322\,
            I => \N__43319\
        );

    \I__8108\ : Span4Mux_h
    port map (
            O => \N__43319\,
            I => \N__43316\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__43316\,
            I => \N__43313\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__43313\,
            I => \ALU.d_RNI9R8EZ0Z_4\
        );

    \I__8105\ : InMux
    port map (
            O => \N__43310\,
            I => \N__43300\
        );

    \I__8104\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43297\
        );

    \I__8103\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43288\
        );

    \I__8102\ : InMux
    port map (
            O => \N__43307\,
            I => \N__43288\
        );

    \I__8101\ : InMux
    port map (
            O => \N__43306\,
            I => \N__43280\
        );

    \I__8100\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43280\
        );

    \I__8099\ : InMux
    port map (
            O => \N__43304\,
            I => \N__43280\
        );

    \I__8098\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43274\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__43300\,
            I => \N__43269\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__43297\,
            I => \N__43269\
        );

    \I__8095\ : InMux
    port map (
            O => \N__43296\,
            I => \N__43260\
        );

    \I__8094\ : InMux
    port map (
            O => \N__43295\,
            I => \N__43260\
        );

    \I__8093\ : InMux
    port map (
            O => \N__43294\,
            I => \N__43260\
        );

    \I__8092\ : InMux
    port map (
            O => \N__43293\,
            I => \N__43260\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__43288\,
            I => \N__43257\
        );

    \I__8090\ : InMux
    port map (
            O => \N__43287\,
            I => \N__43254\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__43280\,
            I => \N__43251\
        );

    \I__8088\ : InMux
    port map (
            O => \N__43279\,
            I => \N__43244\
        );

    \I__8087\ : InMux
    port map (
            O => \N__43278\,
            I => \N__43244\
        );

    \I__8086\ : InMux
    port map (
            O => \N__43277\,
            I => \N__43244\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__43274\,
            I => \N__43239\
        );

    \I__8084\ : Span4Mux_v
    port map (
            O => \N__43269\,
            I => \N__43234\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__43260\,
            I => \N__43231\
        );

    \I__8082\ : Span4Mux_v
    port map (
            O => \N__43257\,
            I => \N__43222\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__43254\,
            I => \N__43222\
        );

    \I__8080\ : Span4Mux_v
    port map (
            O => \N__43251\,
            I => \N__43222\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__43244\,
            I => \N__43222\
        );

    \I__8078\ : InMux
    port map (
            O => \N__43243\,
            I => \N__43217\
        );

    \I__8077\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43217\
        );

    \I__8076\ : Span4Mux_v
    port map (
            O => \N__43239\,
            I => \N__43214\
        );

    \I__8075\ : InMux
    port map (
            O => \N__43238\,
            I => \N__43209\
        );

    \I__8074\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43209\
        );

    \I__8073\ : Span4Mux_h
    port map (
            O => \N__43234\,
            I => \N__43206\
        );

    \I__8072\ : Span4Mux_v
    port map (
            O => \N__43231\,
            I => \N__43201\
        );

    \I__8071\ : Span4Mux_h
    port map (
            O => \N__43222\,
            I => \N__43201\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__43217\,
            I => \N__43198\
        );

    \I__8069\ : Odrv4
    port map (
            O => \N__43214\,
            I => \aluOperand2_2\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__43209\,
            I => \aluOperand2_2\
        );

    \I__8067\ : Odrv4
    port map (
            O => \N__43206\,
            I => \aluOperand2_2\
        );

    \I__8066\ : Odrv4
    port map (
            O => \N__43201\,
            I => \aluOperand2_2\
        );

    \I__8065\ : Odrv4
    port map (
            O => \N__43198\,
            I => \aluOperand2_2\
        );

    \I__8064\ : CascadeMux
    port map (
            O => \N__43187\,
            I => \ALU.N_852_cascade_\
        );

    \I__8063\ : InMux
    port map (
            O => \N__43184\,
            I => \N__43180\
        );

    \I__8062\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43177\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43174\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__43177\,
            I => \ALU.N_966\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__43174\,
            I => \ALU.N_966\
        );

    \I__8058\ : CascadeMux
    port map (
            O => \N__43169\,
            I => \ALU.N_766_cascade_\
        );

    \I__8057\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43161\
        );

    \I__8056\ : CascadeMux
    port map (
            O => \N__43165\,
            I => \N__43157\
        );

    \I__8055\ : CascadeMux
    port map (
            O => \N__43164\,
            I => \N__43154\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__43161\,
            I => \N__43151\
        );

    \I__8053\ : InMux
    port map (
            O => \N__43160\,
            I => \N__43146\
        );

    \I__8052\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43146\
        );

    \I__8051\ : InMux
    port map (
            O => \N__43154\,
            I => \N__43143\
        );

    \I__8050\ : Span12Mux_h
    port map (
            O => \N__43151\,
            I => \N__43140\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__43146\,
            I => \N__43137\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__43143\,
            I => \N__43134\
        );

    \I__8047\ : Odrv12
    port map (
            O => \N__43140\,
            I => \ALU.N_634\
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__43137\,
            I => \ALU.N_634\
        );

    \I__8045\ : Odrv12
    port map (
            O => \N__43134\,
            I => \ALU.N_634\
        );

    \I__8044\ : CascadeMux
    port map (
            O => \N__43127\,
            I => \ALU.N_634_cascade_\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__43124\,
            I => \ALU.N_811_cascade_\
        );

    \I__8042\ : InMux
    port map (
            O => \N__43121\,
            I => \N__43115\
        );

    \I__8041\ : InMux
    port map (
            O => \N__43120\,
            I => \N__43112\
        );

    \I__8040\ : InMux
    port map (
            O => \N__43119\,
            I => \N__43109\
        );

    \I__8039\ : InMux
    port map (
            O => \N__43118\,
            I => \N__43106\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__43115\,
            I => \N__43101\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__43112\,
            I => \N__43096\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__43109\,
            I => \N__43096\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__43106\,
            I => \N__43093\
        );

    \I__8034\ : InMux
    port map (
            O => \N__43105\,
            I => \N__43090\
        );

    \I__8033\ : InMux
    port map (
            O => \N__43104\,
            I => \N__43087\
        );

    \I__8032\ : Span4Mux_h
    port map (
            O => \N__43101\,
            I => \N__43075\
        );

    \I__8031\ : Span4Mux_v
    port map (
            O => \N__43096\,
            I => \N__43075\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__43093\,
            I => \N__43075\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__43090\,
            I => \N__43075\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__43087\,
            I => \N__43075\
        );

    \I__8027\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43072\
        );

    \I__8026\ : Odrv4
    port map (
            O => \N__43075\,
            I => \ALU.d_RNIK8M6K5Z0Z_6\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__43072\,
            I => \ALU.d_RNIK8M6K5Z0Z_6\
        );

    \I__8024\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43062\
        );

    \I__8023\ : InMux
    port map (
            O => \N__43066\,
            I => \N__43059\
        );

    \I__8022\ : InMux
    port map (
            O => \N__43065\,
            I => \N__43056\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__43062\,
            I => \N__43052\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__43059\,
            I => \N__43048\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__43056\,
            I => \N__43045\
        );

    \I__8018\ : InMux
    port map (
            O => \N__43055\,
            I => \N__43042\
        );

    \I__8017\ : Span4Mux_h
    port map (
            O => \N__43052\,
            I => \N__43034\
        );

    \I__8016\ : InMux
    port map (
            O => \N__43051\,
            I => \N__43031\
        );

    \I__8015\ : Span4Mux_v
    port map (
            O => \N__43048\,
            I => \N__43024\
        );

    \I__8014\ : Span4Mux_v
    port map (
            O => \N__43045\,
            I => \N__43024\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__43042\,
            I => \N__43024\
        );

    \I__8012\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43021\
        );

    \I__8011\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43018\
        );

    \I__8010\ : InMux
    port map (
            O => \N__43039\,
            I => \N__43015\
        );

    \I__8009\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43010\
        );

    \I__8008\ : InMux
    port map (
            O => \N__43037\,
            I => \N__43010\
        );

    \I__8007\ : Odrv4
    port map (
            O => \N__43034\,
            I => \ALU.a_15_sZ0Z_11\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__43031\,
            I => \ALU.a_15_sZ0Z_11\
        );

    \I__8005\ : Odrv4
    port map (
            O => \N__43024\,
            I => \ALU.a_15_sZ0Z_11\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__43021\,
            I => \ALU.a_15_sZ0Z_11\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__43018\,
            I => \ALU.a_15_sZ0Z_11\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__43015\,
            I => \ALU.a_15_sZ0Z_11\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__43010\,
            I => \ALU.a_15_sZ0Z_11\
        );

    \I__8000\ : CascadeMux
    port map (
            O => \N__42995\,
            I => \ALU.d_RNIK8M6K5Z0Z_6_cascade_\
        );

    \I__7999\ : InMux
    port map (
            O => \N__42992\,
            I => \N__42987\
        );

    \I__7998\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42984\
        );

    \I__7997\ : InMux
    port map (
            O => \N__42990\,
            I => \N__42979\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__42987\,
            I => \N__42974\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__42984\,
            I => \N__42971\
        );

    \I__7994\ : InMux
    port map (
            O => \N__42983\,
            I => \N__42968\
        );

    \I__7993\ : InMux
    port map (
            O => \N__42982\,
            I => \N__42965\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__42979\,
            I => \N__42962\
        );

    \I__7991\ : InMux
    port map (
            O => \N__42978\,
            I => \N__42959\
        );

    \I__7990\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42956\
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__42974\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0\
        );

    \I__7988\ : Odrv4
    port map (
            O => \N__42971\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__42968\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__42965\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0\
        );

    \I__7985\ : Odrv12
    port map (
            O => \N__42962\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__42959\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__42956\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0\
        );

    \I__7982\ : InMux
    port map (
            O => \N__42941\,
            I => \N__42938\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__42938\,
            I => \N__42934\
        );

    \I__7980\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42931\
        );

    \I__7979\ : Span4Mux_v
    port map (
            O => \N__42934\,
            I => \N__42928\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__42931\,
            I => \N__42925\
        );

    \I__7977\ : Span4Mux_h
    port map (
            O => \N__42928\,
            I => \N__42922\
        );

    \I__7976\ : Span4Mux_v
    port map (
            O => \N__42925\,
            I => \N__42919\
        );

    \I__7975\ : Span4Mux_h
    port map (
            O => \N__42922\,
            I => \N__42916\
        );

    \I__7974\ : Span4Mux_h
    port map (
            O => \N__42919\,
            I => \N__42913\
        );

    \I__7973\ : Odrv4
    port map (
            O => \N__42916\,
            I => \ALU.aZ0Z_6\
        );

    \I__7972\ : Odrv4
    port map (
            O => \N__42913\,
            I => \ALU.aZ0Z_6\
        );

    \I__7971\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42905\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__42905\,
            I => \ALU.N_766\
        );

    \I__7969\ : CascadeMux
    port map (
            O => \N__42902\,
            I => \ALU.N_606_cascade_\
        );

    \I__7968\ : InMux
    port map (
            O => \N__42899\,
            I => \N__42896\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__42896\,
            I => \N__42893\
        );

    \I__7966\ : Span4Mux_h
    port map (
            O => \N__42893\,
            I => \N__42890\
        );

    \I__7965\ : Odrv4
    port map (
            O => \N__42890\,
            I => \ALU.addsub_axb_1_1\
        );

    \I__7964\ : InMux
    port map (
            O => \N__42887\,
            I => \N__42884\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__42884\,
            I => \ALU.N_1026\
        );

    \I__7962\ : InMux
    port map (
            O => \N__42881\,
            I => \N__42878\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__42878\,
            I => \N__42875\
        );

    \I__7960\ : Odrv4
    port map (
            O => \N__42875\,
            I => \ALU.mult_293_c_RNOZ0Z_0\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__7958\ : InMux
    port map (
            O => \N__42869\,
            I => \N__42865\
        );

    \I__7957\ : InMux
    port map (
            O => \N__42868\,
            I => \N__42862\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__42865\,
            I => \N__42859\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__42862\,
            I => \ALU.N_1011\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__42859\,
            I => \ALU.N_1011\
        );

    \I__7953\ : InMux
    port map (
            O => \N__42854\,
            I => \N__42851\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__42851\,
            I => \ALU.mult_323_c_RNIAA0BZ0Z82\
        );

    \I__7951\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42845\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__42845\,
            I => \ALU.d_RNIGD2441Z0Z_8\
        );

    \I__7949\ : CascadeMux
    port map (
            O => \N__42842\,
            I => \ALU.N_639_cascade_\
        );

    \I__7948\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42836\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__42836\,
            I => \N__42833\
        );

    \I__7946\ : Span4Mux_v
    port map (
            O => \N__42833\,
            I => \N__42830\
        );

    \I__7945\ : Sp12to4
    port map (
            O => \N__42830\,
            I => \N__42827\
        );

    \I__7944\ : Odrv12
    port map (
            O => \N__42827\,
            I => \ALU.d_RNIC6EBM2Z0Z_2\
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__42824\,
            I => \ALU.d_RNIFVCT15Z0Z_8_cascade_\
        );

    \I__7942\ : InMux
    port map (
            O => \N__42821\,
            I => \N__42818\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__42818\,
            I => \ALU.lshift_11\
        );

    \I__7940\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42812\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__42812\,
            I => \N__42807\
        );

    \I__7938\ : InMux
    port map (
            O => \N__42811\,
            I => \N__42802\
        );

    \I__7937\ : InMux
    port map (
            O => \N__42810\,
            I => \N__42802\
        );

    \I__7936\ : Odrv4
    port map (
            O => \N__42807\,
            I => \ALU.N_851\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__42802\,
            I => \ALU.N_851\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__42797\,
            I => \ALU.N_851_cascade_\
        );

    \I__7933\ : InMux
    port map (
            O => \N__42794\,
            I => \N__42791\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__42791\,
            I => \ALU.c_RNINT9PO2_0Z0Z_10\
        );

    \I__7931\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42782\
        );

    \I__7930\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42782\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__42782\,
            I => \ALU.N_978\
        );

    \I__7928\ : CascadeMux
    port map (
            O => \N__42779\,
            I => \ALU.N_978_cascade_\
        );

    \I__7927\ : InMux
    port map (
            O => \N__42776\,
            I => \N__42773\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__42773\,
            I => \N__42769\
        );

    \I__7925\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42766\
        );

    \I__7924\ : Span4Mux_h
    port map (
            O => \N__42769\,
            I => \N__42763\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__42766\,
            I => \N__42758\
        );

    \I__7922\ : Span4Mux_h
    port map (
            O => \N__42763\,
            I => \N__42758\
        );

    \I__7921\ : Odrv4
    port map (
            O => \N__42758\,
            I => \ALU.N_836\
        );

    \I__7920\ : CascadeMux
    port map (
            O => \N__42755\,
            I => \N__42752\
        );

    \I__7919\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42749\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__42749\,
            I => \N__42746\
        );

    \I__7917\ : Span4Mux_v
    port map (
            O => \N__42746\,
            I => \N__42743\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__42743\,
            I => \ALU.mult_293_c_RNOZ0\
        );

    \I__7915\ : InMux
    port map (
            O => \N__42740\,
            I => \N__42737\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__42737\,
            I => \N__42734\
        );

    \I__7913\ : Span4Mux_v
    port map (
            O => \N__42734\,
            I => \N__42731\
        );

    \I__7912\ : Odrv4
    port map (
            O => \N__42731\,
            I => \ALU.d_RNI34ECOZ0Z_9\
        );

    \I__7911\ : CascadeMux
    port map (
            O => \N__42728\,
            I => \N__42725\
        );

    \I__7910\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42722\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__42722\,
            I => \N__42719\
        );

    \I__7908\ : Span4Mux_h
    port map (
            O => \N__42719\,
            I => \N__42716\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__42716\,
            I => \N__42713\
        );

    \I__7906\ : Odrv4
    port map (
            O => \N__42713\,
            I => \ALU.d_RNI0PI3E1Z0Z_8\
        );

    \I__7905\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42707\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__42707\,
            I => \ALU.mult_9_10\
        );

    \I__7903\ : InMux
    port map (
            O => \N__42704\,
            I => \ALU.mult_9_c9\
        );

    \I__7902\ : InMux
    port map (
            O => \N__42701\,
            I => \N__42698\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__42698\,
            I => \ALU.d_RNIFCNKLZ0Z_9\
        );

    \I__7900\ : CascadeMux
    port map (
            O => \N__42695\,
            I => \N__42692\
        );

    \I__7899\ : InMux
    port map (
            O => \N__42692\,
            I => \N__42689\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__42689\,
            I => \N__42686\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__42686\,
            I => \ALU.d_RNIDR5C61Z0Z_8\
        );

    \I__7896\ : InMux
    port map (
            O => \N__42683\,
            I => \N__42680\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__42680\,
            I => \ALU.mult_9_11\
        );

    \I__7894\ : InMux
    port map (
            O => \N__42677\,
            I => \ALU.mult_9_c10\
        );

    \I__7893\ : CascadeMux
    port map (
            O => \N__42674\,
            I => \N__42671\
        );

    \I__7892\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42668\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__42668\,
            I => \ALU.d_RNIG61LGZ0Z_9\
        );

    \I__7890\ : InMux
    port map (
            O => \N__42665\,
            I => \N__42662\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__42662\,
            I => \ALU.mult_9_12\
        );

    \I__7888\ : InMux
    port map (
            O => \N__42659\,
            I => \ALU.mult_9_c11\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__42656\,
            I => \N__42653\
        );

    \I__7886\ : InMux
    port map (
            O => \N__42653\,
            I => \N__42650\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__42650\,
            I => \N__42647\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__42647\,
            I => \N__42644\
        );

    \I__7883\ : Odrv4
    port map (
            O => \N__42644\,
            I => \ALU.d_RNI68LSHZ0Z_9\
        );

    \I__7882\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42638\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__42638\,
            I => \ALU.mult_9_13\
        );

    \I__7880\ : InMux
    port map (
            O => \N__42635\,
            I => \ALU.mult_9_c12\
        );

    \I__7879\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42629\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__42629\,
            I => \N__42626\
        );

    \I__7877\ : Span4Mux_v
    port map (
            O => \N__42626\,
            I => \N__42623\
        );

    \I__7876\ : Sp12to4
    port map (
            O => \N__42623\,
            I => \N__42620\
        );

    \I__7875\ : Odrv12
    port map (
            O => \N__42620\,
            I => \ALU.d_RNISSV4IZ0Z_9\
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__42617\,
            I => \N__42614\
        );

    \I__7873\ : InMux
    port map (
            O => \N__42614\,
            I => \N__42611\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__42611\,
            I => \N__42608\
        );

    \I__7871\ : Span12Mux_h
    port map (
            O => \N__42608\,
            I => \N__42605\
        );

    \I__7870\ : Odrv12
    port map (
            O => \N__42605\,
            I => \ALU.d_RNI371041Z0Z_8\
        );

    \I__7869\ : InMux
    port map (
            O => \N__42602\,
            I => \N__42599\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__42599\,
            I => \ALU.mult_9_14\
        );

    \I__7867\ : InMux
    port map (
            O => \N__42596\,
            I => \ALU.mult_9_c13\
        );

    \I__7866\ : InMux
    port map (
            O => \N__42593\,
            I => \N__42590\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__42590\,
            I => \N__42587\
        );

    \I__7864\ : Span4Mux_h
    port map (
            O => \N__42587\,
            I => \N__42584\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__42584\,
            I => \N__42581\
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__42581\,
            I => \ALU.c_RNI0QV651Z0Z_10\
        );

    \I__7861\ : InMux
    port map (
            O => \N__42578\,
            I => \ALU.mult_9_c14\
        );

    \I__7860\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42572\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__42572\,
            I => \ALU.N_862\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__42569\,
            I => \ALU.N_862_cascade_\
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__42566\,
            I => \ALU.N_922_cascade_\
        );

    \I__7856\ : InMux
    port map (
            O => \N__42563\,
            I => \N__42560\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__42560\,
            I => \N__42557\
        );

    \I__7854\ : Span4Mux_h
    port map (
            O => \N__42557\,
            I => \N__42554\
        );

    \I__7853\ : Odrv4
    port map (
            O => \N__42554\,
            I => \ALU.d_RNIR6J013Z0Z_2\
        );

    \I__7852\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42543\
        );

    \I__7851\ : InMux
    port map (
            O => \N__42550\,
            I => \N__42540\
        );

    \I__7850\ : InMux
    port map (
            O => \N__42549\,
            I => \N__42537\
        );

    \I__7849\ : InMux
    port map (
            O => \N__42548\,
            I => \N__42533\
        );

    \I__7848\ : InMux
    port map (
            O => \N__42547\,
            I => \N__42530\
        );

    \I__7847\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42526\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__42543\,
            I => \N__42523\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__42540\,
            I => \N__42520\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__42537\,
            I => \N__42517\
        );

    \I__7843\ : InMux
    port map (
            O => \N__42536\,
            I => \N__42514\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__42533\,
            I => \N__42509\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__42530\,
            I => \N__42509\
        );

    \I__7840\ : InMux
    port map (
            O => \N__42529\,
            I => \N__42506\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__42526\,
            I => \N__42501\
        );

    \I__7838\ : Span4Mux_h
    port map (
            O => \N__42523\,
            I => \N__42501\
        );

    \I__7837\ : Span4Mux_v
    port map (
            O => \N__42520\,
            I => \N__42498\
        );

    \I__7836\ : Span4Mux_v
    port map (
            O => \N__42517\,
            I => \N__42495\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__42514\,
            I => \N__42490\
        );

    \I__7834\ : Span4Mux_v
    port map (
            O => \N__42509\,
            I => \N__42490\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__42506\,
            I => \N__42485\
        );

    \I__7832\ : Span4Mux_h
    port map (
            O => \N__42501\,
            I => \N__42485\
        );

    \I__7831\ : Span4Mux_h
    port map (
            O => \N__42498\,
            I => \N__42482\
        );

    \I__7830\ : Span4Mux_h
    port map (
            O => \N__42495\,
            I => \N__42477\
        );

    \I__7829\ : Span4Mux_v
    port map (
            O => \N__42490\,
            I => \N__42477\
        );

    \I__7828\ : Span4Mux_v
    port map (
            O => \N__42485\,
            I => \N__42474\
        );

    \I__7827\ : Span4Mux_h
    port map (
            O => \N__42482\,
            I => \N__42471\
        );

    \I__7826\ : Odrv4
    port map (
            O => \N__42477\,
            I => \ALU.d_RNI1AHUF8Z0Z_2\
        );

    \I__7825\ : Odrv4
    port map (
            O => \N__42474\,
            I => \ALU.d_RNI1AHUF8Z0Z_2\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__42471\,
            I => \ALU.d_RNI1AHUF8Z0Z_2\
        );

    \I__7823\ : InMux
    port map (
            O => \N__42464\,
            I => \N__42460\
        );

    \I__7822\ : CascadeMux
    port map (
            O => \N__42463\,
            I => \N__42457\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__42460\,
            I => \N__42454\
        );

    \I__7820\ : InMux
    port map (
            O => \N__42457\,
            I => \N__42451\
        );

    \I__7819\ : Odrv12
    port map (
            O => \N__42454\,
            I => \ALU.mult_25_10\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__42451\,
            I => \ALU.mult_25_10\
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__42446\,
            I => \N__42443\
        );

    \I__7816\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42440\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__42440\,
            I => \ALU.mult_11_10\
        );

    \I__7814\ : InMux
    port map (
            O => \N__42437\,
            I => \N__42434\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__42434\,
            I => \N__42431\
        );

    \I__7812\ : Span4Mux_h
    port map (
            O => \N__42431\,
            I => \N__42428\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__42428\,
            I => \ALU.mult_293_c_RNIOCJMDZ0Z9\
        );

    \I__7810\ : CascadeMux
    port map (
            O => \N__42425\,
            I => \N__42422\
        );

    \I__7809\ : InMux
    port map (
            O => \N__42422\,
            I => \N__42419\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__42419\,
            I => \ALU.mult_11_11\
        );

    \I__7807\ : InMux
    port map (
            O => \N__42416\,
            I => \N__42413\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__42413\,
            I => \N__42410\
        );

    \I__7805\ : Span4Mux_h
    port map (
            O => \N__42410\,
            I => \N__42407\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__42407\,
            I => \ALU.mult_21_11\
        );

    \I__7803\ : InMux
    port map (
            O => \N__42404\,
            I => \ALU.mult_21_c10\
        );

    \I__7802\ : InMux
    port map (
            O => \N__42401\,
            I => \N__42397\
        );

    \I__7801\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42394\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__42397\,
            I => \ALU.mult_21_12\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__42394\,
            I => \ALU.mult_21_12\
        );

    \I__7798\ : InMux
    port map (
            O => \N__42389\,
            I => \ALU.mult_21_c11\
        );

    \I__7797\ : InMux
    port map (
            O => \N__42386\,
            I => \N__42383\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__42383\,
            I => \ALU.mult_21_13\
        );

    \I__7795\ : InMux
    port map (
            O => \N__42380\,
            I => \ALU.mult_21_c12\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__42377\,
            I => \N__42374\
        );

    \I__7793\ : InMux
    port map (
            O => \N__42374\,
            I => \N__42371\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__42371\,
            I => \N__42367\
        );

    \I__7791\ : InMux
    port map (
            O => \N__42370\,
            I => \N__42364\
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__42367\,
            I => \ALU.mult_21_14\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__42364\,
            I => \ALU.mult_21_14\
        );

    \I__7788\ : InMux
    port map (
            O => \N__42359\,
            I => \ALU.mult_21_c13\
        );

    \I__7787\ : InMux
    port map (
            O => \N__42356\,
            I => \N__42353\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__42353\,
            I => \ALU.mult_23_15\
        );

    \I__7785\ : InMux
    port map (
            O => \N__42350\,
            I => \ALU.mult_21_c14\
        );

    \I__7784\ : InMux
    port map (
            O => \N__42347\,
            I => \N__42344\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__42344\,
            I => \N__42341\
        );

    \I__7782\ : Span4Mux_v
    port map (
            O => \N__42341\,
            I => \N__42338\
        );

    \I__7781\ : Odrv4
    port map (
            O => \N__42338\,
            I => \ALU.mult_476_c_RNIFLP0OZ0Z7\
        );

    \I__7780\ : InMux
    port map (
            O => \N__42335\,
            I => \N__42329\
        );

    \I__7779\ : InMux
    port map (
            O => \N__42334\,
            I => \N__42329\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__42329\,
            I => \N__42326\
        );

    \I__7777\ : Span4Mux_h
    port map (
            O => \N__42326\,
            I => \N__42323\
        );

    \I__7776\ : Span4Mux_h
    port map (
            O => \N__42323\,
            I => \N__42319\
        );

    \I__7775\ : CascadeMux
    port map (
            O => \N__42322\,
            I => \N__42316\
        );

    \I__7774\ : Span4Mux_h
    port map (
            O => \N__42319\,
            I => \N__42313\
        );

    \I__7773\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42310\
        );

    \I__7772\ : Odrv4
    port map (
            O => \N__42313\,
            I => \CONTROL.addrstack_1_7\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__42310\,
            I => \CONTROL.addrstack_1_7\
        );

    \I__7770\ : InMux
    port map (
            O => \N__42305\,
            I => \N__42299\
        );

    \I__7769\ : InMux
    port map (
            O => \N__42304\,
            I => \N__42299\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__42299\,
            I => \CONTROL.g0_4Z0Z_2\
        );

    \I__7767\ : CascadeMux
    port map (
            O => \N__42296\,
            I => \CONTROL.g0_i_m2_1_cascade_\
        );

    \I__7766\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42290\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__42290\,
            I => \CONTROL.g1_1\
        );

    \I__7764\ : InMux
    port map (
            O => \N__42287\,
            I => \N__42284\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__42284\,
            I => \N__42281\
        );

    \I__7762\ : Span4Mux_v
    port map (
            O => \N__42281\,
            I => \N__42277\
        );

    \I__7761\ : InMux
    port map (
            O => \N__42280\,
            I => \N__42274\
        );

    \I__7760\ : Sp12to4
    port map (
            O => \N__42277\,
            I => \N__42271\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__42274\,
            I => \CONTROL.addrstackptrZ0Z_7\
        );

    \I__7758\ : Odrv12
    port map (
            O => \N__42271\,
            I => \CONTROL.addrstackptrZ0Z_7\
        );

    \I__7757\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42258\
        );

    \I__7756\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42255\
        );

    \I__7755\ : InMux
    port map (
            O => \N__42264\,
            I => \N__42250\
        );

    \I__7754\ : InMux
    port map (
            O => \N__42263\,
            I => \N__42250\
        );

    \I__7753\ : CascadeMux
    port map (
            O => \N__42262\,
            I => \N__42245\
        );

    \I__7752\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42241\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__42258\,
            I => \N__42236\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__42255\,
            I => \N__42236\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__42250\,
            I => \N__42232\
        );

    \I__7748\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42225\
        );

    \I__7747\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42225\
        );

    \I__7746\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42225\
        );

    \I__7745\ : InMux
    port map (
            O => \N__42244\,
            I => \N__42222\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__42241\,
            I => \N__42217\
        );

    \I__7743\ : Span4Mux_h
    port map (
            O => \N__42236\,
            I => \N__42213\
        );

    \I__7742\ : CascadeMux
    port map (
            O => \N__42235\,
            I => \N__42209\
        );

    \I__7741\ : Span4Mux_h
    port map (
            O => \N__42232\,
            I => \N__42203\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__42225\,
            I => \N__42203\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__42222\,
            I => \N__42200\
        );

    \I__7738\ : InMux
    port map (
            O => \N__42221\,
            I => \N__42197\
        );

    \I__7737\ : CascadeMux
    port map (
            O => \N__42220\,
            I => \N__42192\
        );

    \I__7736\ : Span4Mux_h
    port map (
            O => \N__42217\,
            I => \N__42189\
        );

    \I__7735\ : InMux
    port map (
            O => \N__42216\,
            I => \N__42186\
        );

    \I__7734\ : Span4Mux_h
    port map (
            O => \N__42213\,
            I => \N__42183\
        );

    \I__7733\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42176\
        );

    \I__7732\ : InMux
    port map (
            O => \N__42209\,
            I => \N__42176\
        );

    \I__7731\ : InMux
    port map (
            O => \N__42208\,
            I => \N__42176\
        );

    \I__7730\ : Span4Mux_h
    port map (
            O => \N__42203\,
            I => \N__42169\
        );

    \I__7729\ : Span4Mux_h
    port map (
            O => \N__42200\,
            I => \N__42169\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__42197\,
            I => \N__42169\
        );

    \I__7727\ : InMux
    port map (
            O => \N__42196\,
            I => \N__42162\
        );

    \I__7726\ : InMux
    port map (
            O => \N__42195\,
            I => \N__42162\
        );

    \I__7725\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42162\
        );

    \I__7724\ : Odrv4
    port map (
            O => \N__42189\,
            I => \PROM_ROMDATA_dintern_5ro\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__42186\,
            I => \PROM_ROMDATA_dintern_5ro\
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__42183\,
            I => \PROM_ROMDATA_dintern_5ro\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__42176\,
            I => \PROM_ROMDATA_dintern_5ro\
        );

    \I__7720\ : Odrv4
    port map (
            O => \N__42169\,
            I => \PROM_ROMDATA_dintern_5ro\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__42162\,
            I => \PROM_ROMDATA_dintern_5ro\
        );

    \I__7718\ : InMux
    port map (
            O => \N__42149\,
            I => \N__42146\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__42146\,
            I => \N__42143\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__42143\,
            I => \N__42140\
        );

    \I__7715\ : Odrv4
    port map (
            O => \N__42140\,
            I => \CONTROL.g0_2_iZ0Z_1\
        );

    \I__7714\ : InMux
    port map (
            O => \N__42137\,
            I => \N__42134\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__42134\,
            I => \PROM.ROMDATA.m381_am\
        );

    \I__7712\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42128\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__42128\,
            I => \N__42125\
        );

    \I__7710\ : Span4Mux_h
    port map (
            O => \N__42125\,
            I => \N__42122\
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__42122\,
            I => \PROM.ROMDATA.m375_am\
        );

    \I__7708\ : InMux
    port map (
            O => \N__42119\,
            I => \N__42116\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__42116\,
            I => \PROM.ROMDATA.m382_ns_1\
        );

    \I__7706\ : CascadeMux
    port map (
            O => \N__42113\,
            I => \N__42110\
        );

    \I__7705\ : InMux
    port map (
            O => \N__42110\,
            I => \N__42107\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__42107\,
            I => \N__42104\
        );

    \I__7703\ : Span4Mux_h
    port map (
            O => \N__42104\,
            I => \N__42101\
        );

    \I__7702\ : Span4Mux_h
    port map (
            O => \N__42101\,
            I => \N__42098\
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__42098\,
            I => \ALU.rshift_3_ns_1_0\
        );

    \I__7700\ : CascadeMux
    port map (
            O => \N__42095\,
            I => \ALU.N_858_cascade_\
        );

    \I__7699\ : CascadeMux
    port map (
            O => \N__42092\,
            I => \ALU.rshift_15_ns_1_0_cascade_\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__42089\,
            I => \ALU.rshift_3_ns_1_4_cascade_\
        );

    \I__7697\ : InMux
    port map (
            O => \N__42086\,
            I => \N__42083\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__42083\,
            I => \N__42077\
        );

    \I__7695\ : InMux
    port map (
            O => \N__42082\,
            I => \N__42074\
        );

    \I__7694\ : InMux
    port map (
            O => \N__42081\,
            I => \N__42071\
        );

    \I__7693\ : InMux
    port map (
            O => \N__42080\,
            I => \N__42067\
        );

    \I__7692\ : Span4Mux_v
    port map (
            O => \N__42077\,
            I => \N__42060\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__42074\,
            I => \N__42060\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__42071\,
            I => \N__42060\
        );

    \I__7689\ : InMux
    port map (
            O => \N__42070\,
            I => \N__42057\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__42067\,
            I => \N__42054\
        );

    \I__7687\ : Span4Mux_h
    port map (
            O => \N__42060\,
            I => \N__42049\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__42057\,
            I => \N__42049\
        );

    \I__7685\ : Odrv12
    port map (
            O => \N__42054\,
            I => \CONTROL.un1_programCounter9_reto_rep1\
        );

    \I__7684\ : Odrv4
    port map (
            O => \N__42049\,
            I => \CONTROL.un1_programCounter9_reto_rep1\
        );

    \I__7683\ : InMux
    port map (
            O => \N__42044\,
            I => \N__42041\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__42041\,
            I => \N__42038\
        );

    \I__7681\ : Span4Mux_v
    port map (
            O => \N__42038\,
            I => \N__42035\
        );

    \I__7680\ : Span4Mux_h
    port map (
            O => \N__42035\,
            I => \N__42032\
        );

    \I__7679\ : Span4Mux_h
    port map (
            O => \N__42032\,
            I => \N__42029\
        );

    \I__7678\ : Odrv4
    port map (
            O => \N__42029\,
            I => \CONTROL.g0_2Z0Z_1\
        );

    \I__7677\ : InMux
    port map (
            O => \N__42026\,
            I => \N__42023\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__42023\,
            I => \N__42020\
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__42020\,
            I => \CONTROL.N_133_0_0\
        );

    \I__7674\ : InMux
    port map (
            O => \N__42017\,
            I => \N__42014\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__42014\,
            I => \CONTROL.N_114_i\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__42011\,
            I => \N__42008\
        );

    \I__7671\ : InMux
    port map (
            O => \N__42008\,
            I => \N__42005\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__42005\,
            I => \N__42002\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__42002\,
            I => \N__41999\
        );

    \I__7668\ : Span4Mux_h
    port map (
            O => \N__41999\,
            I => \N__41996\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__41996\,
            I => \N__41993\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__41993\,
            I => \CONTROL.g1_1_4\
        );

    \I__7665\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41987\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__41987\,
            I => \N__41983\
        );

    \I__7663\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41978\
        );

    \I__7662\ : Span4Mux_v
    port map (
            O => \N__41983\,
            I => \N__41973\
        );

    \I__7661\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41970\
        );

    \I__7660\ : InMux
    port map (
            O => \N__41981\,
            I => \N__41967\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__41978\,
            I => \N__41964\
        );

    \I__7658\ : InMux
    port map (
            O => \N__41977\,
            I => \N__41961\
        );

    \I__7657\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41955\
        );

    \I__7656\ : Span4Mux_v
    port map (
            O => \N__41973\,
            I => \N__41952\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__41970\,
            I => \N__41949\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__41967\,
            I => \N__41946\
        );

    \I__7653\ : Span4Mux_h
    port map (
            O => \N__41964\,
            I => \N__41941\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__41961\,
            I => \N__41941\
        );

    \I__7651\ : InMux
    port map (
            O => \N__41960\,
            I => \N__41938\
        );

    \I__7650\ : InMux
    port map (
            O => \N__41959\,
            I => \N__41933\
        );

    \I__7649\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41933\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__41955\,
            I => \N__41930\
        );

    \I__7647\ : Span4Mux_v
    port map (
            O => \N__41952\,
            I => \N__41927\
        );

    \I__7646\ : Span4Mux_h
    port map (
            O => \N__41949\,
            I => \N__41924\
        );

    \I__7645\ : Sp12to4
    port map (
            O => \N__41946\,
            I => \N__41916\
        );

    \I__7644\ : Sp12to4
    port map (
            O => \N__41941\,
            I => \N__41916\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__41938\,
            I => \N__41916\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__41933\,
            I => \N__41913\
        );

    \I__7641\ : Span4Mux_v
    port map (
            O => \N__41930\,
            I => \N__41910\
        );

    \I__7640\ : Span4Mux_h
    port map (
            O => \N__41927\,
            I => \N__41905\
        );

    \I__7639\ : Span4Mux_h
    port map (
            O => \N__41924\,
            I => \N__41905\
        );

    \I__7638\ : InMux
    port map (
            O => \N__41923\,
            I => \N__41902\
        );

    \I__7637\ : Span12Mux_v
    port map (
            O => \N__41916\,
            I => \N__41899\
        );

    \I__7636\ : Odrv4
    port map (
            O => \N__41913\,
            I => \CONTROL.un1_busState114_2_0_0\
        );

    \I__7635\ : Odrv4
    port map (
            O => \N__41910\,
            I => \CONTROL.un1_busState114_2_0_0\
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__41905\,
            I => \CONTROL.un1_busState114_2_0_0\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__41902\,
            I => \CONTROL.un1_busState114_2_0_0\
        );

    \I__7632\ : Odrv12
    port map (
            O => \N__41899\,
            I => \CONTROL.un1_busState114_2_0_0\
        );

    \I__7631\ : CascadeMux
    port map (
            O => \N__41888\,
            I => \CONTROL.g1_1_cascade_\
        );

    \I__7630\ : CascadeMux
    port map (
            O => \N__41885\,
            I => \N__41882\
        );

    \I__7629\ : InMux
    port map (
            O => \N__41882\,
            I => \N__41879\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__41879\,
            I => \N__41876\
        );

    \I__7627\ : Span4Mux_v
    port map (
            O => \N__41876\,
            I => \N__41873\
        );

    \I__7626\ : Span4Mux_h
    port map (
            O => \N__41873\,
            I => \N__41870\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__41870\,
            I => \N__41867\
        );

    \I__7624\ : Odrv4
    port map (
            O => \N__41867\,
            I => \CONTROL.addrstackptr_N_7_i\
        );

    \I__7623\ : CascadeMux
    port map (
            O => \N__41864\,
            I => \N__41861\
        );

    \I__7622\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41858\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__41858\,
            I => \N__41855\
        );

    \I__7620\ : Odrv4
    port map (
            O => \N__41855\,
            I => \CONTROL.g1_0_0\
        );

    \I__7619\ : InMux
    port map (
            O => \N__41852\,
            I => \N__41849\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__41849\,
            I => \CONTROL.g0_i_m2_1\
        );

    \I__7617\ : InMux
    port map (
            O => \N__41846\,
            I => \N__41843\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__41843\,
            I => \N__41840\
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__41840\,
            I => \PROM.ROMDATA.m31\
        );

    \I__7614\ : CascadeMux
    port map (
            O => \N__41837\,
            I => \m125_e_cascade_\
        );

    \I__7613\ : InMux
    port map (
            O => \N__41834\,
            I => \N__41830\
        );

    \I__7612\ : InMux
    port map (
            O => \N__41833\,
            I => \N__41827\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__41830\,
            I => \N__41824\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__41827\,
            I => \PROM.ROMDATA.N_557_mux\
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__41824\,
            I => \PROM.ROMDATA.N_557_mux\
        );

    \I__7608\ : InMux
    port map (
            O => \N__41819\,
            I => \N__41816\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__41816\,
            I => \N__41813\
        );

    \I__7606\ : Odrv4
    port map (
            O => \N__41813\,
            I => \PROM.ROMDATA.m77\
        );

    \I__7605\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41807\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__41807\,
            I => \N__41802\
        );

    \I__7603\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41797\
        );

    \I__7602\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41797\
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__41802\,
            I => m93_ns
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__41797\,
            I => m93_ns
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__41792\,
            I => \m93_ns_cascade_\
        );

    \I__7598\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41786\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__41786\,
            I => \N__41783\
        );

    \I__7596\ : Span4Mux_v
    port map (
            O => \N__41783\,
            I => \N__41780\
        );

    \I__7595\ : Span4Mux_h
    port map (
            O => \N__41780\,
            I => \N__41777\
        );

    \I__7594\ : Span4Mux_h
    port map (
            O => \N__41777\,
            I => \N__41774\
        );

    \I__7593\ : Odrv4
    port map (
            O => \N__41774\,
            I => \CONTROL.addrstack_5\
        );

    \I__7592\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41768\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__41768\,
            I => \N__41765\
        );

    \I__7590\ : Span4Mux_h
    port map (
            O => \N__41765\,
            I => \N__41760\
        );

    \I__7589\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41757\
        );

    \I__7588\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41754\
        );

    \I__7587\ : Odrv4
    port map (
            O => \N__41760\,
            I => \CONTROL.addrstack_reto_5\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__41757\,
            I => \CONTROL.addrstack_reto_5\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__41754\,
            I => \CONTROL.addrstack_reto_5\
        );

    \I__7584\ : InMux
    port map (
            O => \N__41747\,
            I => \N__41744\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__41744\,
            I => \N__41741\
        );

    \I__7582\ : Span4Mux_v
    port map (
            O => \N__41741\,
            I => \N__41737\
        );

    \I__7581\ : InMux
    port map (
            O => \N__41740\,
            I => \N__41734\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__41737\,
            I => \N__41729\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__41734\,
            I => \N__41729\
        );

    \I__7578\ : Span4Mux_h
    port map (
            O => \N__41729\,
            I => \N__41726\
        );

    \I__7577\ : Odrv4
    port map (
            O => \N__41726\,
            I => \CONTROL.programCounter_1_5\
        );

    \I__7576\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41720\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__41720\,
            I => \N__41717\
        );

    \I__7574\ : Span4Mux_h
    port map (
            O => \N__41717\,
            I => \N__41713\
        );

    \I__7573\ : InMux
    port map (
            O => \N__41716\,
            I => \N__41710\
        );

    \I__7572\ : Odrv4
    port map (
            O => \N__41713\,
            I => \CONTROL.programCounter_1_reto_5\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__41710\,
            I => \CONTROL.programCounter_1_reto_5\
        );

    \I__7570\ : CascadeMux
    port map (
            O => \N__41705\,
            I => \CONTROL.N_86_0_cascade_\
        );

    \I__7569\ : CascadeMux
    port map (
            O => \N__41702\,
            I => \N__41699\
        );

    \I__7568\ : InMux
    port map (
            O => \N__41699\,
            I => \N__41693\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__41698\,
            I => \N__41690\
        );

    \I__7566\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41685\
        );

    \I__7565\ : CascadeMux
    port map (
            O => \N__41696\,
            I => \N__41682\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__41693\,
            I => \N__41679\
        );

    \I__7563\ : InMux
    port map (
            O => \N__41690\,
            I => \N__41676\
        );

    \I__7562\ : InMux
    port map (
            O => \N__41689\,
            I => \N__41671\
        );

    \I__7561\ : InMux
    port map (
            O => \N__41688\,
            I => \N__41671\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__41685\,
            I => \N__41667\
        );

    \I__7559\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41664\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__41679\,
            I => \N__41659\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__41676\,
            I => \N__41659\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__41671\,
            I => \N__41656\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__41670\,
            I => \N__41652\
        );

    \I__7554\ : Span4Mux_v
    port map (
            O => \N__41667\,
            I => \N__41647\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41642\
        );

    \I__7552\ : Span4Mux_h
    port map (
            O => \N__41659\,
            I => \N__41642\
        );

    \I__7551\ : Span4Mux_h
    port map (
            O => \N__41656\,
            I => \N__41639\
        );

    \I__7550\ : InMux
    port map (
            O => \N__41655\,
            I => \N__41636\
        );

    \I__7549\ : InMux
    port map (
            O => \N__41652\,
            I => \N__41633\
        );

    \I__7548\ : InMux
    port map (
            O => \N__41651\,
            I => \N__41628\
        );

    \I__7547\ : InMux
    port map (
            O => \N__41650\,
            I => \N__41628\
        );

    \I__7546\ : Odrv4
    port map (
            O => \N__41647\,
            I => \controlWord_1\
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__41642\,
            I => \controlWord_1\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__41639\,
            I => \controlWord_1\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__41636\,
            I => \controlWord_1\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__41633\,
            I => \controlWord_1\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__41628\,
            I => \controlWord_1\
        );

    \I__7540\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41612\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__41612\,
            I => \N__41609\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__41609\,
            I => \N__41606\
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__41606\,
            I => \CONTROL.N_135\
        );

    \I__7536\ : InMux
    port map (
            O => \N__41603\,
            I => \N__41597\
        );

    \I__7535\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41597\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__41597\,
            I => \N__41591\
        );

    \I__7533\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41586\
        );

    \I__7532\ : InMux
    port map (
            O => \N__41595\,
            I => \N__41586\
        );

    \I__7531\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41583\
        );

    \I__7530\ : Span4Mux_v
    port map (
            O => \N__41591\,
            I => \N__41577\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__41586\,
            I => \N__41572\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__41583\,
            I => \N__41569\
        );

    \I__7527\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41566\
        );

    \I__7526\ : InMux
    port map (
            O => \N__41581\,
            I => \N__41563\
        );

    \I__7525\ : InMux
    port map (
            O => \N__41580\,
            I => \N__41560\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__41577\,
            I => \N__41555\
        );

    \I__7523\ : InMux
    port map (
            O => \N__41576\,
            I => \N__41550\
        );

    \I__7522\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41550\
        );

    \I__7521\ : Span4Mux_h
    port map (
            O => \N__41572\,
            I => \N__41545\
        );

    \I__7520\ : Span4Mux_h
    port map (
            O => \N__41569\,
            I => \N__41545\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__41566\,
            I => \N__41542\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__41563\,
            I => \N__41539\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__41560\,
            I => \N__41536\
        );

    \I__7516\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41531\
        );

    \I__7515\ : InMux
    port map (
            O => \N__41558\,
            I => \N__41531\
        );

    \I__7514\ : Span4Mux_h
    port map (
            O => \N__41555\,
            I => \N__41526\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__41550\,
            I => \N__41526\
        );

    \I__7512\ : Span4Mux_h
    port map (
            O => \N__41545\,
            I => \N__41523\
        );

    \I__7511\ : Span4Mux_h
    port map (
            O => \N__41542\,
            I => \N__41518\
        );

    \I__7510\ : Span4Mux_h
    port map (
            O => \N__41539\,
            I => \N__41518\
        );

    \I__7509\ : Span12Mux_h
    port map (
            O => \N__41536\,
            I => \N__41515\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__41531\,
            I => \CONTROL.N_74_0\
        );

    \I__7507\ : Odrv4
    port map (
            O => \N__41526\,
            I => \CONTROL.N_74_0\
        );

    \I__7506\ : Odrv4
    port map (
            O => \N__41523\,
            I => \CONTROL.N_74_0\
        );

    \I__7505\ : Odrv4
    port map (
            O => \N__41518\,
            I => \CONTROL.N_74_0\
        );

    \I__7504\ : Odrv12
    port map (
            O => \N__41515\,
            I => \CONTROL.N_74_0\
        );

    \I__7503\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41500\
        );

    \I__7502\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41497\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__41500\,
            I => \N__41493\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__41497\,
            I => \N__41490\
        );

    \I__7499\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41485\
        );

    \I__7498\ : Span4Mux_v
    port map (
            O => \N__41493\,
            I => \N__41480\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__41490\,
            I => \N__41480\
        );

    \I__7496\ : InMux
    port map (
            O => \N__41489\,
            I => \N__41477\
        );

    \I__7495\ : InMux
    port map (
            O => \N__41488\,
            I => \N__41473\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__41485\,
            I => \N__41470\
        );

    \I__7493\ : Span4Mux_h
    port map (
            O => \N__41480\,
            I => \N__41465\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__41477\,
            I => \N__41465\
        );

    \I__7491\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41460\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__41473\,
            I => \N__41457\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__41470\,
            I => \N__41452\
        );

    \I__7488\ : Span4Mux_h
    port map (
            O => \N__41465\,
            I => \N__41452\
        );

    \I__7487\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41449\
        );

    \I__7486\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41446\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__41460\,
            I => \CONTROL.N_249\
        );

    \I__7484\ : Odrv12
    port map (
            O => \N__41457\,
            I => \CONTROL.N_249\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__41452\,
            I => \CONTROL.N_249\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__41449\,
            I => \CONTROL.N_249\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__41446\,
            I => \CONTROL.N_249\
        );

    \I__7480\ : CascadeMux
    port map (
            O => \N__41435\,
            I => \N__41425\
        );

    \I__7479\ : InMux
    port map (
            O => \N__41434\,
            I => \N__41420\
        );

    \I__7478\ : CascadeMux
    port map (
            O => \N__41433\,
            I => \N__41417\
        );

    \I__7477\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41412\
        );

    \I__7476\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41409\
        );

    \I__7475\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41405\
        );

    \I__7474\ : InMux
    port map (
            O => \N__41429\,
            I => \N__41398\
        );

    \I__7473\ : InMux
    port map (
            O => \N__41428\,
            I => \N__41398\
        );

    \I__7472\ : InMux
    port map (
            O => \N__41425\,
            I => \N__41398\
        );

    \I__7471\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41388\
        );

    \I__7470\ : InMux
    port map (
            O => \N__41423\,
            I => \N__41385\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__41420\,
            I => \N__41382\
        );

    \I__7468\ : InMux
    port map (
            O => \N__41417\,
            I => \N__41379\
        );

    \I__7467\ : CascadeMux
    port map (
            O => \N__41416\,
            I => \N__41376\
        );

    \I__7466\ : CascadeMux
    port map (
            O => \N__41415\,
            I => \N__41373\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__41412\,
            I => \N__41366\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__41409\,
            I => \N__41366\
        );

    \I__7463\ : InMux
    port map (
            O => \N__41408\,
            I => \N__41363\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__41405\,
            I => \N__41358\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__41398\,
            I => \N__41358\
        );

    \I__7460\ : CascadeMux
    port map (
            O => \N__41397\,
            I => \N__41353\
        );

    \I__7459\ : InMux
    port map (
            O => \N__41396\,
            I => \N__41350\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__41395\,
            I => \N__41347\
        );

    \I__7457\ : InMux
    port map (
            O => \N__41394\,
            I => \N__41340\
        );

    \I__7456\ : InMux
    port map (
            O => \N__41393\,
            I => \N__41340\
        );

    \I__7455\ : InMux
    port map (
            O => \N__41392\,
            I => \N__41340\
        );

    \I__7454\ : InMux
    port map (
            O => \N__41391\,
            I => \N__41337\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__41388\,
            I => \N__41328\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__41385\,
            I => \N__41328\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__41382\,
            I => \N__41328\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__41379\,
            I => \N__41328\
        );

    \I__7449\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41319\
        );

    \I__7448\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41319\
        );

    \I__7447\ : InMux
    port map (
            O => \N__41372\,
            I => \N__41319\
        );

    \I__7446\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41319\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__41366\,
            I => \N__41312\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__41363\,
            I => \N__41312\
        );

    \I__7443\ : Span4Mux_v
    port map (
            O => \N__41358\,
            I => \N__41312\
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__41357\,
            I => \N__41309\
        );

    \I__7441\ : CascadeMux
    port map (
            O => \N__41356\,
            I => \N__41306\
        );

    \I__7440\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41302\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__41350\,
            I => \N__41299\
        );

    \I__7438\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41296\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__41340\,
            I => \N__41289\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__41337\,
            I => \N__41289\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__41328\,
            I => \N__41289\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__41319\,
            I => \N__41284\
        );

    \I__7433\ : Span4Mux_h
    port map (
            O => \N__41312\,
            I => \N__41284\
        );

    \I__7432\ : InMux
    port map (
            O => \N__41309\,
            I => \N__41277\
        );

    \I__7431\ : InMux
    port map (
            O => \N__41306\,
            I => \N__41277\
        );

    \I__7430\ : InMux
    port map (
            O => \N__41305\,
            I => \N__41277\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__41302\,
            I => \controlWord_5\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__41299\,
            I => \controlWord_5\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__41296\,
            I => \controlWord_5\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__41289\,
            I => \controlWord_5\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__41284\,
            I => \controlWord_5\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__41277\,
            I => \controlWord_5\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__41264\,
            I => \CONTROL.N_74_0_cascade_\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__41261\,
            I => \N__41253\
        );

    \I__7421\ : InMux
    port map (
            O => \N__41260\,
            I => \N__41250\
        );

    \I__7420\ : CascadeMux
    port map (
            O => \N__41259\,
            I => \N__41242\
        );

    \I__7419\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41236\
        );

    \I__7418\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41236\
        );

    \I__7417\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41230\
        );

    \I__7416\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41227\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__41250\,
            I => \N__41224\
        );

    \I__7414\ : InMux
    port map (
            O => \N__41249\,
            I => \N__41211\
        );

    \I__7413\ : InMux
    port map (
            O => \N__41248\,
            I => \N__41211\
        );

    \I__7412\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41211\
        );

    \I__7411\ : InMux
    port map (
            O => \N__41246\,
            I => \N__41211\
        );

    \I__7410\ : InMux
    port map (
            O => \N__41245\,
            I => \N__41211\
        );

    \I__7409\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41211\
        );

    \I__7408\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41207\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__41236\,
            I => \N__41204\
        );

    \I__7406\ : CascadeMux
    port map (
            O => \N__41235\,
            I => \N__41198\
        );

    \I__7405\ : InMux
    port map (
            O => \N__41234\,
            I => \N__41195\
        );

    \I__7404\ : InMux
    port map (
            O => \N__41233\,
            I => \N__41188\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__41230\,
            I => \N__41185\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__41227\,
            I => \N__41182\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__41224\,
            I => \N__41177\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__41211\,
            I => \N__41177\
        );

    \I__7399\ : InMux
    port map (
            O => \N__41210\,
            I => \N__41174\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__41207\,
            I => \N__41171\
        );

    \I__7397\ : Span4Mux_h
    port map (
            O => \N__41204\,
            I => \N__41168\
        );

    \I__7396\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41163\
        );

    \I__7395\ : InMux
    port map (
            O => \N__41202\,
            I => \N__41163\
        );

    \I__7394\ : InMux
    port map (
            O => \N__41201\,
            I => \N__41158\
        );

    \I__7393\ : InMux
    port map (
            O => \N__41198\,
            I => \N__41158\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__41195\,
            I => \N__41155\
        );

    \I__7391\ : InMux
    port map (
            O => \N__41194\,
            I => \N__41146\
        );

    \I__7390\ : InMux
    port map (
            O => \N__41193\,
            I => \N__41146\
        );

    \I__7389\ : InMux
    port map (
            O => \N__41192\,
            I => \N__41146\
        );

    \I__7388\ : InMux
    port map (
            O => \N__41191\,
            I => \N__41146\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__41188\,
            I => \N__41137\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__41185\,
            I => \N__41137\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__41182\,
            I => \N__41137\
        );

    \I__7384\ : Span4Mux_h
    port map (
            O => \N__41177\,
            I => \N__41137\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__41174\,
            I => \controlWord_6\
        );

    \I__7382\ : Odrv12
    port map (
            O => \N__41171\,
            I => \controlWord_6\
        );

    \I__7381\ : Odrv4
    port map (
            O => \N__41168\,
            I => \controlWord_6\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__41163\,
            I => \controlWord_6\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__41158\,
            I => \controlWord_6\
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__41155\,
            I => \controlWord_6\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__41146\,
            I => \controlWord_6\
        );

    \I__7376\ : Odrv4
    port map (
            O => \N__41137\,
            I => \controlWord_6\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__41120\,
            I => \CONTROL.un1_busState96_1_i_i_232_1_cascade_\
        );

    \I__7374\ : InMux
    port map (
            O => \N__41117\,
            I => \N__41114\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__41114\,
            I => \CONTROL.programCounter_ret_36_RNINU4NARZ0Z_7\
        );

    \I__7372\ : CascadeMux
    port map (
            O => \N__41111\,
            I => \PROM.ROMDATA.m23_cascade_\
        );

    \I__7371\ : InMux
    port map (
            O => \N__41108\,
            I => \N__41105\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__41105\,
            I => \N__41102\
        );

    \I__7369\ : Span4Mux_v
    port map (
            O => \N__41102\,
            I => \N__41097\
        );

    \I__7368\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41092\
        );

    \I__7367\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41092\
        );

    \I__7366\ : Span4Mux_h
    port map (
            O => \N__41097\,
            I => \N__41089\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__41092\,
            I => \N__41086\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__41089\,
            I => \PROM_ROMDATA_dintern_31_0__N_556_mux\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__41086\,
            I => \PROM_ROMDATA_dintern_31_0__N_556_mux\
        );

    \I__7362\ : InMux
    port map (
            O => \N__41081\,
            I => \N__41078\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__41078\,
            I => \N__41075\
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__41075\,
            I => \PROM.ROMDATA.m294_am\
        );

    \I__7359\ : CascadeMux
    port map (
            O => \N__41072\,
            I => \N__41069\
        );

    \I__7358\ : InMux
    port map (
            O => \N__41069\,
            I => \N__41066\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__41066\,
            I => \N__41063\
        );

    \I__7356\ : Span4Mux_h
    port map (
            O => \N__41063\,
            I => \N__41060\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__41060\,
            I => \PROM.ROMDATA.m271_1\
        );

    \I__7354\ : CascadeMux
    port map (
            O => \N__41057\,
            I => \PROM.ROMDATA.m271_1_cascade_\
        );

    \I__7353\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41046\
        );

    \I__7352\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41046\
        );

    \I__7351\ : InMux
    port map (
            O => \N__41052\,
            I => \N__41041\
        );

    \I__7350\ : InMux
    port map (
            O => \N__41051\,
            I => \N__41041\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__41046\,
            I => \N__41036\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__41041\,
            I => \N__41036\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__41036\,
            I => \N__41033\
        );

    \I__7346\ : Span4Mux_v
    port map (
            O => \N__41033\,
            I => \N__41030\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__41030\,
            I => \N__41027\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__41027\,
            I => \PROM.ROMDATA.m258_ns\
        );

    \I__7343\ : CascadeMux
    port map (
            O => \N__41024\,
            I => \PROM.ROMDATA.m258_ns_cascade_\
        );

    \I__7342\ : CascadeMux
    port map (
            O => \N__41021\,
            I => \PROM_ROMDATA_dintern_9ro_cascade_\
        );

    \I__7341\ : InMux
    port map (
            O => \N__41018\,
            I => \N__41015\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__41015\,
            I => \CONTROL.increment28lto5_1Z0Z_0\
        );

    \I__7339\ : CascadeMux
    port map (
            O => \N__41012\,
            I => \N__41009\
        );

    \I__7338\ : InMux
    port map (
            O => \N__41009\,
            I => \N__41005\
        );

    \I__7337\ : InMux
    port map (
            O => \N__41008\,
            I => \N__41002\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__41005\,
            I => \N__40999\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__41002\,
            I => \N__40996\
        );

    \I__7334\ : Span4Mux_v
    port map (
            O => \N__40999\,
            I => \N__40993\
        );

    \I__7333\ : Span4Mux_v
    port map (
            O => \N__40996\,
            I => \N__40988\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__40993\,
            I => \N__40988\
        );

    \I__7331\ : Odrv4
    port map (
            O => \N__40988\,
            I => \PROM.ROMDATA.N_566_mux\
        );

    \I__7330\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40982\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__40982\,
            I => \N__40979\
        );

    \I__7328\ : Span4Mux_v
    port map (
            O => \N__40979\,
            I => \N__40976\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__40976\,
            I => \N__40973\
        );

    \I__7326\ : Span4Mux_h
    port map (
            O => \N__40973\,
            I => \N__40970\
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__40970\,
            I => \PROM.ROMDATA.m470_bm\
        );

    \I__7324\ : CascadeMux
    port map (
            O => \N__40967\,
            I => \N__40964\
        );

    \I__7323\ : InMux
    port map (
            O => \N__40964\,
            I => \N__40959\
        );

    \I__7322\ : InMux
    port map (
            O => \N__40963\,
            I => \N__40955\
        );

    \I__7321\ : CascadeMux
    port map (
            O => \N__40962\,
            I => \N__40952\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__40959\,
            I => \N__40949\
        );

    \I__7319\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40946\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__40955\,
            I => \N__40943\
        );

    \I__7317\ : InMux
    port map (
            O => \N__40952\,
            I => \N__40940\
        );

    \I__7316\ : Span12Mux_h
    port map (
            O => \N__40949\,
            I => \N__40935\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__40946\,
            I => \N__40935\
        );

    \I__7314\ : Span4Mux_v
    port map (
            O => \N__40943\,
            I => \N__40930\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__40940\,
            I => \N__40930\
        );

    \I__7312\ : Odrv12
    port map (
            O => \N__40935\,
            I => \CONTROL.N_215\
        );

    \I__7311\ : Odrv4
    port map (
            O => \N__40930\,
            I => \CONTROL.N_215\
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__40925\,
            I => \N__40921\
        );

    \I__7309\ : CascadeMux
    port map (
            O => \N__40924\,
            I => \N__40917\
        );

    \I__7308\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40906\
        );

    \I__7307\ : InMux
    port map (
            O => \N__40920\,
            I => \N__40906\
        );

    \I__7306\ : InMux
    port map (
            O => \N__40917\,
            I => \N__40901\
        );

    \I__7305\ : InMux
    port map (
            O => \N__40916\,
            I => \N__40901\
        );

    \I__7304\ : InMux
    port map (
            O => \N__40915\,
            I => \N__40896\
        );

    \I__7303\ : InMux
    port map (
            O => \N__40914\,
            I => \N__40896\
        );

    \I__7302\ : InMux
    port map (
            O => \N__40913\,
            I => \N__40893\
        );

    \I__7301\ : InMux
    port map (
            O => \N__40912\,
            I => \N__40884\
        );

    \I__7300\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40884\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__40906\,
            I => \N__40881\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__40901\,
            I => \N__40878\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__40896\,
            I => \N__40875\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__40893\,
            I => \N__40872\
        );

    \I__7295\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40863\
        );

    \I__7294\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40863\
        );

    \I__7293\ : InMux
    port map (
            O => \N__40890\,
            I => \N__40863\
        );

    \I__7292\ : InMux
    port map (
            O => \N__40889\,
            I => \N__40863\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__40884\,
            I => \N__40860\
        );

    \I__7290\ : Span4Mux_v
    port map (
            O => \N__40881\,
            I => \N__40857\
        );

    \I__7289\ : Span4Mux_v
    port map (
            O => \N__40878\,
            I => \N__40850\
        );

    \I__7288\ : Span4Mux_v
    port map (
            O => \N__40875\,
            I => \N__40850\
        );

    \I__7287\ : Span4Mux_v
    port map (
            O => \N__40872\,
            I => \N__40850\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__40863\,
            I => \N__40847\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__40860\,
            I => \N__40844\
        );

    \I__7284\ : Sp12to4
    port map (
            O => \N__40857\,
            I => \N__40839\
        );

    \I__7283\ : Sp12to4
    port map (
            O => \N__40850\,
            I => \N__40839\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__40847\,
            I => \PROM.ROMDATA.dintern_12dfltZ0Z_0\
        );

    \I__7281\ : Odrv4
    port map (
            O => \N__40844\,
            I => \PROM.ROMDATA.dintern_12dfltZ0Z_0\
        );

    \I__7280\ : Odrv12
    port map (
            O => \N__40839\,
            I => \PROM.ROMDATA.dintern_12dfltZ0Z_0\
        );

    \I__7279\ : CascadeMux
    port map (
            O => \N__40832\,
            I => \PROM.ROMDATA.m284_cascade_\
        );

    \I__7278\ : CascadeMux
    port map (
            O => \N__40829\,
            I => \controlWord_12_cascade_\
        );

    \I__7277\ : InMux
    port map (
            O => \N__40826\,
            I => \N__40823\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__40823\,
            I => \N__40820\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__40820\,
            I => \N__40815\
        );

    \I__7274\ : InMux
    port map (
            O => \N__40819\,
            I => \N__40812\
        );

    \I__7273\ : InMux
    port map (
            O => \N__40818\,
            I => \N__40809\
        );

    \I__7272\ : Odrv4
    port map (
            O => \N__40815\,
            I => \CONTROL.increment28lto5_0\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__40812\,
            I => \CONTROL.increment28lto5_0\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__40809\,
            I => \CONTROL.increment28lto5_0\
        );

    \I__7269\ : CascadeMux
    port map (
            O => \N__40802\,
            I => \N__40797\
        );

    \I__7268\ : InMux
    port map (
            O => \N__40801\,
            I => \N__40787\
        );

    \I__7267\ : InMux
    port map (
            O => \N__40800\,
            I => \N__40787\
        );

    \I__7266\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40787\
        );

    \I__7265\ : InMux
    port map (
            O => \N__40796\,
            I => \N__40787\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__40787\,
            I => \N__40784\
        );

    \I__7263\ : Odrv12
    port map (
            O => \N__40784\,
            I => \PROM.ROMDATA.m273\
        );

    \I__7262\ : CascadeMux
    port map (
            O => \N__40781\,
            I => \PROM.ROMDATA.m273_cascade_\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__40778\,
            I => \PROM_ROMDATA_dintern_11ro_cascade_\
        );

    \I__7260\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40772\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__40772\,
            I => \CONTROL.increment28lto5_0_xZ0Z1\
        );

    \I__7258\ : InMux
    port map (
            O => \N__40769\,
            I => \N__40766\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__40766\,
            I => \CONTROL.increment28lto5_0_xZ0Z0\
        );

    \I__7256\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40757\
        );

    \I__7255\ : InMux
    port map (
            O => \N__40762\,
            I => \N__40757\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__40757\,
            I => \PROM_ROMDATA_dintern_11ro\
        );

    \I__7253\ : CascadeMux
    port map (
            O => \N__40754\,
            I => \N__40751\
        );

    \I__7252\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40746\
        );

    \I__7251\ : InMux
    port map (
            O => \N__40750\,
            I => \N__40741\
        );

    \I__7250\ : InMux
    port map (
            O => \N__40749\,
            I => \N__40741\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__40746\,
            I => \N__40736\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__40741\,
            I => \N__40736\
        );

    \I__7247\ : Span4Mux_h
    port map (
            O => \N__40736\,
            I => \N__40733\
        );

    \I__7246\ : Span4Mux_h
    port map (
            O => \N__40733\,
            I => \N__40730\
        );

    \I__7245\ : Span4Mux_h
    port map (
            O => \N__40730\,
            I => \N__40726\
        );

    \I__7244\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40723\
        );

    \I__7243\ : Span4Mux_v
    port map (
            O => \N__40726\,
            I => \N__40720\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__40723\,
            I => \aluStatus_4\
        );

    \I__7241\ : Odrv4
    port map (
            O => \N__40720\,
            I => \aluStatus_4\
        );

    \I__7240\ : InMux
    port map (
            O => \N__40715\,
            I => \N__40712\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__40712\,
            I => \controlWord_12\
        );

    \I__7238\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40706\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__40706\,
            I => \N__40703\
        );

    \I__7236\ : Span4Mux_h
    port map (
            O => \N__40703\,
            I => \N__40700\
        );

    \I__7235\ : Sp12to4
    port map (
            O => \N__40700\,
            I => \N__40697\
        );

    \I__7234\ : Span12Mux_v
    port map (
            O => \N__40697\,
            I => \N__40694\
        );

    \I__7233\ : Odrv12
    port map (
            O => \N__40694\,
            I => \CONTROL.g0_1_i_a6Z0Z_0\
        );

    \I__7232\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40688\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__40688\,
            I => \N__40685\
        );

    \I__7230\ : Span4Mux_h
    port map (
            O => \N__40685\,
            I => \N__40682\
        );

    \I__7229\ : Span4Mux_v
    port map (
            O => \N__40682\,
            I => \N__40679\
        );

    \I__7228\ : Odrv4
    port map (
            O => \N__40679\,
            I => \CONTROL.g0_1_i_a6Z0Z_1\
        );

    \I__7227\ : InMux
    port map (
            O => \N__40676\,
            I => \N__40673\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__40673\,
            I => \N__40670\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__40670\,
            I => \N__40667\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__40667\,
            I => \N__40664\
        );

    \I__7223\ : Span4Mux_h
    port map (
            O => \N__40664\,
            I => \N__40661\
        );

    \I__7222\ : Odrv4
    port map (
            O => \N__40661\,
            I => \CONTROL.g0_3_i_a7Z0Z_0\
        );

    \I__7221\ : CEMux
    port map (
            O => \N__40658\,
            I => \N__40654\
        );

    \I__7220\ : CEMux
    port map (
            O => \N__40657\,
            I => \N__40651\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__40654\,
            I => \N__40648\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__40651\,
            I => \N__40644\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__40648\,
            I => \N__40641\
        );

    \I__7216\ : CEMux
    port map (
            O => \N__40647\,
            I => \N__40638\
        );

    \I__7215\ : Span4Mux_v
    port map (
            O => \N__40644\,
            I => \N__40629\
        );

    \I__7214\ : Span4Mux_h
    port map (
            O => \N__40641\,
            I => \N__40629\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__40638\,
            I => \N__40629\
        );

    \I__7212\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40626\
        );

    \I__7211\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40622\
        );

    \I__7210\ : Span4Mux_h
    port map (
            O => \N__40629\,
            I => \N__40619\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__40626\,
            I => \N__40616\
        );

    \I__7208\ : InMux
    port map (
            O => \N__40625\,
            I => \N__40613\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__40622\,
            I => \N__40610\
        );

    \I__7206\ : Odrv4
    port map (
            O => \N__40619\,
            I => \CONTROL.aluReadBus_1_sqmuxa\
        );

    \I__7205\ : Odrv4
    port map (
            O => \N__40616\,
            I => \CONTROL.aluReadBus_1_sqmuxa\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__40613\,
            I => \CONTROL.aluReadBus_1_sqmuxa\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__40610\,
            I => \CONTROL.aluReadBus_1_sqmuxa\
        );

    \I__7202\ : InMux
    port map (
            O => \N__40601\,
            I => \N__40598\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__40598\,
            I => \N__40595\
        );

    \I__7200\ : Span4Mux_v
    port map (
            O => \N__40595\,
            I => \N__40589\
        );

    \I__7199\ : InMux
    port map (
            O => \N__40594\,
            I => \N__40586\
        );

    \I__7198\ : InMux
    port map (
            O => \N__40593\,
            I => \N__40582\
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__40592\,
            I => \N__40577\
        );

    \I__7196\ : Span4Mux_h
    port map (
            O => \N__40589\,
            I => \N__40571\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__40586\,
            I => \N__40571\
        );

    \I__7194\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40568\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__40582\,
            I => \N__40565\
        );

    \I__7192\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40560\
        );

    \I__7191\ : InMux
    port map (
            O => \N__40580\,
            I => \N__40560\
        );

    \I__7190\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40555\
        );

    \I__7189\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40555\
        );

    \I__7188\ : Span4Mux_h
    port map (
            O => \N__40571\,
            I => \N__40550\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__40568\,
            I => \N__40550\
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__40565\,
            I => \ALU.un14_log_a0_2Z0Z_15\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__40560\,
            I => \ALU.un14_log_a0_2Z0Z_15\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__40555\,
            I => \ALU.un14_log_a0_2Z0Z_15\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__40550\,
            I => \ALU.un14_log_a0_2Z0Z_15\
        );

    \I__7182\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40537\
        );

    \I__7181\ : InMux
    port map (
            O => \N__40540\,
            I => \N__40534\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__40537\,
            I => \N__40531\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__40534\,
            I => \N__40528\
        );

    \I__7178\ : Span4Mux_v
    port map (
            O => \N__40531\,
            I => \N__40523\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__40528\,
            I => \N__40523\
        );

    \I__7176\ : Odrv4
    port map (
            O => \N__40523\,
            I => \ALU.d_RNIN8NU4Z0Z_9\
        );

    \I__7175\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40517\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__40517\,
            I => \N__40514\
        );

    \I__7173\ : Span4Mux_v
    port map (
            O => \N__40514\,
            I => \N__40510\
        );

    \I__7172\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40507\
        );

    \I__7171\ : Span4Mux_h
    port map (
            O => \N__40510\,
            I => \N__40504\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__40507\,
            I => \ALU.combOperand2_0_0_9\
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__40504\,
            I => \ALU.combOperand2_0_0_9\
        );

    \I__7168\ : CascadeMux
    port map (
            O => \N__40499\,
            I => \N__40495\
        );

    \I__7167\ : InMux
    port map (
            O => \N__40498\,
            I => \N__40491\
        );

    \I__7166\ : InMux
    port map (
            O => \N__40495\,
            I => \N__40488\
        );

    \I__7165\ : CascadeMux
    port map (
            O => \N__40494\,
            I => \N__40485\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__40491\,
            I => \N__40480\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__40488\,
            I => \N__40480\
        );

    \I__7162\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40477\
        );

    \I__7161\ : Span4Mux_h
    port map (
            O => \N__40480\,
            I => \N__40474\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__40477\,
            I => \N__40471\
        );

    \I__7159\ : Span4Mux_h
    port map (
            O => \N__40474\,
            I => \N__40466\
        );

    \I__7158\ : Span4Mux_v
    port map (
            O => \N__40471\,
            I => \N__40466\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__40466\,
            I => \DROM_ROMDATA_dintern_9ro\
        );

    \I__7156\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40460\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__40460\,
            I => \N__40457\
        );

    \I__7154\ : Span4Mux_h
    port map (
            O => \N__40457\,
            I => \N__40454\
        );

    \I__7153\ : Span4Mux_v
    port map (
            O => \N__40454\,
            I => \N__40451\
        );

    \I__7152\ : Span4Mux_v
    port map (
            O => \N__40451\,
            I => \N__40448\
        );

    \I__7151\ : Span4Mux_v
    port map (
            O => \N__40448\,
            I => \N__40445\
        );

    \I__7150\ : Span4Mux_h
    port map (
            O => \N__40445\,
            I => \N__40442\
        );

    \I__7149\ : Span4Mux_h
    port map (
            O => \N__40442\,
            I => \N__40439\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__40439\,
            I => \N__40436\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__40436\,
            I => \gpuOut_c_9\
        );

    \I__7146\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40430\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__40430\,
            I => \N__40427\
        );

    \I__7144\ : Span4Mux_h
    port map (
            O => \N__40427\,
            I => \N__40424\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__40424\,
            I => \N__40421\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__40421\,
            I => \N__40418\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__40418\,
            I => \N__40415\
        );

    \I__7140\ : Span4Mux_v
    port map (
            O => \N__40415\,
            I => \N__40412\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__40412\,
            I => \N__40409\
        );

    \I__7138\ : IoSpan4Mux
    port map (
            O => \N__40409\,
            I => \N__40406\
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__40406\,
            I => \D9_in_c\
        );

    \I__7136\ : CascadeMux
    port map (
            O => \N__40403\,
            I => \CONTROL.N_170_cascade_\
        );

    \I__7135\ : InMux
    port map (
            O => \N__40400\,
            I => \N__40397\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__40397\,
            I => \N_186\
        );

    \I__7133\ : InMux
    port map (
            O => \N__40394\,
            I => \N__40391\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__40391\,
            I => \CONTROL.N_202\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__40388\,
            I => \N_186_cascade_\
        );

    \I__7130\ : IoInMux
    port map (
            O => \N__40385\,
            I => \N__40381\
        );

    \I__7129\ : IoInMux
    port map (
            O => \N__40384\,
            I => \N__40378\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__40381\,
            I => \N__40375\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__40378\,
            I => \N__40372\
        );

    \I__7126\ : IoSpan4Mux
    port map (
            O => \N__40375\,
            I => \N__40369\
        );

    \I__7125\ : IoSpan4Mux
    port map (
            O => \N__40372\,
            I => \N__40366\
        );

    \I__7124\ : Span4Mux_s1_h
    port map (
            O => \N__40369\,
            I => \N__40363\
        );

    \I__7123\ : Span4Mux_s2_h
    port map (
            O => \N__40366\,
            I => \N__40360\
        );

    \I__7122\ : Span4Mux_h
    port map (
            O => \N__40363\,
            I => \N__40357\
        );

    \I__7121\ : Span4Mux_h
    port map (
            O => \N__40360\,
            I => \N__40354\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__40357\,
            I => \N__40350\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__40354\,
            I => \N__40347\
        );

    \I__7118\ : InMux
    port map (
            O => \N__40353\,
            I => \N__40344\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__40350\,
            I => \N__40341\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__40347\,
            I => \N__40336\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__40344\,
            I => \N__40336\
        );

    \I__7114\ : Span4Mux_h
    port map (
            O => \N__40341\,
            I => \N__40333\
        );

    \I__7113\ : Span4Mux_v
    port map (
            O => \N__40336\,
            I => \N__40330\
        );

    \I__7112\ : Span4Mux_v
    port map (
            O => \N__40333\,
            I => \N__40325\
        );

    \I__7111\ : Span4Mux_v
    port map (
            O => \N__40330\,
            I => \N__40325\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__40325\,
            I => bus_9
        );

    \I__7109\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40319\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__40319\,
            I => \N__40316\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__40316\,
            I => \N__40313\
        );

    \I__7106\ : Span4Mux_v
    port map (
            O => \N__40313\,
            I => \N__40310\
        );

    \I__7105\ : Span4Mux_h
    port map (
            O => \N__40310\,
            I => \N__40306\
        );

    \I__7104\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40303\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__40306\,
            I => \CONTROL.ctrlOut_9\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__40303\,
            I => \CONTROL.ctrlOut_9\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__40298\,
            I => \N__40293\
        );

    \I__7100\ : InMux
    port map (
            O => \N__40297\,
            I => \N__40287\
        );

    \I__7099\ : InMux
    port map (
            O => \N__40296\,
            I => \N__40287\
        );

    \I__7098\ : InMux
    port map (
            O => \N__40293\,
            I => \N__40282\
        );

    \I__7097\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40282\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__40287\,
            I => \N__40279\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__40282\,
            I => \N__40276\
        );

    \I__7094\ : Span4Mux_v
    port map (
            O => \N__40279\,
            I => \N__40273\
        );

    \I__7093\ : Odrv4
    port map (
            O => \N__40276\,
            I => \PROM.ROMDATA.m284\
        );

    \I__7092\ : Odrv4
    port map (
            O => \N__40273\,
            I => \PROM.ROMDATA.m284\
        );

    \I__7091\ : InMux
    port map (
            O => \N__40268\,
            I => \N__40264\
        );

    \I__7090\ : CascadeMux
    port map (
            O => \N__40267\,
            I => \N__40261\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__40264\,
            I => \N__40258\
        );

    \I__7088\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40255\
        );

    \I__7087\ : Span4Mux_v
    port map (
            O => \N__40258\,
            I => \N__40252\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__40255\,
            I => \N__40249\
        );

    \I__7085\ : Span4Mux_h
    port map (
            O => \N__40252\,
            I => \N__40246\
        );

    \I__7084\ : Span4Mux_v
    port map (
            O => \N__40249\,
            I => \N__40243\
        );

    \I__7083\ : Span4Mux_v
    port map (
            O => \N__40246\,
            I => \N__40240\
        );

    \I__7082\ : Span4Mux_v
    port map (
            O => \N__40243\,
            I => \N__40236\
        );

    \I__7081\ : Span4Mux_v
    port map (
            O => \N__40240\,
            I => \N__40233\
        );

    \I__7080\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40230\
        );

    \I__7079\ : Span4Mux_h
    port map (
            O => \N__40236\,
            I => \N__40227\
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__40233\,
            I => h_5
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__40230\,
            I => h_5
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__40227\,
            I => h_5
        );

    \I__7075\ : InMux
    port map (
            O => \N__40220\,
            I => \N__40216\
        );

    \I__7074\ : InMux
    port map (
            O => \N__40219\,
            I => \N__40213\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__40216\,
            I => \N__40210\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__40213\,
            I => \N__40207\
        );

    \I__7071\ : Span12Mux_v
    port map (
            O => \N__40210\,
            I => \N__40204\
        );

    \I__7070\ : Span4Mux_h
    port map (
            O => \N__40207\,
            I => \N__40201\
        );

    \I__7069\ : Odrv12
    port map (
            O => \N__40204\,
            I => \ALU.dZ0Z_5\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__40201\,
            I => \ALU.dZ0Z_5\
        );

    \I__7067\ : InMux
    port map (
            O => \N__40196\,
            I => \N__40193\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__40193\,
            I => \ALU.d_RNIBT8EZ0Z_5\
        );

    \I__7065\ : CascadeMux
    port map (
            O => \N__40190\,
            I => \PROM.ROMDATA.m407_cascade_\
        );

    \I__7064\ : CascadeMux
    port map (
            O => \N__40187\,
            I => \PROM.ROMDATA.m488_ns_cascade_\
        );

    \I__7063\ : InMux
    port map (
            O => \N__40184\,
            I => \N__40181\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__40181\,
            I => \ALU.lshift_15_0_1\
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__40178\,
            I => \ALU.mult_1_cascade_\
        );

    \I__7060\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40172\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__40172\,
            I => \N__40169\
        );

    \I__7058\ : Span4Mux_v
    port map (
            O => \N__40169\,
            I => \N__40166\
        );

    \I__7057\ : Odrv4
    port map (
            O => \N__40166\,
            I => \ALU.a_15_m3_d_ns_1_1\
        );

    \I__7056\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40160\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__40160\,
            I => \N__40157\
        );

    \I__7054\ : Span4Mux_h
    port map (
            O => \N__40157\,
            I => \N__40154\
        );

    \I__7053\ : Span4Mux_v
    port map (
            O => \N__40154\,
            I => \N__40151\
        );

    \I__7052\ : Odrv4
    port map (
            O => \N__40151\,
            I => \ALU.d_RNIJOQE21Z0Z_0\
        );

    \I__7051\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40145\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__40145\,
            I => \N__40141\
        );

    \I__7049\ : InMux
    port map (
            O => \N__40144\,
            I => \N__40138\
        );

    \I__7048\ : Span4Mux_v
    port map (
            O => \N__40141\,
            I => \N__40135\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__40138\,
            I => \N__40131\
        );

    \I__7046\ : Span4Mux_h
    port map (
            O => \N__40135\,
            I => \N__40128\
        );

    \I__7045\ : InMux
    port map (
            O => \N__40134\,
            I => \N__40125\
        );

    \I__7044\ : Span4Mux_v
    port map (
            O => \N__40131\,
            I => \N__40122\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__40128\,
            I => \N__40119\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__40125\,
            I => \N__40116\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__40122\,
            I => \N__40113\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__40119\,
            I => \N__40108\
        );

    \I__7039\ : Span4Mux_h
    port map (
            O => \N__40116\,
            I => \N__40108\
        );

    \I__7038\ : Span4Mux_h
    port map (
            O => \N__40113\,
            I => \N__40105\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__40108\,
            I => \N__40102\
        );

    \I__7036\ : Odrv4
    port map (
            O => \N__40105\,
            I => g_5
        );

    \I__7035\ : Odrv4
    port map (
            O => \N__40102\,
            I => g_5
        );

    \I__7034\ : InMux
    port map (
            O => \N__40097\,
            I => \N__40094\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__40094\,
            I => \N__40091\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__40091\,
            I => \N__40087\
        );

    \I__7031\ : InMux
    port map (
            O => \N__40090\,
            I => \N__40084\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__40087\,
            I => \N__40081\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__40084\,
            I => \N__40078\
        );

    \I__7028\ : Span4Mux_h
    port map (
            O => \N__40081\,
            I => \N__40073\
        );

    \I__7027\ : Span4Mux_v
    port map (
            O => \N__40078\,
            I => \N__40073\
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__40073\,
            I => \ALU.cZ0Z_5\
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__40070\,
            I => \N__40066\
        );

    \I__7024\ : InMux
    port map (
            O => \N__40069\,
            I => \N__40063\
        );

    \I__7023\ : InMux
    port map (
            O => \N__40066\,
            I => \N__40060\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__40063\,
            I => \N__40057\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__40060\,
            I => \N__40054\
        );

    \I__7020\ : Span12Mux_h
    port map (
            O => \N__40057\,
            I => \N__40051\
        );

    \I__7019\ : Span4Mux_h
    port map (
            O => \N__40054\,
            I => \N__40048\
        );

    \I__7018\ : Odrv12
    port map (
            O => \N__40051\,
            I => \ALU.eZ0Z_5\
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__40048\,
            I => \ALU.eZ0Z_5\
        );

    \I__7016\ : InMux
    port map (
            O => \N__40043\,
            I => \N__40040\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__40040\,
            I => \N__40037\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__40037\,
            I => \N__40033\
        );

    \I__7013\ : InMux
    port map (
            O => \N__40036\,
            I => \N__40030\
        );

    \I__7012\ : Span4Mux_v
    port map (
            O => \N__40033\,
            I => \N__40027\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__40030\,
            I => \N__40024\
        );

    \I__7010\ : Span4Mux_h
    port map (
            O => \N__40027\,
            I => \N__40021\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__40024\,
            I => \N__40018\
        );

    \I__7008\ : Odrv4
    port map (
            O => \N__40021\,
            I => \ALU.aZ0Z_5\
        );

    \I__7007\ : Odrv4
    port map (
            O => \N__40018\,
            I => \ALU.aZ0Z_5\
        );

    \I__7006\ : InMux
    port map (
            O => \N__40013\,
            I => \N__40010\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__40010\,
            I => \ALU.c_RNI8KVQZ0Z_5\
        );

    \I__7004\ : CascadeMux
    port map (
            O => \N__40007\,
            I => \ALU.e_RNI48JMZ0Z_5_cascade_\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__40004\,
            I => \ALU.operand2_7_ns_1_5_cascade_\
        );

    \I__7002\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39998\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__39998\,
            I => \N__39995\
        );

    \I__7000\ : Span4Mux_v
    port map (
            O => \N__39995\,
            I => \N__39992\
        );

    \I__6999\ : Span4Mux_h
    port map (
            O => \N__39992\,
            I => \N__39989\
        );

    \I__6998\ : Odrv4
    port map (
            O => \N__39989\,
            I => \ALU.operand2_5\
        );

    \I__6997\ : InMux
    port map (
            O => \N__39986\,
            I => \N__39983\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__39983\,
            I => \N__39980\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__39980\,
            I => \N__39977\
        );

    \I__6994\ : Span4Mux_v
    port map (
            O => \N__39977\,
            I => \N__39974\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__39974\,
            I => \N__39969\
        );

    \I__6992\ : InMux
    port map (
            O => \N__39973\,
            I => \N__39966\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__39972\,
            I => \N__39963\
        );

    \I__6990\ : Span4Mux_v
    port map (
            O => \N__39969\,
            I => \N__39960\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__39966\,
            I => \N__39957\
        );

    \I__6988\ : InMux
    port map (
            O => \N__39963\,
            I => \N__39954\
        );

    \I__6987\ : Span4Mux_v
    port map (
            O => \N__39960\,
            I => \N__39949\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__39957\,
            I => \N__39949\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__39954\,
            I => \N__39946\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__39949\,
            I => \N__39943\
        );

    \I__6983\ : Span12Mux_v
    port map (
            O => \N__39946\,
            I => \N__39940\
        );

    \I__6982\ : Span4Mux_v
    port map (
            O => \N__39943\,
            I => \N__39937\
        );

    \I__6981\ : Odrv12
    port map (
            O => \N__39940\,
            I => f_5
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__39937\,
            I => f_5
        );

    \I__6979\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39929\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__39929\,
            I => \N__39926\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__39926\,
            I => \N__39923\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__39923\,
            I => \N__39919\
        );

    \I__6975\ : InMux
    port map (
            O => \N__39922\,
            I => \N__39916\
        );

    \I__6974\ : Sp12to4
    port map (
            O => \N__39919\,
            I => \N__39913\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__39916\,
            I => \N__39910\
        );

    \I__6972\ : Odrv12
    port map (
            O => \N__39913\,
            I => \ALU.bZ0Z_5\
        );

    \I__6971\ : Odrv12
    port map (
            O => \N__39910\,
            I => \ALU.bZ0Z_5\
        );

    \I__6970\ : InMux
    port map (
            O => \N__39905\,
            I => \N__39902\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__39902\,
            I => \ALU.b_RNI7HSPZ0Z_5\
        );

    \I__6968\ : InMux
    port map (
            O => \N__39899\,
            I => \N__39896\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__39896\,
            I => \N__39892\
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__39895\,
            I => \N__39889\
        );

    \I__6965\ : Span4Mux_v
    port map (
            O => \N__39892\,
            I => \N__39886\
        );

    \I__6964\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39883\
        );

    \I__6963\ : Sp12to4
    port map (
            O => \N__39886\,
            I => \N__39880\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__39883\,
            I => \N__39877\
        );

    \I__6961\ : Span12Mux_h
    port map (
            O => \N__39880\,
            I => \N__39874\
        );

    \I__6960\ : Span4Mux_h
    port map (
            O => \N__39877\,
            I => \N__39871\
        );

    \I__6959\ : Odrv12
    port map (
            O => \N__39874\,
            I => \ALU.bZ0Z_6\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__39871\,
            I => \ALU.bZ0Z_6\
        );

    \I__6957\ : InMux
    port map (
            O => \N__39866\,
            I => \N__39863\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__39863\,
            I => \N__39859\
        );

    \I__6955\ : InMux
    port map (
            O => \N__39862\,
            I => \N__39856\
        );

    \I__6954\ : Span4Mux_h
    port map (
            O => \N__39859\,
            I => \N__39851\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__39856\,
            I => \N__39851\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__39851\,
            I => \N__39848\
        );

    \I__6951\ : Sp12to4
    port map (
            O => \N__39848\,
            I => \N__39845\
        );

    \I__6950\ : Odrv12
    port map (
            O => \N__39845\,
            I => \ALU.bZ0Z_3\
        );

    \I__6949\ : InMux
    port map (
            O => \N__39842\,
            I => \N__39836\
        );

    \I__6948\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39836\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__39836\,
            I => \N__39833\
        );

    \I__6946\ : Span4Mux_h
    port map (
            O => \N__39833\,
            I => \N__39830\
        );

    \I__6945\ : Span4Mux_h
    port map (
            O => \N__39830\,
            I => \N__39827\
        );

    \I__6944\ : Sp12to4
    port map (
            O => \N__39827\,
            I => \N__39824\
        );

    \I__6943\ : Span12Mux_v
    port map (
            O => \N__39824\,
            I => \N__39821\
        );

    \I__6942\ : Odrv12
    port map (
            O => \N__39821\,
            I => \ALU.bZ0Z_11\
        );

    \I__6941\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39814\
        );

    \I__6940\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39811\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__39814\,
            I => \N__39808\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__39811\,
            I => \N__39805\
        );

    \I__6937\ : Span4Mux_v
    port map (
            O => \N__39808\,
            I => \N__39802\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__39805\,
            I => \N__39799\
        );

    \I__6935\ : Span4Mux_h
    port map (
            O => \N__39802\,
            I => \N__39796\
        );

    \I__6934\ : Span4Mux_h
    port map (
            O => \N__39799\,
            I => \N__39793\
        );

    \I__6933\ : Span4Mux_h
    port map (
            O => \N__39796\,
            I => \N__39790\
        );

    \I__6932\ : Sp12to4
    port map (
            O => \N__39793\,
            I => \N__39787\
        );

    \I__6931\ : Sp12to4
    port map (
            O => \N__39790\,
            I => \N__39782\
        );

    \I__6930\ : Span12Mux_s7_h
    port map (
            O => \N__39787\,
            I => \N__39782\
        );

    \I__6929\ : Odrv12
    port map (
            O => \N__39782\,
            I => \ALU.bZ0Z_12\
        );

    \I__6928\ : InMux
    port map (
            O => \N__39779\,
            I => \N__39776\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__39776\,
            I => \N__39773\
        );

    \I__6926\ : Span4Mux_v
    port map (
            O => \N__39773\,
            I => \N__39770\
        );

    \I__6925\ : Span4Mux_v
    port map (
            O => \N__39770\,
            I => \N__39767\
        );

    \I__6924\ : Odrv4
    port map (
            O => \N__39767\,
            I => \CONTROL.gZ0Z3\
        );

    \I__6923\ : InMux
    port map (
            O => \N__39764\,
            I => \N__39761\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__39761\,
            I => \N__39758\
        );

    \I__6921\ : Span4Mux_v
    port map (
            O => \N__39758\,
            I => \N__39755\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__39755\,
            I => \ALU.lshift_15_0_sx_1\
        );

    \I__6919\ : IoInMux
    port map (
            O => \N__39752\,
            I => \N__39748\
        );

    \I__6918\ : IoInMux
    port map (
            O => \N__39751\,
            I => \N__39745\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__39748\,
            I => \N__39742\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__39745\,
            I => \N__39739\
        );

    \I__6915\ : Span4Mux_s0_h
    port map (
            O => \N__39742\,
            I => \N__39736\
        );

    \I__6914\ : IoSpan4Mux
    port map (
            O => \N__39739\,
            I => \N__39733\
        );

    \I__6913\ : Sp12to4
    port map (
            O => \N__39736\,
            I => \N__39729\
        );

    \I__6912\ : Sp12to4
    port map (
            O => \N__39733\,
            I => \N__39726\
        );

    \I__6911\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39723\
        );

    \I__6910\ : Span12Mux_v
    port map (
            O => \N__39729\,
            I => \N__39720\
        );

    \I__6909\ : Span12Mux_s7_h
    port map (
            O => \N__39726\,
            I => \N__39715\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__39723\,
            I => \N__39715\
        );

    \I__6907\ : Span12Mux_h
    port map (
            O => \N__39720\,
            I => \N__39710\
        );

    \I__6906\ : Span12Mux_h
    port map (
            O => \N__39715\,
            I => \N__39710\
        );

    \I__6905\ : Odrv12
    port map (
            O => \N__39710\,
            I => bus_14
        );

    \I__6904\ : CascadeMux
    port map (
            O => \N__39707\,
            I => \ALU.lshift_15_0_1_cascade_\
        );

    \I__6903\ : InMux
    port map (
            O => \N__39704\,
            I => \N__39701\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__39701\,
            I => \ALU.a_15_m0_sx_14\
        );

    \I__6901\ : InMux
    port map (
            O => \N__39698\,
            I => \N__39695\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__39695\,
            I => \ALU.c_RNI890LZ0Z_13\
        );

    \I__6899\ : CascadeMux
    port map (
            O => \N__39692\,
            I => \ALU.a_RNI4P741Z0Z_13_cascade_\
        );

    \I__6898\ : InMux
    port map (
            O => \N__39689\,
            I => \N__39686\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__39686\,
            I => \ALU.d_RNIAHCTZ0Z_13\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__39683\,
            I => \ALU.operand2_7_ns_1_13_cascade_\
        );

    \I__6895\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39677\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__39677\,
            I => \ALU.b_RNI61KC1Z0Z_13\
        );

    \I__6893\ : InMux
    port map (
            O => \N__39674\,
            I => \N__39671\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__39671\,
            I => \N__39668\
        );

    \I__6891\ : Span4Mux_h
    port map (
            O => \N__39668\,
            I => \N__39665\
        );

    \I__6890\ : Span4Mux_h
    port map (
            O => \N__39665\,
            I => \N__39662\
        );

    \I__6889\ : Span4Mux_v
    port map (
            O => \N__39662\,
            I => \N__39659\
        );

    \I__6888\ : Odrv4
    port map (
            O => \N__39659\,
            I => \ALU.operand2_13\
        );

    \I__6887\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39653\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__39653\,
            I => \N__39648\
        );

    \I__6885\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39645\
        );

    \I__6884\ : InMux
    port map (
            O => \N__39651\,
            I => \N__39642\
        );

    \I__6883\ : Span4Mux_v
    port map (
            O => \N__39648\,
            I => \N__39637\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__39645\,
            I => \N__39637\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__39642\,
            I => \N__39634\
        );

    \I__6880\ : Span4Mux_v
    port map (
            O => \N__39637\,
            I => \N__39631\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__39634\,
            I => \N__39628\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__39631\,
            I => \N__39625\
        );

    \I__6877\ : Span4Mux_v
    port map (
            O => \N__39628\,
            I => \N__39622\
        );

    \I__6876\ : Span4Mux_h
    port map (
            O => \N__39625\,
            I => \N__39619\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__39622\,
            I => bus_0_13
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__39619\,
            I => bus_0_13
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__39614\,
            I => \ALU.operand2_13_cascade_\
        );

    \I__6872\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39608\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__39608\,
            I => \N__39600\
        );

    \I__6870\ : InMux
    port map (
            O => \N__39607\,
            I => \N__39595\
        );

    \I__6869\ : InMux
    port map (
            O => \N__39606\,
            I => \N__39592\
        );

    \I__6868\ : InMux
    port map (
            O => \N__39605\,
            I => \N__39589\
        );

    \I__6867\ : InMux
    port map (
            O => \N__39604\,
            I => \N__39586\
        );

    \I__6866\ : InMux
    port map (
            O => \N__39603\,
            I => \N__39583\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__39600\,
            I => \N__39580\
        );

    \I__6864\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39577\
        );

    \I__6863\ : InMux
    port map (
            O => \N__39598\,
            I => \N__39574\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__39595\,
            I => \N__39571\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__39592\,
            I => \N__39568\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__39589\,
            I => \N__39565\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__39586\,
            I => \N__39558\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__39583\,
            I => \N__39558\
        );

    \I__6857\ : Span4Mux_v
    port map (
            O => \N__39580\,
            I => \N__39558\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__39577\,
            I => \N__39551\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__39574\,
            I => \N__39551\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__39571\,
            I => \N__39551\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__39568\,
            I => \N__39544\
        );

    \I__6852\ : Span4Mux_v
    port map (
            O => \N__39565\,
            I => \N__39544\
        );

    \I__6851\ : Span4Mux_h
    port map (
            O => \N__39558\,
            I => \N__39544\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__39551\,
            I => \ALU.d_RNI02EVNBZ0Z_4\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__39544\,
            I => \ALU.d_RNI02EVNBZ0Z_4\
        );

    \I__6848\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39536\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__39536\,
            I => \N__39532\
        );

    \I__6846\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39527\
        );

    \I__6845\ : Span4Mux_h
    port map (
            O => \N__39532\,
            I => \N__39524\
        );

    \I__6844\ : InMux
    port map (
            O => \N__39531\,
            I => \N__39521\
        );

    \I__6843\ : InMux
    port map (
            O => \N__39530\,
            I => \N__39518\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__39527\,
            I => \N__39511\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__39524\,
            I => \N__39504\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__39521\,
            I => \N__39504\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__39518\,
            I => \N__39504\
        );

    \I__6838\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39501\
        );

    \I__6837\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39498\
        );

    \I__6836\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39495\
        );

    \I__6835\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39492\
        );

    \I__6834\ : Odrv4
    port map (
            O => \N__39511\,
            I => \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__39504\,
            I => \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__39501\,
            I => \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__39498\,
            I => \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__39495\,
            I => \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__39492\,
            I => \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\
        );

    \I__6828\ : InMux
    port map (
            O => \N__39479\,
            I => \N__39476\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__39476\,
            I => \N__39472\
        );

    \I__6826\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39469\
        );

    \I__6825\ : Span4Mux_v
    port map (
            O => \N__39472\,
            I => \N__39465\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__39469\,
            I => \N__39462\
        );

    \I__6823\ : InMux
    port map (
            O => \N__39468\,
            I => \N__39459\
        );

    \I__6822\ : Span4Mux_h
    port map (
            O => \N__39465\,
            I => \N__39450\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__39462\,
            I => \N__39450\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__39459\,
            I => \N__39447\
        );

    \I__6819\ : InMux
    port map (
            O => \N__39458\,
            I => \N__39444\
        );

    \I__6818\ : InMux
    port map (
            O => \N__39457\,
            I => \N__39441\
        );

    \I__6817\ : InMux
    port map (
            O => \N__39456\,
            I => \N__39438\
        );

    \I__6816\ : InMux
    port map (
            O => \N__39455\,
            I => \N__39435\
        );

    \I__6815\ : Odrv4
    port map (
            O => \N__39450\,
            I => \ALU.addsub_cry_1_c_RNIICPECZ0Z7\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__39447\,
            I => \ALU.addsub_cry_1_c_RNIICPECZ0Z7\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__39444\,
            I => \ALU.addsub_cry_1_c_RNIICPECZ0Z7\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__39441\,
            I => \ALU.addsub_cry_1_c_RNIICPECZ0Z7\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__39438\,
            I => \ALU.addsub_cry_1_c_RNIICPECZ0Z7\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__39435\,
            I => \ALU.addsub_cry_1_c_RNIICPECZ0Z7\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__39422\,
            I => \N__39419\
        );

    \I__6808\ : InMux
    port map (
            O => \N__39419\,
            I => \N__39416\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__39416\,
            I => \N__39412\
        );

    \I__6806\ : InMux
    port map (
            O => \N__39415\,
            I => \N__39409\
        );

    \I__6805\ : Span4Mux_v
    port map (
            O => \N__39412\,
            I => \N__39404\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__39409\,
            I => \N__39404\
        );

    \I__6803\ : Span4Mux_h
    port map (
            O => \N__39404\,
            I => \N__39401\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__39401\,
            I => \N__39398\
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__39398\,
            I => \ALU.bZ0Z_2\
        );

    \I__6800\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39388\
        );

    \I__6799\ : InMux
    port map (
            O => \N__39394\,
            I => \N__39384\
        );

    \I__6798\ : InMux
    port map (
            O => \N__39393\,
            I => \N__39381\
        );

    \I__6797\ : InMux
    port map (
            O => \N__39392\,
            I => \N__39378\
        );

    \I__6796\ : InMux
    port map (
            O => \N__39391\,
            I => \N__39374\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__39388\,
            I => \N__39371\
        );

    \I__6794\ : InMux
    port map (
            O => \N__39387\,
            I => \N__39368\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__39384\,
            I => \N__39365\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__39381\,
            I => \N__39360\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__39378\,
            I => \N__39360\
        );

    \I__6790\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39357\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__39374\,
            I => \N__39354\
        );

    \I__6788\ : Span4Mux_v
    port map (
            O => \N__39371\,
            I => \N__39351\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__39368\,
            I => \N__39346\
        );

    \I__6786\ : Span4Mux_v
    port map (
            O => \N__39365\,
            I => \N__39346\
        );

    \I__6785\ : Span4Mux_v
    port map (
            O => \N__39360\,
            I => \N__39343\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__39357\,
            I => \N__39340\
        );

    \I__6783\ : Span4Mux_v
    port map (
            O => \N__39354\,
            I => \N__39335\
        );

    \I__6782\ : Span4Mux_h
    port map (
            O => \N__39351\,
            I => \N__39335\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__39346\,
            I => \N__39330\
        );

    \I__6780\ : Span4Mux_h
    port map (
            O => \N__39343\,
            I => \N__39330\
        );

    \I__6779\ : Odrv4
    port map (
            O => \N__39340\,
            I => \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9\
        );

    \I__6778\ : Odrv4
    port map (
            O => \N__39335\,
            I => \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9\
        );

    \I__6777\ : Odrv4
    port map (
            O => \N__39330\,
            I => \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9\
        );

    \I__6776\ : InMux
    port map (
            O => \N__39323\,
            I => \N__39316\
        );

    \I__6775\ : InMux
    port map (
            O => \N__39322\,
            I => \N__39311\
        );

    \I__6774\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39308\
        );

    \I__6773\ : InMux
    port map (
            O => \N__39320\,
            I => \N__39305\
        );

    \I__6772\ : InMux
    port map (
            O => \N__39319\,
            I => \N__39302\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__39316\,
            I => \N__39298\
        );

    \I__6770\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39295\
        );

    \I__6769\ : InMux
    port map (
            O => \N__39314\,
            I => \N__39292\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__39311\,
            I => \N__39289\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__39308\,
            I => \N__39286\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__39305\,
            I => \N__39283\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__39302\,
            I => \N__39280\
        );

    \I__6764\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39277\
        );

    \I__6763\ : Span4Mux_h
    port map (
            O => \N__39298\,
            I => \N__39274\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__39295\,
            I => \N__39265\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__39292\,
            I => \N__39265\
        );

    \I__6760\ : Span4Mux_h
    port map (
            O => \N__39289\,
            I => \N__39265\
        );

    \I__6759\ : Span4Mux_v
    port map (
            O => \N__39286\,
            I => \N__39265\
        );

    \I__6758\ : Span4Mux_h
    port map (
            O => \N__39283\,
            I => \N__39260\
        );

    \I__6757\ : Span4Mux_h
    port map (
            O => \N__39280\,
            I => \N__39260\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__39277\,
            I => \ALU.addsub_cry_4_c_RNI5L6IQAZ0\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__39274\,
            I => \ALU.addsub_cry_4_c_RNI5L6IQAZ0\
        );

    \I__6754\ : Odrv4
    port map (
            O => \N__39265\,
            I => \ALU.addsub_cry_4_c_RNI5L6IQAZ0\
        );

    \I__6753\ : Odrv4
    port map (
            O => \N__39260\,
            I => \ALU.addsub_cry_4_c_RNI5L6IQAZ0\
        );

    \I__6752\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39248\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__39248\,
            I => \N__39245\
        );

    \I__6750\ : Span4Mux_v
    port map (
            O => \N__39245\,
            I => \N__39241\
        );

    \I__6749\ : InMux
    port map (
            O => \N__39244\,
            I => \N__39238\
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__39241\,
            I => \ALU.N_1025\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__39238\,
            I => \ALU.N_1025\
        );

    \I__6746\ : InMux
    port map (
            O => \N__39233\,
            I => \N__39230\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__39230\,
            I => \N__39226\
        );

    \I__6744\ : InMux
    port map (
            O => \N__39229\,
            I => \N__39223\
        );

    \I__6743\ : Span4Mux_h
    port map (
            O => \N__39226\,
            I => \N__39218\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__39223\,
            I => \N__39218\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__39218\,
            I => \N__39215\
        );

    \I__6740\ : Odrv4
    port map (
            O => \N__39215\,
            I => \ALU.N_864\
        );

    \I__6739\ : CascadeMux
    port map (
            O => \N__39212\,
            I => \ALU.N_965_cascade_\
        );

    \I__6738\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39206\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__39206\,
            I => \N__39203\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__39203\,
            I => \ALU.d_RNIFHCRU4Z0Z_2\
        );

    \I__6735\ : InMux
    port map (
            O => \N__39200\,
            I => \N__39197\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__39197\,
            I => \N__39194\
        );

    \I__6733\ : Span4Mux_v
    port map (
            O => \N__39194\,
            I => \N__39191\
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__39191\,
            I => \ALU.mult_15_15\
        );

    \I__6731\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39185\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__39185\,
            I => \ALU.c_RNINT9PO2Z0Z_10\
        );

    \I__6729\ : InMux
    port map (
            O => \N__39182\,
            I => \N__39179\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__39179\,
            I => \ALU.mult_13\
        );

    \I__6727\ : InMux
    port map (
            O => \N__39176\,
            I => \N__39172\
        );

    \I__6726\ : InMux
    port map (
            O => \N__39175\,
            I => \N__39169\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__39172\,
            I => \N__39166\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__39169\,
            I => \N__39163\
        );

    \I__6723\ : Span4Mux_h
    port map (
            O => \N__39166\,
            I => \N__39160\
        );

    \I__6722\ : Span4Mux_h
    port map (
            O => \N__39163\,
            I => \N__39155\
        );

    \I__6721\ : Span4Mux_h
    port map (
            O => \N__39160\,
            I => \N__39155\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__39155\,
            I => \ALU.N_642\
        );

    \I__6719\ : CascadeMux
    port map (
            O => \N__39152\,
            I => \ALU.d_RNIULN025Z0Z_2_cascade_\
        );

    \I__6718\ : InMux
    port map (
            O => \N__39149\,
            I => \N__39146\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__39146\,
            I => \ALU.d_RNIULN025_0Z0Z_2\
        );

    \I__6716\ : CascadeMux
    port map (
            O => \N__39143\,
            I => \ALU.lshift_10_cascade_\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__39140\,
            I => \ALU.c_RNIO0KOKEZ0Z_10_cascade_\
        );

    \I__6714\ : InMux
    port map (
            O => \N__39137\,
            I => \N__39134\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__39134\,
            I => \N__39130\
        );

    \I__6712\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39127\
        );

    \I__6711\ : Span4Mux_v
    port map (
            O => \N__39130\,
            I => \N__39122\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__39127\,
            I => \N__39122\
        );

    \I__6709\ : Span4Mux_h
    port map (
            O => \N__39122\,
            I => \N__39119\
        );

    \I__6708\ : Span4Mux_h
    port map (
            O => \N__39119\,
            I => \N__39116\
        );

    \I__6707\ : Sp12to4
    port map (
            O => \N__39116\,
            I => \N__39113\
        );

    \I__6706\ : Span12Mux_v
    port map (
            O => \N__39113\,
            I => \N__39110\
        );

    \I__6705\ : Span12Mux_h
    port map (
            O => \N__39110\,
            I => \N__39107\
        );

    \I__6704\ : Odrv12
    port map (
            O => \N__39107\,
            I => \ALU.bZ0Z_10\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__39104\,
            I => \ALU.lshift_3_ns_1_15_cascade_\
        );

    \I__6702\ : InMux
    port map (
            O => \N__39101\,
            I => \N__39097\
        );

    \I__6701\ : InMux
    port map (
            O => \N__39100\,
            I => \N__39092\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__39097\,
            I => \N__39083\
        );

    \I__6699\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39078\
        );

    \I__6698\ : InMux
    port map (
            O => \N__39095\,
            I => \N__39078\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__39092\,
            I => \N__39075\
        );

    \I__6696\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39068\
        );

    \I__6695\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39068\
        );

    \I__6694\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39068\
        );

    \I__6693\ : InMux
    port map (
            O => \N__39088\,
            I => \N__39061\
        );

    \I__6692\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39061\
        );

    \I__6691\ : InMux
    port map (
            O => \N__39086\,
            I => \N__39061\
        );

    \I__6690\ : Span4Mux_h
    port map (
            O => \N__39083\,
            I => \N__39058\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__39078\,
            I => \ALU.d_RNI64MA6Z0Z_0\
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__39075\,
            I => \ALU.d_RNI64MA6Z0Z_0\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__39068\,
            I => \ALU.d_RNI64MA6Z0Z_0\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__39061\,
            I => \ALU.d_RNI64MA6Z0Z_0\
        );

    \I__6685\ : Odrv4
    port map (
            O => \N__39058\,
            I => \ALU.d_RNI64MA6Z0Z_0\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__39047\,
            I => \N__39041\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__39046\,
            I => \N__39037\
        );

    \I__6682\ : CascadeMux
    port map (
            O => \N__39045\,
            I => \N__39034\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__39044\,
            I => \N__39031\
        );

    \I__6680\ : InMux
    port map (
            O => \N__39041\,
            I => \N__39028\
        );

    \I__6679\ : InMux
    port map (
            O => \N__39040\,
            I => \N__39020\
        );

    \I__6678\ : InMux
    port map (
            O => \N__39037\,
            I => \N__39013\
        );

    \I__6677\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39013\
        );

    \I__6676\ : InMux
    port map (
            O => \N__39031\,
            I => \N__39013\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__39028\,
            I => \N__39010\
        );

    \I__6674\ : InMux
    port map (
            O => \N__39027\,
            I => \N__39005\
        );

    \I__6673\ : InMux
    port map (
            O => \N__39026\,
            I => \N__39005\
        );

    \I__6672\ : InMux
    port map (
            O => \N__39025\,
            I => \N__38998\
        );

    \I__6671\ : InMux
    port map (
            O => \N__39024\,
            I => \N__38998\
        );

    \I__6670\ : InMux
    port map (
            O => \N__39023\,
            I => \N__38998\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__39020\,
            I => \N__38993\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__39013\,
            I => \N__38993\
        );

    \I__6667\ : Span4Mux_h
    port map (
            O => \N__39010\,
            I => \N__38990\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__39005\,
            I => \N_225_0\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__38998\,
            I => \N_225_0\
        );

    \I__6664\ : Odrv4
    port map (
            O => \N__38993\,
            I => \N_225_0\
        );

    \I__6663\ : Odrv4
    port map (
            O => \N__38990\,
            I => \N_225_0\
        );

    \I__6662\ : InMux
    port map (
            O => \N__38981\,
            I => \N__38978\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__38978\,
            I => \N__38974\
        );

    \I__6660\ : CascadeMux
    port map (
            O => \N__38977\,
            I => \N__38971\
        );

    \I__6659\ : Span4Mux_v
    port map (
            O => \N__38974\,
            I => \N__38968\
        );

    \I__6658\ : InMux
    port map (
            O => \N__38971\,
            I => \N__38965\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__38968\,
            I => \ALU.mult_25_12\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__38965\,
            I => \ALU.mult_25_12\
        );

    \I__6655\ : CascadeMux
    port map (
            O => \N__38960\,
            I => \ALU.mult_13_12_cascade_\
        );

    \I__6654\ : InMux
    port map (
            O => \N__38957\,
            I => \N__38954\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__38954\,
            I => \ALU.mult_467_c_RNICRDK6BZ0\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__38951\,
            I => \N__38948\
        );

    \I__6651\ : InMux
    port map (
            O => \N__38948\,
            I => \N__38945\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__38945\,
            I => \ALU.mult_13_12\
        );

    \I__6649\ : CascadeMux
    port map (
            O => \N__38942\,
            I => \N__38939\
        );

    \I__6648\ : InMux
    port map (
            O => \N__38939\,
            I => \N__38936\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__38936\,
            I => \N__38933\
        );

    \I__6646\ : Odrv12
    port map (
            O => \N__38933\,
            I => \ALU.mult_13_13\
        );

    \I__6645\ : CascadeMux
    port map (
            O => \N__38930\,
            I => \N__38927\
        );

    \I__6644\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38924\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__38924\,
            I => \ALU.mult_27_13\
        );

    \I__6642\ : InMux
    port map (
            O => \N__38921\,
            I => \ALU.mult_27_c12\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__38918\,
            I => \N__38915\
        );

    \I__6640\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38912\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__38912\,
            I => \ALU.mult_365_c_RNI8ALOZ0Z96\
        );

    \I__6638\ : CascadeMux
    port map (
            O => \N__38909\,
            I => \N__38906\
        );

    \I__6637\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38903\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__38903\,
            I => \ALU.mult_27_14\
        );

    \I__6635\ : InMux
    port map (
            O => \N__38900\,
            I => \ALU.mult_27_c13\
        );

    \I__6634\ : InMux
    port map (
            O => \N__38897\,
            I => \ALU.mult_27_c14\
        );

    \I__6633\ : CascadeMux
    port map (
            O => \N__38894\,
            I => \N__38891\
        );

    \I__6632\ : InMux
    port map (
            O => \N__38891\,
            I => \N__38888\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__38888\,
            I => \N__38885\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__38885\,
            I => \ALU.mult_27_c14_THRU_CO\
        );

    \I__6629\ : CascadeMux
    port map (
            O => \N__38882\,
            I => \N__38879\
        );

    \I__6628\ : InMux
    port map (
            O => \N__38879\,
            I => \N__38876\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__38876\,
            I => \ALU.mult_9\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__38873\,
            I => \N__38870\
        );

    \I__6625\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38864\
        );

    \I__6624\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38864\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__38864\,
            I => \N__38861\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__38861\,
            I => \N__38858\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__38858\,
            I => \PROM.ROMDATA.m382_ns\
        );

    \I__6620\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38852\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__38852\,
            I => \N__38849\
        );

    \I__6618\ : Span12Mux_v
    port map (
            O => \N__38849\,
            I => \N__38844\
        );

    \I__6617\ : InMux
    port map (
            O => \N__38848\,
            I => \N__38839\
        );

    \I__6616\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38839\
        );

    \I__6615\ : Odrv12
    port map (
            O => \N__38844\,
            I => \busState_1_RNIAR0U1_2\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__38839\,
            I => \busState_1_RNIAR0U1_2\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__38834\,
            I => \N_225_0_cascade_\
        );

    \I__6612\ : InMux
    port map (
            O => \N__38831\,
            I => \N__38828\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__38828\,
            I => \ALU.mult_13_15\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__38825\,
            I => \ALU.mult_15_14_cascade_\
        );

    \I__6609\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38818\
        );

    \I__6608\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38815\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__38818\,
            I => \ALU.mult_13_14\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__38815\,
            I => \ALU.mult_13_14\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__38810\,
            I => \N__38807\
        );

    \I__6604\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38804\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__38804\,
            I => \CONTROL.N_304_0\
        );

    \I__6602\ : InMux
    port map (
            O => \N__38801\,
            I => \N__38795\
        );

    \I__6601\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38795\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__38795\,
            I => \N__38792\
        );

    \I__6599\ : Span4Mux_h
    port map (
            O => \N__38792\,
            I => \N__38789\
        );

    \I__6598\ : Span4Mux_h
    port map (
            O => \N__38789\,
            I => \N__38786\
        );

    \I__6597\ : Sp12to4
    port map (
            O => \N__38786\,
            I => \N__38783\
        );

    \I__6596\ : Odrv12
    port map (
            O => \N__38783\,
            I => \PROM.ROMDATA.m433_ns\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__38780\,
            I => \PROM.ROMDATA.m294_bm_cascade_\
        );

    \I__6594\ : CascadeMux
    port map (
            O => \N__38777\,
            I => \PROM.ROMDATA.m31_cascade_\
        );

    \I__6593\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38771\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__38771\,
            I => \N__38768\
        );

    \I__6591\ : Span4Mux_v
    port map (
            O => \N__38768\,
            I => \N__38765\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__38765\,
            I => \N__38761\
        );

    \I__6589\ : InMux
    port map (
            O => \N__38764\,
            I => \N__38758\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__38761\,
            I => \CONTROL.ctrlOut_12\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__38758\,
            I => \CONTROL.ctrlOut_12\
        );

    \I__6586\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38750\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__38750\,
            I => \CONTROL.dout_reto_12\
        );

    \I__6584\ : CascadeMux
    port map (
            O => \N__38747\,
            I => \PROM.ROMDATA.m391_cascade_\
        );

    \I__6583\ : InMux
    port map (
            O => \N__38744\,
            I => \N__38741\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__38741\,
            I => \PROM.ROMDATA.m433_bm\
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__38738\,
            I => \controlWord_4_cascade_\
        );

    \I__6580\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38731\
        );

    \I__6579\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38728\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__38731\,
            I => \CONTROL.N_5_0\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__38728\,
            I => \CONTROL.N_5_0\
        );

    \I__6576\ : InMux
    port map (
            O => \N__38723\,
            I => \N__38720\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__38720\,
            I => \CONTROL.g0_12_1\
        );

    \I__6574\ : InMux
    port map (
            O => \N__38717\,
            I => \N__38710\
        );

    \I__6573\ : InMux
    port map (
            O => \N__38716\,
            I => \N__38707\
        );

    \I__6572\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38700\
        );

    \I__6571\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38700\
        );

    \I__6570\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38700\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__38710\,
            I => \N__38696\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__38707\,
            I => \N__38693\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__38700\,
            I => \N__38690\
        );

    \I__6566\ : InMux
    port map (
            O => \N__38699\,
            I => \N__38687\
        );

    \I__6565\ : Span4Mux_h
    port map (
            O => \N__38696\,
            I => \N__38684\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__38693\,
            I => \N__38679\
        );

    \I__6563\ : Span4Mux_v
    port map (
            O => \N__38690\,
            I => \N__38679\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__38687\,
            I => \N__38675\
        );

    \I__6561\ : Span4Mux_v
    port map (
            O => \N__38684\,
            I => \N__38672\
        );

    \I__6560\ : Span4Mux_h
    port map (
            O => \N__38679\,
            I => \N__38669\
        );

    \I__6559\ : InMux
    port map (
            O => \N__38678\,
            I => \N__38666\
        );

    \I__6558\ : Odrv12
    port map (
            O => \N__38675\,
            I => \CONTROL.N_360\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__38672\,
            I => \CONTROL.N_360\
        );

    \I__6556\ : Odrv4
    port map (
            O => \N__38669\,
            I => \CONTROL.N_360\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__38666\,
            I => \CONTROL.N_360\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__38657\,
            I => \N__38654\
        );

    \I__6553\ : InMux
    port map (
            O => \N__38654\,
            I => \N__38651\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__38651\,
            I => \N__38648\
        );

    \I__6551\ : Span4Mux_h
    port map (
            O => \N__38648\,
            I => \N__38645\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__38645\,
            I => \N__38641\
        );

    \I__6549\ : InMux
    port map (
            O => \N__38644\,
            I => \N__38638\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__38641\,
            I => \CONTROL.N_362\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__38638\,
            I => \CONTROL.N_362\
        );

    \I__6546\ : InMux
    port map (
            O => \N__38633\,
            I => \N__38630\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__38627\,
            I => \CONTROL.m28_0_120_i_i_0\
        );

    \I__6543\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38620\
        );

    \I__6542\ : InMux
    port map (
            O => \N__38623\,
            I => \N__38617\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__38620\,
            I => \N__38614\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__38617\,
            I => \N__38611\
        );

    \I__6539\ : Odrv12
    port map (
            O => \N__38614\,
            I => \CONTROL.N_321\
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__38611\,
            I => \CONTROL.N_321\
        );

    \I__6537\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38603\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__38603\,
            I => \N__38600\
        );

    \I__6535\ : Odrv12
    port map (
            O => \N__38600\,
            I => \CONTROL.N_338\
        );

    \I__6534\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38588\
        );

    \I__6533\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38588\
        );

    \I__6532\ : InMux
    port map (
            O => \N__38595\,
            I => \N__38588\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__38588\,
            I => \N__38585\
        );

    \I__6530\ : Span4Mux_v
    port map (
            O => \N__38585\,
            I => \N__38576\
        );

    \I__6529\ : InMux
    port map (
            O => \N__38584\,
            I => \N__38571\
        );

    \I__6528\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38571\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__38582\,
            I => \N__38568\
        );

    \I__6526\ : InMux
    port map (
            O => \N__38581\,
            I => \N__38559\
        );

    \I__6525\ : InMux
    port map (
            O => \N__38580\,
            I => \N__38559\
        );

    \I__6524\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38559\
        );

    \I__6523\ : Span4Mux_h
    port map (
            O => \N__38576\,
            I => \N__38556\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38553\
        );

    \I__6521\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38550\
        );

    \I__6520\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38545\
        );

    \I__6519\ : InMux
    port map (
            O => \N__38566\,
            I => \N__38545\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__38559\,
            I => \N__38542\
        );

    \I__6517\ : Odrv4
    port map (
            O => \N__38556\,
            I => \PROM_ROMDATA_dintern_0ro\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__38553\,
            I => \PROM_ROMDATA_dintern_0ro\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__38550\,
            I => \PROM_ROMDATA_dintern_0ro\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__38545\,
            I => \PROM_ROMDATA_dintern_0ro\
        );

    \I__6513\ : Odrv4
    port map (
            O => \N__38542\,
            I => \PROM_ROMDATA_dintern_0ro\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__38531\,
            I => \PROM_ROMDATA_dintern_0ro_cascade_\
        );

    \I__6511\ : CascadeMux
    port map (
            O => \N__38528\,
            I => \N__38525\
        );

    \I__6510\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38522\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__38522\,
            I => \N__38519\
        );

    \I__6508\ : Odrv12
    port map (
            O => \N__38519\,
            I => \CONTROL.un1_busState_0_sqmuxa_i_a2_0\
        );

    \I__6507\ : InMux
    port map (
            O => \N__38516\,
            I => \N__38513\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__38513\,
            I => \N__38510\
        );

    \I__6505\ : Span12Mux_s11_v
    port map (
            O => \N__38510\,
            I => \N__38507\
        );

    \I__6504\ : Odrv12
    port map (
            O => \N__38507\,
            I => \CONTROL.N_133_0_1\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__38504\,
            I => \PROM_ROMDATA_dintern_3ro_cascade_\
        );

    \I__6502\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38498\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__38498\,
            I => \N__38495\
        );

    \I__6500\ : Span4Mux_h
    port map (
            O => \N__38495\,
            I => \N__38492\
        );

    \I__6499\ : Span4Mux_h
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__38489\,
            I => \CONTROL.g0_3_i_2_0\
        );

    \I__6497\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38483\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__38483\,
            I => \N__38480\
        );

    \I__6495\ : Odrv12
    port map (
            O => \N__38480\,
            I => \CONTROL.g0_2_i_a7Z0Z_3\
        );

    \I__6494\ : InMux
    port map (
            O => \N__38477\,
            I => \N__38474\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__38474\,
            I => \CONTROL.g0_2_i_a7Z0Z_2\
        );

    \I__6492\ : CascadeMux
    port map (
            O => \N__38471\,
            I => \CONTROL.g0_2_i_2_cascade_\
        );

    \I__6491\ : InMux
    port map (
            O => \N__38468\,
            I => \N__38465\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__38465\,
            I => \N__38462\
        );

    \I__6489\ : Span4Mux_v
    port map (
            O => \N__38462\,
            I => \N__38458\
        );

    \I__6488\ : CascadeMux
    port map (
            O => \N__38461\,
            I => \N__38455\
        );

    \I__6487\ : Span4Mux_h
    port map (
            O => \N__38458\,
            I => \N__38452\
        );

    \I__6486\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38449\
        );

    \I__6485\ : Odrv4
    port map (
            O => \N__38452\,
            I => \CONTROL.addrstack_1_2\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__38449\,
            I => \CONTROL.addrstack_1_2\
        );

    \I__6483\ : InMux
    port map (
            O => \N__38444\,
            I => \N__38438\
        );

    \I__6482\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38432\
        );

    \I__6481\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38432\
        );

    \I__6480\ : InMux
    port map (
            O => \N__38441\,
            I => \N__38428\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__38438\,
            I => \N__38425\
        );

    \I__6478\ : InMux
    port map (
            O => \N__38437\,
            I => \N__38422\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__38432\,
            I => \N__38419\
        );

    \I__6476\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38416\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__38428\,
            I => \N__38412\
        );

    \I__6474\ : Span4Mux_v
    port map (
            O => \N__38425\,
            I => \N__38408\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__38422\,
            I => \N__38405\
        );

    \I__6472\ : Span4Mux_v
    port map (
            O => \N__38419\,
            I => \N__38400\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38400\
        );

    \I__6470\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38397\
        );

    \I__6469\ : Span4Mux_v
    port map (
            O => \N__38412\,
            I => \N__38394\
        );

    \I__6468\ : InMux
    port map (
            O => \N__38411\,
            I => \N__38391\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__38408\,
            I => \N__38384\
        );

    \I__6466\ : Span4Mux_h
    port map (
            O => \N__38405\,
            I => \N__38384\
        );

    \I__6465\ : Span4Mux_h
    port map (
            O => \N__38400\,
            I => \N__38384\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__38397\,
            I => \CONTROL.addrstackptrZ0Z_1\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__38394\,
            I => \CONTROL.addrstackptrZ0Z_1\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__38391\,
            I => \CONTROL.addrstackptrZ0Z_1\
        );

    \I__6461\ : Odrv4
    port map (
            O => \N__38384\,
            I => \CONTROL.addrstackptrZ0Z_1\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__38375\,
            I => \CONTROL.N_5_0_cascade_\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__38372\,
            I => \CONTROL.g0_12_1_cascade_\
        );

    \I__6458\ : CascadeMux
    port map (
            O => \N__38369\,
            I => \N__38366\
        );

    \I__6457\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38363\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__38363\,
            I => \N__38360\
        );

    \I__6455\ : Span12Mux_h
    port map (
            O => \N__38360\,
            I => \N__38357\
        );

    \I__6454\ : Odrv12
    port map (
            O => \N__38357\,
            I => \CONTROL.addrstackptr_8_2\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__38354\,
            I => \controlWord_6_cascade_\
        );

    \I__6452\ : InMux
    port map (
            O => \N__38351\,
            I => \N__38348\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__38348\,
            I => \CONTROL.N_140_0\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__38345\,
            I => \CONTROL.un1_busState96_1_i_i_a2_1Z0Z_1_cascade_\
        );

    \I__6449\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38339\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__38339\,
            I => \CONTROL.un1_busState96_1_i_i_a2_0Z0Z_1\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__38336\,
            I => \CONTROL.un1_busState96_1_i_iZ0Z_0_cascade_\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__38333\,
            I => \controlWord_5_cascade_\
        );

    \I__6445\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38327\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__38327\,
            I => \CONTROL.N_134_0\
        );

    \I__6443\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38320\
        );

    \I__6442\ : InMux
    port map (
            O => \N__38323\,
            I => \N__38317\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__38320\,
            I => \N__38314\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__38317\,
            I => \N__38309\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__38314\,
            I => \N__38309\
        );

    \I__6438\ : Span4Mux_h
    port map (
            O => \N__38309\,
            I => \N__38306\
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__38306\,
            I => \CONTROL.N_327\
        );

    \I__6436\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38300\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__38300\,
            I => \N__38297\
        );

    \I__6434\ : Span4Mux_v
    port map (
            O => \N__38297\,
            I => \N__38294\
        );

    \I__6433\ : Span4Mux_v
    port map (
            O => \N__38294\,
            I => \N__38291\
        );

    \I__6432\ : Span4Mux_v
    port map (
            O => \N__38291\,
            I => \N__38288\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__38288\,
            I => \ALU.status_RNO_2Z0Z_0\
        );

    \I__6430\ : CascadeMux
    port map (
            O => \N__38285\,
            I => \N__38282\
        );

    \I__6429\ : InMux
    port map (
            O => \N__38282\,
            I => \N__38279\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__38279\,
            I => \ALU.status_e_1_0\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__38276\,
            I => \CONTROL.increment28lto5_1Z0Z_1_cascade_\
        );

    \I__6426\ : InMux
    port map (
            O => \N__38273\,
            I => \N__38269\
        );

    \I__6425\ : InMux
    port map (
            O => \N__38272\,
            I => \N__38266\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__38269\,
            I => \N__38261\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__38266\,
            I => \N__38258\
        );

    \I__6422\ : InMux
    port map (
            O => \N__38265\,
            I => \N__38253\
        );

    \I__6421\ : InMux
    port map (
            O => \N__38264\,
            I => \N__38253\
        );

    \I__6420\ : Span4Mux_v
    port map (
            O => \N__38261\,
            I => \N__38250\
        );

    \I__6419\ : Span4Mux_v
    port map (
            O => \N__38258\,
            I => \N__38244\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__38253\,
            I => \N__38241\
        );

    \I__6417\ : Span4Mux_h
    port map (
            O => \N__38250\,
            I => \N__38238\
        );

    \I__6416\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38231\
        );

    \I__6415\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38231\
        );

    \I__6414\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38231\
        );

    \I__6413\ : Span4Mux_h
    port map (
            O => \N__38244\,
            I => \N__38226\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__38241\,
            I => \N__38226\
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__38238\,
            I => \PROM_ROMDATA_dintern_8ro\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__38231\,
            I => \PROM_ROMDATA_dintern_8ro\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__38226\,
            I => \PROM_ROMDATA_dintern_8ro\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__38219\,
            I => \CONTROL.increment28lto5_1_1_2_cascade_\
        );

    \I__6407\ : InMux
    port map (
            O => \N__38216\,
            I => \N__38213\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__38213\,
            I => \N__38210\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__38210\,
            I => \N__38206\
        );

    \I__6404\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38201\
        );

    \I__6403\ : Span4Mux_h
    port map (
            O => \N__38206\,
            I => \N__38198\
        );

    \I__6402\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38193\
        );

    \I__6401\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38193\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__38201\,
            I => \PROM_ROMDATA_dintern_7ro\
        );

    \I__6399\ : Odrv4
    port map (
            O => \N__38198\,
            I => \PROM_ROMDATA_dintern_7ro\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__38193\,
            I => \PROM_ROMDATA_dintern_7ro\
        );

    \I__6397\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38181\
        );

    \I__6396\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38178\
        );

    \I__6395\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38175\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__38181\,
            I => \N__38172\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__38178\,
            I => \N__38167\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__38175\,
            I => \N__38167\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__38172\,
            I => \N__38164\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__38167\,
            I => \N__38161\
        );

    \I__6389\ : Span4Mux_h
    port map (
            O => \N__38164\,
            I => \N__38157\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__38161\,
            I => \N__38154\
        );

    \I__6387\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38151\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__38157\,
            I => \CONTROL.increment28lto5_1Z0Z_2\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__38154\,
            I => \CONTROL.increment28lto5_1Z0Z_2\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__38151\,
            I => \CONTROL.increment28lto5_1Z0Z_2\
        );

    \I__6383\ : CEMux
    port map (
            O => \N__38144\,
            I => \N__38141\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__38141\,
            I => \N__38137\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__38140\,
            I => \N__38134\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__38137\,
            I => \N__38131\
        );

    \I__6379\ : InMux
    port map (
            O => \N__38134\,
            I => \N__38128\
        );

    \I__6378\ : Span4Mux_h
    port map (
            O => \N__38131\,
            I => \N__38122\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__38128\,
            I => \N__38119\
        );

    \I__6376\ : InMux
    port map (
            O => \N__38127\,
            I => \N__38116\
        );

    \I__6375\ : CEMux
    port map (
            O => \N__38126\,
            I => \N__38113\
        );

    \I__6374\ : CEMux
    port map (
            O => \N__38125\,
            I => \N__38110\
        );

    \I__6373\ : Sp12to4
    port map (
            O => \N__38122\,
            I => \N__38105\
        );

    \I__6372\ : Span12Mux_v
    port map (
            O => \N__38119\,
            I => \N__38105\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__38116\,
            I => \N__38102\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__38113\,
            I => \CONTROL.N_48_0\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__38110\,
            I => \CONTROL.N_48_0\
        );

    \I__6368\ : Odrv12
    port map (
            O => \N__38105\,
            I => \CONTROL.N_48_0\
        );

    \I__6367\ : Odrv4
    port map (
            O => \N__38102\,
            I => \CONTROL.N_48_0\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__38093\,
            I => \ALU.N_1200_cascade_\
        );

    \I__6365\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38087\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__38087\,
            I => \ALU.N_1248\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__38084\,
            I => \ALU.d_RNIGMEO4Z0Z_3_cascade_\
        );

    \I__6362\ : InMux
    port map (
            O => \N__38081\,
            I => \N__38078\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__38078\,
            I => \N__38075\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__38075\,
            I => \N__38072\
        );

    \I__6359\ : Span4Mux_h
    port map (
            O => \N__38072\,
            I => \N__38069\
        );

    \I__6358\ : Odrv4
    port map (
            O => \N__38069\,
            I => \ALU.combOperand2_d_bmZ0Z_3\
        );

    \I__6357\ : InMux
    port map (
            O => \N__38066\,
            I => \N__38062\
        );

    \I__6356\ : InMux
    port map (
            O => \N__38065\,
            I => \N__38059\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__38062\,
            I => \N__38054\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__38059\,
            I => \N__38051\
        );

    \I__6353\ : InMux
    port map (
            O => \N__38058\,
            I => \N__38046\
        );

    \I__6352\ : InMux
    port map (
            O => \N__38057\,
            I => \N__38046\
        );

    \I__6351\ : Span4Mux_v
    port map (
            O => \N__38054\,
            I => \N__38043\
        );

    \I__6350\ : Span4Mux_v
    port map (
            O => \N__38051\,
            I => \N__38040\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__38046\,
            I => \N__38037\
        );

    \I__6348\ : Span4Mux_h
    port map (
            O => \N__38043\,
            I => \N__38032\
        );

    \I__6347\ : Span4Mux_h
    port map (
            O => \N__38040\,
            I => \N__38032\
        );

    \I__6346\ : Odrv12
    port map (
            O => \N__38037\,
            I => \ALU.d_RNI2CUG6Z0Z_3\
        );

    \I__6345\ : Odrv4
    port map (
            O => \N__38032\,
            I => \ALU.d_RNI2CUG6Z0Z_3\
        );

    \I__6344\ : InMux
    port map (
            O => \N__38027\,
            I => \N__38024\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__38024\,
            I => \N__38021\
        );

    \I__6342\ : Span4Mux_v
    port map (
            O => \N__38021\,
            I => \N__38018\
        );

    \I__6341\ : Span4Mux_v
    port map (
            O => \N__38018\,
            I => \N__38015\
        );

    \I__6340\ : Span4Mux_v
    port map (
            O => \N__38015\,
            I => \N__38012\
        );

    \I__6339\ : Span4Mux_v
    port map (
            O => \N__38012\,
            I => \N__38009\
        );

    \I__6338\ : Span4Mux_h
    port map (
            O => \N__38009\,
            I => \N__38006\
        );

    \I__6337\ : Span4Mux_h
    port map (
            O => \N__38006\,
            I => \N__38003\
        );

    \I__6336\ : Span4Mux_h
    port map (
            O => \N__38003\,
            I => \N__38000\
        );

    \I__6335\ : Span4Mux_h
    port map (
            O => \N__38000\,
            I => \N__37997\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__37997\,
            I => \gpuOut_c_4\
        );

    \I__6333\ : InMux
    port map (
            O => \N__37994\,
            I => \N__37990\
        );

    \I__6332\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37987\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__37990\,
            I => \N__37984\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__37987\,
            I => \N__37981\
        );

    \I__6329\ : Span4Mux_h
    port map (
            O => \N__37984\,
            I => \N__37978\
        );

    \I__6328\ : Span4Mux_v
    port map (
            O => \N__37981\,
            I => \N__37973\
        );

    \I__6327\ : Span4Mux_v
    port map (
            O => \N__37978\,
            I => \N__37973\
        );

    \I__6326\ : Odrv4
    port map (
            O => \N__37973\,
            I => \CONTROL.N_165\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__37970\,
            I => \N__37967\
        );

    \I__6324\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37964\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__37964\,
            I => \N__37961\
        );

    \I__6322\ : Span4Mux_v
    port map (
            O => \N__37961\,
            I => \N__37957\
        );

    \I__6321\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37954\
        );

    \I__6320\ : Span4Mux_v
    port map (
            O => \N__37957\,
            I => \N__37951\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__37954\,
            I => \N__37948\
        );

    \I__6318\ : Sp12to4
    port map (
            O => \N__37951\,
            I => \N__37945\
        );

    \I__6317\ : Span4Mux_h
    port map (
            O => \N__37948\,
            I => \N__37942\
        );

    \I__6316\ : Span12Mux_h
    port map (
            O => \N__37945\,
            I => \N__37938\
        );

    \I__6315\ : Span4Mux_h
    port map (
            O => \N__37942\,
            I => \N__37935\
        );

    \I__6314\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37932\
        );

    \I__6313\ : Odrv12
    port map (
            O => \N__37938\,
            I => h_9
        );

    \I__6312\ : Odrv4
    port map (
            O => \N__37935\,
            I => h_9
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__37932\,
            I => h_9
        );

    \I__6310\ : InMux
    port map (
            O => \N__37925\,
            I => \N__37922\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__37922\,
            I => \N__37919\
        );

    \I__6308\ : Odrv4
    port map (
            O => \N__37919\,
            I => \ALU.e_RNICGJMZ0Z_9\
        );

    \I__6307\ : InMux
    port map (
            O => \N__37916\,
            I => \N__37913\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__37913\,
            I => \ALU.d_RNIKKNJZ0Z_9\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__37910\,
            I => \ALU.operand2_7_ns_1_9_cascade_\
        );

    \I__6304\ : InMux
    port map (
            O => \N__37907\,
            I => \N__37904\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__37904\,
            I => \ALU.b_RNIG8BVZ0Z_9\
        );

    \I__6302\ : CascadeMux
    port map (
            O => \N__37901\,
            I => \ALU.operand2_9_cascade_\
        );

    \I__6301\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37895\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__37895\,
            I => \ALU.e_RNI933SZ0Z_0\
        );

    \I__6299\ : CascadeMux
    port map (
            O => \N__37892\,
            I => \ALU.c_RNIDFF01Z0Z_0_cascade_\
        );

    \I__6298\ : InMux
    port map (
            O => \N__37889\,
            I => \N__37886\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__37886\,
            I => \ALU.d_RNI0G5DZ0Z_0\
        );

    \I__6296\ : CascadeMux
    port map (
            O => \N__37883\,
            I => \ALU.b_RNIS3POZ0Z_0_cascade_\
        );

    \I__6295\ : InMux
    port map (
            O => \N__37880\,
            I => \N__37877\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__37877\,
            I => \ALU.operand2_7_ns_1_0\
        );

    \I__6293\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37871\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__37871\,
            I => \N__37867\
        );

    \I__6291\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37864\
        );

    \I__6290\ : Span4Mux_v
    port map (
            O => \N__37867\,
            I => \N__37861\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__37864\,
            I => \N__37858\
        );

    \I__6288\ : Span4Mux_v
    port map (
            O => \N__37861\,
            I => \N__37853\
        );

    \I__6287\ : Span4Mux_h
    port map (
            O => \N__37858\,
            I => \N__37853\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__37853\,
            I => \ALU.operand2_0\
        );

    \I__6285\ : InMux
    port map (
            O => \N__37850\,
            I => \N__37847\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__37847\,
            I => \N__37844\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__37844\,
            I => \N__37840\
        );

    \I__6282\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37837\
        );

    \I__6281\ : Span4Mux_v
    port map (
            O => \N__37840\,
            I => \N__37832\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__37837\,
            I => \N__37832\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__37832\,
            I => \ALU.dZ0Z_3\
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__37829\,
            I => \ALU.operand2_6_ns_1_3_cascade_\
        );

    \I__6277\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37823\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__37823\,
            I => \N__37819\
        );

    \I__6275\ : InMux
    port map (
            O => \N__37822\,
            I => \N__37816\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__37819\,
            I => \N__37813\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__37816\,
            I => \N__37810\
        );

    \I__6272\ : Span4Mux_v
    port map (
            O => \N__37813\,
            I => \N__37807\
        );

    \I__6271\ : Odrv12
    port map (
            O => \N__37810\,
            I => \ALU.aZ0Z_3\
        );

    \I__6270\ : Odrv4
    port map (
            O => \N__37807\,
            I => \ALU.aZ0Z_3\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__37802\,
            I => \N__37798\
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__37801\,
            I => \N__37795\
        );

    \I__6267\ : InMux
    port map (
            O => \N__37798\,
            I => \N__37792\
        );

    \I__6266\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37789\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__37792\,
            I => \N__37786\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__37789\,
            I => \N__37783\
        );

    \I__6263\ : Span4Mux_h
    port map (
            O => \N__37786\,
            I => \N__37780\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__37783\,
            I => \N__37777\
        );

    \I__6261\ : Span4Mux_h
    port map (
            O => \N__37780\,
            I => \N__37774\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__37777\,
            I => \ALU.eZ0Z_3\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__37774\,
            I => \ALU.eZ0Z_3\
        );

    \I__6258\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37765\
        );

    \I__6257\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37762\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__37765\,
            I => \N__37759\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__37762\,
            I => \N__37756\
        );

    \I__6254\ : Span4Mux_v
    port map (
            O => \N__37759\,
            I => \N__37753\
        );

    \I__6253\ : Sp12to4
    port map (
            O => \N__37756\,
            I => \N__37750\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__37753\,
            I => \ALU.cZ0Z_3\
        );

    \I__6251\ : Odrv12
    port map (
            O => \N__37750\,
            I => \ALU.cZ0Z_3\
        );

    \I__6250\ : InMux
    port map (
            O => \N__37745\,
            I => \N__37742\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__37742\,
            I => \N__37738\
        );

    \I__6248\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37734\
        );

    \I__6247\ : Span4Mux_v
    port map (
            O => \N__37738\,
            I => \N__37731\
        );

    \I__6246\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37728\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__37734\,
            I => \N__37725\
        );

    \I__6244\ : Span4Mux_v
    port map (
            O => \N__37731\,
            I => \N__37722\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37719\
        );

    \I__6242\ : Span4Mux_v
    port map (
            O => \N__37725\,
            I => \N__37716\
        );

    \I__6241\ : Span4Mux_v
    port map (
            O => \N__37722\,
            I => \N__37713\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__37719\,
            I => \N__37710\
        );

    \I__6239\ : Span4Mux_h
    port map (
            O => \N__37716\,
            I => \N__37707\
        );

    \I__6238\ : Span4Mux_h
    port map (
            O => \N__37713\,
            I => \N__37702\
        );

    \I__6237\ : Span4Mux_v
    port map (
            O => \N__37710\,
            I => \N__37702\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__37707\,
            I => \N__37699\
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__37702\,
            I => g_3
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__37699\,
            I => g_3
        );

    \I__6233\ : CascadeMux
    port map (
            O => \N__37694\,
            I => \ALU.operand2_3_ns_1_3_cascade_\
        );

    \I__6232\ : CascadeMux
    port map (
            O => \N__37691\,
            I => \ALU.a_15_m2_d_d_ns_1_0_0_cascade_\
        );

    \I__6231\ : IoInMux
    port map (
            O => \N__37688\,
            I => \N__37685\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__37685\,
            I => \N__37681\
        );

    \I__6229\ : IoInMux
    port map (
            O => \N__37684\,
            I => \N__37678\
        );

    \I__6228\ : IoSpan4Mux
    port map (
            O => \N__37681\,
            I => \N__37675\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__37678\,
            I => \N__37672\
        );

    \I__6226\ : IoSpan4Mux
    port map (
            O => \N__37675\,
            I => \N__37669\
        );

    \I__6225\ : IoSpan4Mux
    port map (
            O => \N__37672\,
            I => \N__37666\
        );

    \I__6224\ : Sp12to4
    port map (
            O => \N__37669\,
            I => \N__37663\
        );

    \I__6223\ : Span4Mux_s0_h
    port map (
            O => \N__37666\,
            I => \N__37660\
        );

    \I__6222\ : Span12Mux_s7_h
    port map (
            O => \N__37663\,
            I => \N__37656\
        );

    \I__6221\ : Sp12to4
    port map (
            O => \N__37660\,
            I => \N__37653\
        );

    \I__6220\ : InMux
    port map (
            O => \N__37659\,
            I => \N__37650\
        );

    \I__6219\ : Span12Mux_h
    port map (
            O => \N__37656\,
            I => \N__37645\
        );

    \I__6218\ : Span12Mux_h
    port map (
            O => \N__37653\,
            I => \N__37645\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__37650\,
            I => \N__37642\
        );

    \I__6216\ : Odrv12
    port map (
            O => \N__37645\,
            I => bus_0
        );

    \I__6215\ : Odrv12
    port map (
            O => \N__37642\,
            I => bus_0
        );

    \I__6214\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37633\
        );

    \I__6213\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37630\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__37633\,
            I => \N__37627\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__37630\,
            I => \N__37624\
        );

    \I__6210\ : Span4Mux_v
    port map (
            O => \N__37627\,
            I => \N__37621\
        );

    \I__6209\ : Span4Mux_v
    port map (
            O => \N__37624\,
            I => \N__37618\
        );

    \I__6208\ : Span4Mux_h
    port map (
            O => \N__37621\,
            I => \N__37615\
        );

    \I__6207\ : Span4Mux_h
    port map (
            O => \N__37618\,
            I => \N__37612\
        );

    \I__6206\ : Span4Mux_v
    port map (
            O => \N__37615\,
            I => \N__37609\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__37612\,
            I => \ALU.lshift62\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__37609\,
            I => \ALU.lshift62\
        );

    \I__6203\ : CascadeMux
    port map (
            O => \N__37604\,
            I => \ALU.d_RNI4D6E01Z0Z_0_cascade_\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__37601\,
            I => \ALU.d_RNIQQ9O83Z0Z_0_cascade_\
        );

    \I__6201\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37595\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__37595\,
            I => \ALU.d_RNI4HL061Z0Z_0\
        );

    \I__6199\ : CascadeMux
    port map (
            O => \N__37592\,
            I => \ALU.d_RNINUGCF4Z0Z_0_cascade_\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__37589\,
            I => \N__37586\
        );

    \I__6197\ : InMux
    port map (
            O => \N__37586\,
            I => \N__37583\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__37583\,
            I => \N__37580\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__37580\,
            I => \N__37576\
        );

    \I__6194\ : InMux
    port map (
            O => \N__37579\,
            I => \N__37573\
        );

    \I__6193\ : Span4Mux_h
    port map (
            O => \N__37576\,
            I => \N__37570\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__37573\,
            I => \ALU.aZ0Z_0\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__37570\,
            I => \ALU.aZ0Z_0\
        );

    \I__6190\ : InMux
    port map (
            O => \N__37565\,
            I => \N__37562\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__37562\,
            I => \N__37558\
        );

    \I__6188\ : CascadeMux
    port map (
            O => \N__37561\,
            I => \N__37555\
        );

    \I__6187\ : Span4Mux_v
    port map (
            O => \N__37558\,
            I => \N__37552\
        );

    \I__6186\ : InMux
    port map (
            O => \N__37555\,
            I => \N__37549\
        );

    \I__6185\ : Span4Mux_h
    port map (
            O => \N__37552\,
            I => \N__37543\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__37549\,
            I => \N__37543\
        );

    \I__6183\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37540\
        );

    \I__6182\ : Span4Mux_h
    port map (
            O => \N__37543\,
            I => \N__37537\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__37540\,
            I => h_0
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__37537\,
            I => h_0
        );

    \I__6179\ : InMux
    port map (
            O => \N__37532\,
            I => \N__37528\
        );

    \I__6178\ : InMux
    port map (
            O => \N__37531\,
            I => \N__37525\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__37528\,
            I => \ALU.a_15_am_snZ0Z_11\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__37525\,
            I => \ALU.a_15_am_snZ0Z_11\
        );

    \I__6175\ : InMux
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__37517\,
            I => \N__37513\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__37516\,
            I => \N__37509\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__37513\,
            I => \N__37506\
        );

    \I__6171\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37503\
        );

    \I__6170\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37500\
        );

    \I__6169\ : Span4Mux_h
    port map (
            O => \N__37506\,
            I => \N__37495\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__37503\,
            I => \N__37495\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__37500\,
            I => \N__37492\
        );

    \I__6166\ : Span4Mux_h
    port map (
            O => \N__37495\,
            I => \N__37487\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__37492\,
            I => \N__37487\
        );

    \I__6164\ : Span4Mux_v
    port map (
            O => \N__37487\,
            I => \N__37484\
        );

    \I__6163\ : Span4Mux_h
    port map (
            O => \N__37484\,
            I => \N__37481\
        );

    \I__6162\ : Odrv4
    port map (
            O => \N__37481\,
            I => h_1
        );

    \I__6161\ : InMux
    port map (
            O => \N__37478\,
            I => \N__37475\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__37475\,
            I => \N__37472\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__37469\,
            I => \ALU.mult_6\
        );

    \I__6157\ : CascadeMux
    port map (
            O => \N__37466\,
            I => \ALU.mult_489_c_RNIGEUL1AZ0_cascade_\
        );

    \I__6156\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37460\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__37460\,
            I => \ALU.mult_489_c_RNIGEUL1AZ0\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__37457\,
            I => \ALU.mult_489_c_RNIPGBQMCZ0Z_0_cascade_\
        );

    \I__6153\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37451\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__37451\,
            I => \ALU.mult_489_c_RNIPGBQMCZ0\
        );

    \I__6151\ : CascadeMux
    port map (
            O => \N__37448\,
            I => \ALU.mult_489_c_RNI1J3GCUZ0_cascade_\
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__6149\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37439\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__37439\,
            I => \N__37435\
        );

    \I__6147\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37431\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__37435\,
            I => \N__37428\
        );

    \I__6145\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37425\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__37431\,
            I => \N__37422\
        );

    \I__6143\ : Span4Mux_v
    port map (
            O => \N__37428\,
            I => \N__37417\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__37425\,
            I => \N__37417\
        );

    \I__6141\ : Span4Mux_v
    port map (
            O => \N__37422\,
            I => \N__37414\
        );

    \I__6140\ : Span4Mux_h
    port map (
            O => \N__37417\,
            I => \N__37411\
        );

    \I__6139\ : Sp12to4
    port map (
            O => \N__37414\,
            I => \N__37408\
        );

    \I__6138\ : Odrv4
    port map (
            O => \N__37411\,
            I => h_6
        );

    \I__6137\ : Odrv12
    port map (
            O => \N__37408\,
            I => h_6
        );

    \I__6136\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37400\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__37400\,
            I => \N__37397\
        );

    \I__6134\ : Span4Mux_v
    port map (
            O => \N__37397\,
            I => \N__37394\
        );

    \I__6133\ : Span4Mux_h
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__6132\ : Span4Mux_h
    port map (
            O => \N__37391\,
            I => \N__37388\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__37388\,
            I => \ALU.status_17_I_39_c_RNOZ0\
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__37385\,
            I => \N__37382\
        );

    \I__6129\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__37379\,
            I => \N__37376\
        );

    \I__6127\ : Odrv12
    port map (
            O => \N__37376\,
            I => \ALU.mult_365_c_RNOZ0Z_0\
        );

    \I__6126\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37370\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__37370\,
            I => \N__37366\
        );

    \I__6124\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37363\
        );

    \I__6123\ : Odrv12
    port map (
            O => \N__37366\,
            I => \ALU.N_572\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__37363\,
            I => \ALU.N_572\
        );

    \I__6121\ : IoInMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37351\
        );

    \I__6119\ : IoInMux
    port map (
            O => \N__37354\,
            I => \N__37348\
        );

    \I__6118\ : IoSpan4Mux
    port map (
            O => \N__37351\,
            I => \N__37345\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__37348\,
            I => \N__37342\
        );

    \I__6116\ : Sp12to4
    port map (
            O => \N__37345\,
            I => \N__37338\
        );

    \I__6115\ : IoSpan4Mux
    port map (
            O => \N__37342\,
            I => \N__37335\
        );

    \I__6114\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37332\
        );

    \I__6113\ : Span12Mux_s7_h
    port map (
            O => \N__37338\,
            I => \N__37329\
        );

    \I__6112\ : Sp12to4
    port map (
            O => \N__37335\,
            I => \N__37326\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__37332\,
            I => \N__37323\
        );

    \I__6110\ : Span12Mux_h
    port map (
            O => \N__37329\,
            I => \N__37318\
        );

    \I__6109\ : Span12Mux_h
    port map (
            O => \N__37326\,
            I => \N__37318\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__37323\,
            I => \N__37315\
        );

    \I__6107\ : Span12Mux_v
    port map (
            O => \N__37318\,
            I => \N__37312\
        );

    \I__6106\ : Span4Mux_v
    port map (
            O => \N__37315\,
            I => \N__37309\
        );

    \I__6105\ : Odrv12
    port map (
            O => \N__37312\,
            I => bus_11
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__37309\,
            I => bus_11
        );

    \I__6103\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37301\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__37301\,
            I => \N__37298\
        );

    \I__6101\ : Odrv4
    port map (
            O => \N__37298\,
            I => \ALU.mult_11\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__37295\,
            I => \ALU.mult_552_c_RNI70R9DAZ0_cascade_\
        );

    \I__6099\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37289\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__37289\,
            I => \ALU.rshift_11\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__37286\,
            I => \N__37282\
        );

    \I__6096\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37277\
        );

    \I__6095\ : InMux
    port map (
            O => \N__37282\,
            I => \N__37277\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__37277\,
            I => \ALU.a_15_am_rn_0_11\
        );

    \I__6093\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37271\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__37271\,
            I => \ALU.mult_552_c_RNI70R9DAZ0\
        );

    \I__6091\ : CascadeMux
    port map (
            O => \N__37268\,
            I => \ALU.mult_552_c_RNIOT7VLFZ0_cascade_\
        );

    \I__6090\ : CascadeMux
    port map (
            O => \N__37265\,
            I => \N__37262\
        );

    \I__6089\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37256\
        );

    \I__6088\ : InMux
    port map (
            O => \N__37261\,
            I => \N__37256\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__37256\,
            I => \N__37253\
        );

    \I__6086\ : Span4Mux_v
    port map (
            O => \N__37253\,
            I => \N__37250\
        );

    \I__6085\ : Span4Mux_h
    port map (
            O => \N__37250\,
            I => \N__37247\
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__37247\,
            I => \ALU.aZ0Z_11\
        );

    \I__6083\ : CascadeMux
    port map (
            O => \N__37244\,
            I => \ALU.a_15_m3_sZ0Z_13_cascade_\
        );

    \I__6082\ : CascadeMux
    port map (
            O => \N__37241\,
            I => \ALU.a32Z0Z_0_cascade_\
        );

    \I__6081\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37235\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37231\
        );

    \I__6079\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37228\
        );

    \I__6078\ : Span4Mux_h
    port map (
            O => \N__37231\,
            I => \N__37225\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__37228\,
            I => \N__37222\
        );

    \I__6076\ : Span4Mux_v
    port map (
            O => \N__37225\,
            I => \N__37217\
        );

    \I__6075\ : Span4Mux_h
    port map (
            O => \N__37222\,
            I => \N__37217\
        );

    \I__6074\ : Span4Mux_h
    port map (
            O => \N__37217\,
            I => \N__37214\
        );

    \I__6073\ : Span4Mux_v
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__6072\ : Odrv4
    port map (
            O => \N__37211\,
            I => \ALU.aZ0Z_1\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__37208\,
            I => \ALU.d_RNICUA7B5Z0Z_0_cascade_\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__37205\,
            I => \N__37202\
        );

    \I__6069\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37199\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__37199\,
            I => \N__37196\
        );

    \I__6067\ : Odrv12
    port map (
            O => \N__37196\,
            I => \ALU.d_RNIL3JT71Z0Z_0\
        );

    \I__6066\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__6064\ : Span4Mux_h
    port map (
            O => \N__37187\,
            I => \N__37184\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__37184\,
            I => \ALU.N_556\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__37181\,
            I => \ALU.N_556_cascade_\
        );

    \I__6061\ : InMux
    port map (
            O => \N__37178\,
            I => \N__37175\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__37175\,
            I => \ALU.d_RNI3MGBH1Z0Z_1\
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__37172\,
            I => \N__37169\
        );

    \I__6058\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37166\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__37166\,
            I => \ALU.mult_25_11\
        );

    \I__6056\ : InMux
    port map (
            O => \N__37163\,
            I => \ALU.mult_29_c10\
        );

    \I__6055\ : InMux
    port map (
            O => \N__37160\,
            I => \ALU.mult_29_c11\
        );

    \I__6054\ : InMux
    port map (
            O => \N__37157\,
            I => \N__37154\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__37154\,
            I => \ALU.mult_25_13\
        );

    \I__6052\ : InMux
    port map (
            O => \N__37151\,
            I => \ALU.mult_29_c12\
        );

    \I__6051\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37145\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__37145\,
            I => \ALU.mult_25_14\
        );

    \I__6049\ : InMux
    port map (
            O => \N__37142\,
            I => \ALU.mult_29_c13\
        );

    \I__6048\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__37136\,
            I => \ALU.mult_516_c_RNI98SKDCZ0\
        );

    \I__6046\ : InMux
    port map (
            O => \N__37133\,
            I => \ALU.mult_29_c14\
        );

    \I__6045\ : InMux
    port map (
            O => \N__37130\,
            I => \N__37127\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__37121\,
            I => \N__37117\
        );

    \I__6041\ : InMux
    port map (
            O => \N__37120\,
            I => \N__37114\
        );

    \I__6040\ : Span4Mux_h
    port map (
            O => \N__37117\,
            I => \N__37107\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__37114\,
            I => \N__37107\
        );

    \I__6038\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37104\
        );

    \I__6037\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37101\
        );

    \I__6036\ : Odrv4
    port map (
            O => \N__37107\,
            I => bus_0_10
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__37104\,
            I => bus_0_10
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__37101\,
            I => bus_0_10
        );

    \I__6033\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__37091\,
            I => \ALU.mult_10\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__37088\,
            I => \ALU.mult_549_c_RNIB6TIDGZ0_cascade_\
        );

    \I__6030\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37082\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__37082\,
            I => \ALU.a_15_am_1_10\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__37079\,
            I => \ALU.mult_549_c_RNIE7260OZ0_cascade_\
        );

    \I__6027\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37072\
        );

    \I__6026\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37069\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__37072\,
            I => \N__37064\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__37069\,
            I => \N__37064\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__6022\ : Span4Mux_v
    port map (
            O => \N__37061\,
            I => \N__37058\
        );

    \I__6021\ : Sp12to4
    port map (
            O => \N__37058\,
            I => \N__37055\
        );

    \I__6020\ : Odrv12
    port map (
            O => \N__37055\,
            I => \ALU.aZ0Z_10\
        );

    \I__6019\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37049\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__37049\,
            I => \N__37046\
        );

    \I__6017\ : Span4Mux_h
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__37043\,
            I => \ALU.mult_365_c_RNOZ0\
        );

    \I__6015\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37037\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__6013\ : Span4Mux_h
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__6012\ : Odrv4
    port map (
            O => \N__37031\,
            I => \ALU.c_RNIF6GEF1Z0Z_12\
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__37028\,
            I => \N__37025\
        );

    \I__6010\ : InMux
    port map (
            O => \N__37025\,
            I => \N__37022\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__37022\,
            I => \N__37019\
        );

    \I__6008\ : Odrv4
    port map (
            O => \N__37019\,
            I => \ALU.c_RNINUT6PZ0Z_13\
        );

    \I__6007\ : InMux
    port map (
            O => \N__37016\,
            I => \ALU.mult_13_c13\
        );

    \I__6006\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__37007\,
            I => \ALU.c_RNIS83N71Z0Z_12\
        );

    \I__6003\ : InMux
    port map (
            O => \N__37004\,
            I => \ALU.mult_13_c14\
        );

    \I__6002\ : CascadeMux
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__6001\ : InMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__5999\ : Span4Mux_h
    port map (
            O => \N__36992\,
            I => \N__36989\
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__36989\,
            I => \ALU.d_RNIL4PC21Z0Z_6\
        );

    \I__5997\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__36983\,
            I => \ALU.mult_5_5\
        );

    \I__5995\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36977\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__5993\ : Span4Mux_h
    port map (
            O => \N__36974\,
            I => \N__36971\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__36971\,
            I => \ALU.mult_9_9\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__36968\,
            I => \N__36965\
        );

    \I__5990\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36962\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__36962\,
            I => \ALU.mult_25_9\
        );

    \I__5988\ : InMux
    port map (
            O => \N__36959\,
            I => \ALU.mult_29_c8\
        );

    \I__5987\ : InMux
    port map (
            O => \N__36956\,
            I => \ALU.mult_29_c9\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__36953\,
            I => \PROM.ROMDATA.m506_cascade_\
        );

    \I__5985\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36944\
        );

    \I__5984\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36944\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__36944\,
            I => \N__36941\
        );

    \I__5982\ : Span4Mux_h
    port map (
            O => \N__36941\,
            I => \N__36938\
        );

    \I__5981\ : Span4Mux_v
    port map (
            O => \N__36938\,
            I => \N__36935\
        );

    \I__5980\ : Odrv4
    port map (
            O => \N__36935\,
            I => \PROM.ROMDATA.N_571_mux\
        );

    \I__5979\ : InMux
    port map (
            O => \N__36932\,
            I => \N__36929\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__36929\,
            I => \N__36926\
        );

    \I__5977\ : Span4Mux_v
    port map (
            O => \N__36926\,
            I => \N__36922\
        );

    \I__5976\ : CascadeMux
    port map (
            O => \N__36925\,
            I => \N__36919\
        );

    \I__5975\ : Span4Mux_h
    port map (
            O => \N__36922\,
            I => \N__36915\
        );

    \I__5974\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36910\
        );

    \I__5973\ : InMux
    port map (
            O => \N__36918\,
            I => \N__36910\
        );

    \I__5972\ : Span4Mux_v
    port map (
            O => \N__36915\,
            I => \N__36905\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__36910\,
            I => \N__36905\
        );

    \I__5970\ : Span4Mux_v
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__36902\,
            I => \N_177\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__36899\,
            I => \ALU.d_RNI64MA6Z0Z_0_cascade_\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__36896\,
            I => \ALU.log_1_3_ns_1_1_0_cascade_\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__36893\,
            I => \ALU.log_1_3_ns_1_0_cascade_\
        );

    \I__5965\ : CascadeMux
    port map (
            O => \N__36890\,
            I => \ALU.log_1_0_cascade_\
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__36887\,
            I => \ALU.status_8_5_0_cascade_\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__36884\,
            I => \N__36880\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__36883\,
            I => \N__36875\
        );

    \I__5961\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36872\
        );

    \I__5960\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36869\
        );

    \I__5959\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36866\
        );

    \I__5958\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36863\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__36872\,
            I => \N__36860\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__36869\,
            I => \N__36857\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__36866\,
            I => \N__36854\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__36863\,
            I => \N__36851\
        );

    \I__5953\ : Span4Mux_h
    port map (
            O => \N__36860\,
            I => \N__36848\
        );

    \I__5952\ : Span4Mux_h
    port map (
            O => \N__36857\,
            I => \N__36841\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__36854\,
            I => \N__36841\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__36851\,
            I => \N__36841\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__36848\,
            I => \CONTROL.N_384_0\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__36841\,
            I => \CONTROL.N_384_0\
        );

    \I__5947\ : CascadeMux
    port map (
            O => \N__36836\,
            I => \CONTROL.N_209_cascade_\
        );

    \I__5946\ : CascadeMux
    port map (
            O => \N__36833\,
            I => \N__36830\
        );

    \I__5945\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36827\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__36827\,
            I => \CONTROL.un1_busState114_1_0_0_0\
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__36824\,
            I => \CONTROL.N_349_cascade_\
        );

    \I__5942\ : InMux
    port map (
            O => \N__36821\,
            I => \N__36818\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__36818\,
            I => \N__36814\
        );

    \I__5940\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36810\
        );

    \I__5939\ : Span4Mux_h
    port map (
            O => \N__36814\,
            I => \N__36807\
        );

    \I__5938\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36804\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__36810\,
            I => \CONTROL.N_246\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__36807\,
            I => \CONTROL.N_246\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__36804\,
            I => \CONTROL.N_246\
        );

    \I__5934\ : InMux
    port map (
            O => \N__36797\,
            I => \N__36794\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__36794\,
            I => \N__36791\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__36791\,
            I => \CONTROL.m38_i_1\
        );

    \I__5931\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36785\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__36785\,
            I => \CONTROL.N_348\
        );

    \I__5929\ : InMux
    port map (
            O => \N__36782\,
            I => \N__36779\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__36779\,
            I => \N__36775\
        );

    \I__5927\ : InMux
    port map (
            O => \N__36778\,
            I => \N__36772\
        );

    \I__5926\ : Span4Mux_h
    port map (
            O => \N__36775\,
            I => \N__36769\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__36772\,
            I => \N__36766\
        );

    \I__5924\ : Span4Mux_h
    port map (
            O => \N__36769\,
            I => \N__36763\
        );

    \I__5923\ : Span4Mux_h
    port map (
            O => \N__36766\,
            I => \N__36760\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__36763\,
            I => \CONTROL.programCounter_1_12\
        );

    \I__5921\ : Odrv4
    port map (
            O => \N__36760\,
            I => \CONTROL.programCounter_1_12\
        );

    \I__5920\ : InMux
    port map (
            O => \N__36755\,
            I => \N__36752\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__36752\,
            I => \CONTROL.programCounter_1_reto_12\
        );

    \I__5918\ : CascadeMux
    port map (
            O => \N__36749\,
            I => \controlWord_1_cascade_\
        );

    \I__5917\ : CascadeMux
    port map (
            O => \N__36746\,
            I => \CONTROL.N_420_cascade_\
        );

    \I__5916\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36740\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__36740\,
            I => \N__36737\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__36737\,
            I => \N__36734\
        );

    \I__5913\ : Sp12to4
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__5912\ : Odrv12
    port map (
            O => \N__36731\,
            I => \CONTROL.programCounter_1_axb_5\
        );

    \I__5911\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__5909\ : Span4Mux_v
    port map (
            O => \N__36722\,
            I => \N__36719\
        );

    \I__5908\ : Sp12to4
    port map (
            O => \N__36719\,
            I => \N__36716\
        );

    \I__5907\ : Odrv12
    port map (
            O => \N__36716\,
            I => \CONTROL.programCounter_1_axb_0\
        );

    \I__5906\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__36710\,
            I => \N__36707\
        );

    \I__5904\ : Span12Mux_h
    port map (
            O => \N__36707\,
            I => \N__36704\
        );

    \I__5903\ : Odrv12
    port map (
            O => \N__36704\,
            I => \CONTROL.N_105_i\
        );

    \I__5902\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36698\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36695\
        );

    \I__5900\ : Odrv12
    port map (
            O => \N__36695\,
            I => \CONTROL.N_427\
        );

    \I__5899\ : CascadeMux
    port map (
            O => \N__36692\,
            I => \PROM_ROMDATA_dintern_5ro_cascade_\
        );

    \I__5898\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36685\
        );

    \I__5897\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36681\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__36685\,
            I => \N__36677\
        );

    \I__5895\ : InMux
    port map (
            O => \N__36684\,
            I => \N__36674\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36671\
        );

    \I__5893\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36668\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__36677\,
            I => \N__36663\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__36674\,
            I => \N__36663\
        );

    \I__5890\ : Span4Mux_v
    port map (
            O => \N__36671\,
            I => \N__36658\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__36668\,
            I => \N__36658\
        );

    \I__5888\ : Span4Mux_h
    port map (
            O => \N__36663\,
            I => \N__36655\
        );

    \I__5887\ : Odrv4
    port map (
            O => \N__36658\,
            I => \CONTROL.N_80_0\
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__36655\,
            I => \CONTROL.N_80_0\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__36650\,
            I => \N__36647\
        );

    \I__5884\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36644\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__36644\,
            I => \N__36641\
        );

    \I__5882\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36638\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__36638\,
            I => \CONTROL.g0_1_i_3Z0Z_1\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__36635\,
            I => \CONTROL.N_48_0_cascade_\
        );

    \I__5879\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36629\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__36629\,
            I => \CONTROL.un1_controlWord_14_i_0\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__36626\,
            I => \N__36622\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__36625\,
            I => \N__36618\
        );

    \I__5875\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36613\
        );

    \I__5874\ : InMux
    port map (
            O => \N__36621\,
            I => \N__36613\
        );

    \I__5873\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36610\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__36613\,
            I => \N__36606\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__36610\,
            I => \N__36602\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__36609\,
            I => \N__36599\
        );

    \I__5869\ : Span4Mux_v
    port map (
            O => \N__36606\,
            I => \N__36596\
        );

    \I__5868\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36593\
        );

    \I__5867\ : Span4Mux_v
    port map (
            O => \N__36602\,
            I => \N__36590\
        );

    \I__5866\ : InMux
    port map (
            O => \N__36599\,
            I => \N__36587\
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__36596\,
            I => \CONTROL.N_87_0\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__36593\,
            I => \CONTROL.N_87_0\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__36590\,
            I => \CONTROL.N_87_0\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__36587\,
            I => \CONTROL.N_87_0\
        );

    \I__5861\ : InMux
    port map (
            O => \N__36578\,
            I => \N__36575\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__36575\,
            I => \N__36572\
        );

    \I__5859\ : Span4Mux_h
    port map (
            O => \N__36572\,
            I => \N__36569\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__36569\,
            I => \CONTROL.un1_busState97_1_0_1_0\
        );

    \I__5857\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36563\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__36560\,
            I => \N__36557\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__36557\,
            I => \CONTROL.dout_reto_7\
        );

    \I__5853\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36551\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__36551\,
            I => \N__36548\
        );

    \I__5851\ : Span4Mux_h
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__36545\,
            I => \N__36542\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__36542\,
            I => \CONTROL.addrstack_reto_7\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__36539\,
            I => \CONTROL.N_422_cascade_\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__36536\,
            I => \progRomAddress_7_cascade_\
        );

    \I__5846\ : CascadeMux
    port map (
            O => \N__36533\,
            I => \CONTROL.N_340_cascade_\
        );

    \I__5845\ : CEMux
    port map (
            O => \N__36530\,
            I => \N__36527\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__36527\,
            I => \N__36524\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__36524\,
            I => \N__36521\
        );

    \I__5842\ : Odrv4
    port map (
            O => \N__36521\,
            I => \CONTROL.un1_busState103_0_0\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__36518\,
            I => \CONTROL.un1_busState114_2_0_0_xZ0Z0_cascade_\
        );

    \I__5840\ : InMux
    port map (
            O => \N__36515\,
            I => \N__36512\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__36512\,
            I => \CONTROL.un1_busState114_2_0_0_xZ0Z1\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__36509\,
            I => \CONTROL.un1_busState114_2_0_0_0_cascade_\
        );

    \I__5837\ : InMux
    port map (
            O => \N__36506\,
            I => \N__36503\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__36503\,
            I => \N__36500\
        );

    \I__5835\ : Span4Mux_h
    port map (
            O => \N__36500\,
            I => \N__36497\
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__36497\,
            I => \CONTROL.aluReadBus_1_sqmuxa_0_a2_2Z0Z_0\
        );

    \I__5833\ : InMux
    port map (
            O => \N__36494\,
            I => \N__36491\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__36491\,
            I => \N__36488\
        );

    \I__5831\ : Span4Mux_h
    port map (
            O => \N__36488\,
            I => \N__36484\
        );

    \I__5830\ : CascadeMux
    port map (
            O => \N__36487\,
            I => \N__36481\
        );

    \I__5829\ : Span4Mux_v
    port map (
            O => \N__36484\,
            I => \N__36478\
        );

    \I__5828\ : InMux
    port map (
            O => \N__36481\,
            I => \N__36475\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__36478\,
            I => \CONTROL.N_83_0\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__36475\,
            I => \CONTROL.N_83_0\
        );

    \I__5825\ : InMux
    port map (
            O => \N__36470\,
            I => \N__36467\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__5823\ : Span4Mux_v
    port map (
            O => \N__36464\,
            I => \N__36461\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__36461\,
            I => \N__36458\
        );

    \I__5821\ : Span4Mux_h
    port map (
            O => \N__36458\,
            I => \N__36455\
        );

    \I__5820\ : Odrv4
    port map (
            O => \N__36455\,
            I => \CONTROL.increment28lto5_1_1_0\
        );

    \I__5819\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36449\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__36449\,
            I => \N__36444\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__36448\,
            I => \N__36440\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__36447\,
            I => \N__36437\
        );

    \I__5815\ : Span4Mux_v
    port map (
            O => \N__36444\,
            I => \N__36434\
        );

    \I__5814\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36426\
        );

    \I__5813\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36426\
        );

    \I__5812\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36426\
        );

    \I__5811\ : Sp12to4
    port map (
            O => \N__36434\,
            I => \N__36423\
        );

    \I__5810\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36420\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__36426\,
            I => \N__36417\
        );

    \I__5808\ : Odrv12
    port map (
            O => \N__36423\,
            I => \CONTROL.N_101_0\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__36420\,
            I => \CONTROL.N_101_0\
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__36417\,
            I => \CONTROL.N_101_0\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__36410\,
            I => \CONTROL.N_320_cascade_\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__36407\,
            I => \CONTROL.un1_busState103_0_0_cascade_\
        );

    \I__5803\ : CascadeMux
    port map (
            O => \N__36404\,
            I => \N__36401\
        );

    \I__5802\ : InMux
    port map (
            O => \N__36401\,
            I => \N__36398\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__36398\,
            I => \N__36394\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__36397\,
            I => \N__36391\
        );

    \I__5799\ : Span4Mux_h
    port map (
            O => \N__36394\,
            I => \N__36388\
        );

    \I__5798\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36385\
        );

    \I__5797\ : Span4Mux_h
    port map (
            O => \N__36388\,
            I => \N__36382\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__36385\,
            I => \CONTROL.N_95_0\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__36382\,
            I => \CONTROL.N_95_0\
        );

    \I__5794\ : InMux
    port map (
            O => \N__36377\,
            I => \N__36374\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__36374\,
            I => \CONTROL.N_318\
        );

    \I__5792\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36365\
        );

    \I__5791\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36365\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__36365\,
            I => \N__36358\
        );

    \I__5789\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36353\
        );

    \I__5788\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36353\
        );

    \I__5787\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36348\
        );

    \I__5786\ : InMux
    port map (
            O => \N__36361\,
            I => \N__36348\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__36358\,
            I => \aluOperand1_fast_2\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__36353\,
            I => \aluOperand1_fast_2\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__36348\,
            I => \aluOperand1_fast_2\
        );

    \I__5782\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36333\
        );

    \I__5781\ : InMux
    port map (
            O => \N__36340\,
            I => \N__36333\
        );

    \I__5780\ : InMux
    port map (
            O => \N__36339\,
            I => \N__36328\
        );

    \I__5779\ : InMux
    port map (
            O => \N__36338\,
            I => \N__36328\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__36333\,
            I => \N__36319\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__36328\,
            I => \N__36319\
        );

    \I__5776\ : InMux
    port map (
            O => \N__36327\,
            I => \N__36310\
        );

    \I__5775\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36310\
        );

    \I__5774\ : InMux
    port map (
            O => \N__36325\,
            I => \N__36305\
        );

    \I__5773\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36305\
        );

    \I__5772\ : Span4Mux_h
    port map (
            O => \N__36319\,
            I => \N__36302\
        );

    \I__5771\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36297\
        );

    \I__5770\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36297\
        );

    \I__5769\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36292\
        );

    \I__5768\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36292\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__36310\,
            I => \aluOperand1_fast_1\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__36305\,
            I => \aluOperand1_fast_1\
        );

    \I__5765\ : Odrv4
    port map (
            O => \N__36302\,
            I => \aluOperand1_fast_1\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__36297\,
            I => \aluOperand1_fast_1\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__36292\,
            I => \aluOperand1_fast_1\
        );

    \I__5762\ : InMux
    port map (
            O => \N__36281\,
            I => \N__36278\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__36278\,
            I => \N__36275\
        );

    \I__5760\ : Span4Mux_h
    port map (
            O => \N__36275\,
            I => \N__36272\
        );

    \I__5759\ : Span4Mux_v
    port map (
            O => \N__36272\,
            I => \N__36269\
        );

    \I__5758\ : Odrv4
    port map (
            O => \N__36269\,
            I => \CONTROL.increment28lto5_1_1_3\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__36266\,
            I => \CONTROL.increment28lto5_1_1_1_cascade_\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__36263\,
            I => \N__36260\
        );

    \I__5755\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36257\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__36257\,
            I => \N__36254\
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__36254\,
            I => \CONTROL.g0_3_i_a7Z0Z_3\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__36251\,
            I => \PROM.ROMDATA.m221cf1_cascade_\
        );

    \I__5751\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36245\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__36245\,
            I => \PROM.ROMDATA.m221cf1\
        );

    \I__5749\ : CEMux
    port map (
            O => \N__36242\,
            I => \N__36237\
        );

    \I__5748\ : CEMux
    port map (
            O => \N__36241\,
            I => \N__36234\
        );

    \I__5747\ : CEMux
    port map (
            O => \N__36240\,
            I => \N__36231\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__36237\,
            I => \N__36228\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__36234\,
            I => \N__36225\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__36231\,
            I => \N__36222\
        );

    \I__5743\ : Span4Mux_v
    port map (
            O => \N__36228\,
            I => \N__36219\
        );

    \I__5742\ : Span4Mux_v
    port map (
            O => \N__36225\,
            I => \N__36216\
        );

    \I__5741\ : Span4Mux_h
    port map (
            O => \N__36222\,
            I => \N__36213\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__36219\,
            I => \CONTROL.un1_busState98_1_0_0_0\
        );

    \I__5739\ : Odrv4
    port map (
            O => \N__36216\,
            I => \CONTROL.un1_busState98_1_0_0_0\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__36213\,
            I => \CONTROL.un1_busState98_1_0_0_0\
        );

    \I__5737\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36200\
        );

    \I__5736\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36200\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__36200\,
            I => \PROM.ROMDATA.m217\
        );

    \I__5734\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36191\
        );

    \I__5733\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36191\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__36191\,
            I => \PROM.ROMDATA.m221cf0\
        );

    \I__5731\ : InMux
    port map (
            O => \N__36188\,
            I => \N__36185\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__36185\,
            I => \N__36181\
        );

    \I__5729\ : InMux
    port map (
            O => \N__36184\,
            I => \N__36178\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__36181\,
            I => \N__36175\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__36178\,
            I => \ALU.dZ0Z_11\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__36175\,
            I => \ALU.dZ0Z_11\
        );

    \I__5725\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36167\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__36167\,
            I => \N__36164\
        );

    \I__5723\ : Span4Mux_v
    port map (
            O => \N__36164\,
            I => \N__36161\
        );

    \I__5722\ : Odrv4
    port map (
            O => \N__36161\,
            I => \ALU.d_RNI6DCTZ0Z_11\
        );

    \I__5721\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36155\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__36155\,
            I => \N__36152\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__36152\,
            I => \N__36149\
        );

    \I__5718\ : Odrv4
    port map (
            O => \N__36149\,
            I => \ALU.N_920\
        );

    \I__5717\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36143\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__36143\,
            I => \ALU.operand2_3_ns_1_15\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__36140\,
            I => \ALU.dout_3_ns_1_15_cascade_\
        );

    \I__5714\ : InMux
    port map (
            O => \N__36137\,
            I => \N__36133\
        );

    \I__5713\ : InMux
    port map (
            O => \N__36136\,
            I => \N__36130\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__36133\,
            I => \N__36127\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__36130\,
            I => \N__36124\
        );

    \I__5710\ : Span4Mux_v
    port map (
            O => \N__36127\,
            I => \N__36121\
        );

    \I__5709\ : Span4Mux_v
    port map (
            O => \N__36124\,
            I => \N__36118\
        );

    \I__5708\ : Span4Mux_h
    port map (
            O => \N__36121\,
            I => \N__36115\
        );

    \I__5707\ : Sp12to4
    port map (
            O => \N__36118\,
            I => \N__36110\
        );

    \I__5706\ : Sp12to4
    port map (
            O => \N__36115\,
            I => \N__36110\
        );

    \I__5705\ : Span12Mux_h
    port map (
            O => \N__36110\,
            I => \N__36107\
        );

    \I__5704\ : Odrv12
    port map (
            O => \N__36107\,
            I => \ALU.cZ0Z_10\
        );

    \I__5703\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36100\
        );

    \I__5702\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36097\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__36100\,
            I => \N__36092\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__36097\,
            I => \N__36092\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__36092\,
            I => \N__36089\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__36089\,
            I => \N__36086\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__36086\,
            I => \ALU.cZ0Z_11\
        );

    \I__5696\ : InMux
    port map (
            O => \N__36083\,
            I => \N__36080\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__36080\,
            I => \N__36077\
        );

    \I__5694\ : Span4Mux_h
    port map (
            O => \N__36077\,
            I => \N__36074\
        );

    \I__5693\ : Span4Mux_v
    port map (
            O => \N__36074\,
            I => \N__36070\
        );

    \I__5692\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36067\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__36070\,
            I => \ALU.dZ0Z_2\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__36067\,
            I => \ALU.dZ0Z_2\
        );

    \I__5689\ : InMux
    port map (
            O => \N__36062\,
            I => \N__36059\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__36056\,
            I => \N__36052\
        );

    \I__5686\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36049\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__36052\,
            I => \N__36046\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__36049\,
            I => \N__36043\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__36046\,
            I => \N__36040\
        );

    \I__5682\ : Odrv12
    port map (
            O => \N__36043\,
            I => \ALU.dZ0Z_6\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__36040\,
            I => \ALU.dZ0Z_6\
        );

    \I__5680\ : InMux
    port map (
            O => \N__36035\,
            I => \N__36031\
        );

    \I__5679\ : CascadeMux
    port map (
            O => \N__36034\,
            I => \N__36028\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__36031\,
            I => \N__36025\
        );

    \I__5677\ : InMux
    port map (
            O => \N__36028\,
            I => \N__36022\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__36025\,
            I => \N__36019\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__36022\,
            I => \N__36016\
        );

    \I__5674\ : Span4Mux_h
    port map (
            O => \N__36019\,
            I => \N__36013\
        );

    \I__5673\ : Odrv12
    port map (
            O => \N__36016\,
            I => \ALU.dZ0Z_10\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__36013\,
            I => \ALU.dZ0Z_10\
        );

    \I__5671\ : CascadeMux
    port map (
            O => \N__36008\,
            I => \N__36005\
        );

    \I__5670\ : InMux
    port map (
            O => \N__36005\,
            I => \N__36000\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__36004\,
            I => \N__35997\
        );

    \I__5668\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35994\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__36000\,
            I => \N__35991\
        );

    \I__5666\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35988\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__35994\,
            I => \N__35985\
        );

    \I__5664\ : Span4Mux_v
    port map (
            O => \N__35991\,
            I => \N__35980\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__35988\,
            I => \N__35980\
        );

    \I__5662\ : Span4Mux_h
    port map (
            O => \N__35985\,
            I => \N__35975\
        );

    \I__5661\ : Span4Mux_v
    port map (
            O => \N__35980\,
            I => \N__35975\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__35975\,
            I => \N__35972\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__35972\,
            I => f_10
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__35969\,
            I => \N__35964\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__35968\,
            I => \N__35961\
        );

    \I__5656\ : InMux
    port map (
            O => \N__35967\,
            I => \N__35958\
        );

    \I__5655\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35953\
        );

    \I__5654\ : InMux
    port map (
            O => \N__35961\,
            I => \N__35953\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__35958\,
            I => \N__35950\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__35953\,
            I => \N__35947\
        );

    \I__5651\ : Sp12to4
    port map (
            O => \N__35950\,
            I => \N__35944\
        );

    \I__5650\ : Span4Mux_h
    port map (
            O => \N__35947\,
            I => \N__35941\
        );

    \I__5649\ : Span12Mux_v
    port map (
            O => \N__35944\,
            I => \N__35938\
        );

    \I__5648\ : Span4Mux_h
    port map (
            O => \N__35941\,
            I => \N__35935\
        );

    \I__5647\ : Odrv12
    port map (
            O => \N__35938\,
            I => f_11
        );

    \I__5646\ : Odrv4
    port map (
            O => \N__35935\,
            I => f_11
        );

    \I__5645\ : CEMux
    port map (
            O => \N__35930\,
            I => \N__35924\
        );

    \I__5644\ : CEMux
    port map (
            O => \N__35929\,
            I => \N__35921\
        );

    \I__5643\ : CEMux
    port map (
            O => \N__35928\,
            I => \N__35918\
        );

    \I__5642\ : CEMux
    port map (
            O => \N__35927\,
            I => \N__35915\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__35924\,
            I => \N__35912\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__35921\,
            I => \N__35909\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__35918\,
            I => \N__35904\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__35915\,
            I => \N__35904\
        );

    \I__5637\ : Span4Mux_v
    port map (
            O => \N__35912\,
            I => \N__35901\
        );

    \I__5636\ : Span4Mux_v
    port map (
            O => \N__35909\,
            I => \N__35898\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__35904\,
            I => \N__35895\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__35901\,
            I => \N__35888\
        );

    \I__5633\ : Span4Mux_v
    port map (
            O => \N__35898\,
            I => \N__35888\
        );

    \I__5632\ : Span4Mux_h
    port map (
            O => \N__35895\,
            I => \N__35888\
        );

    \I__5631\ : Span4Mux_h
    port map (
            O => \N__35888\,
            I => \N__35885\
        );

    \I__5630\ : Sp12to4
    port map (
            O => \N__35885\,
            I => \N__35882\
        );

    \I__5629\ : Span12Mux_v
    port map (
            O => \N__35882\,
            I => \N__35879\
        );

    \I__5628\ : Odrv12
    port map (
            O => \N__35879\,
            I => \CONSTANT_ZERO_NET\
        );

    \I__5627\ : InMux
    port map (
            O => \N__35876\,
            I => \N__35873\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__35873\,
            I => \N__35869\
        );

    \I__5625\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35866\
        );

    \I__5624\ : Span4Mux_v
    port map (
            O => \N__35869\,
            I => \N__35863\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__35866\,
            I => \N__35858\
        );

    \I__5622\ : Span4Mux_h
    port map (
            O => \N__35863\,
            I => \N__35858\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__35858\,
            I => \N__35855\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__35855\,
            I => \ALU.cZ0Z_2\
        );

    \I__5619\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35848\
        );

    \I__5618\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35845\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__35848\,
            I => \N__35842\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__35845\,
            I => \N__35837\
        );

    \I__5615\ : Span12Mux_v
    port map (
            O => \N__35842\,
            I => \N__35837\
        );

    \I__5614\ : Odrv12
    port map (
            O => \N__35837\,
            I => \ALU.cZ0Z_4\
        );

    \I__5613\ : InMux
    port map (
            O => \N__35834\,
            I => \N__35830\
        );

    \I__5612\ : InMux
    port map (
            O => \N__35833\,
            I => \N__35827\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__35830\,
            I => \N__35824\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__35827\,
            I => \N__35821\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__35824\,
            I => \N__35818\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__35821\,
            I => \N__35815\
        );

    \I__5607\ : Span4Mux_h
    port map (
            O => \N__35818\,
            I => \N__35812\
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__35815\,
            I => \ALU.cZ0Z_6\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__35812\,
            I => \ALU.cZ0Z_6\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__35807\,
            I => \N__35804\
        );

    \I__5603\ : InMux
    port map (
            O => \N__35804\,
            I => \N__35801\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__35801\,
            I => \N__35798\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__35798\,
            I => \N__35793\
        );

    \I__5600\ : InMux
    port map (
            O => \N__35797\,
            I => \N__35790\
        );

    \I__5599\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35787\
        );

    \I__5598\ : Span4Mux_h
    port map (
            O => \N__35793\,
            I => \N__35784\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__35790\,
            I => \N__35779\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__35787\,
            I => \N__35779\
        );

    \I__5595\ : Sp12to4
    port map (
            O => \N__35784\,
            I => \N__35776\
        );

    \I__5594\ : Span12Mux_v
    port map (
            O => \N__35779\,
            I => \N__35773\
        );

    \I__5593\ : Odrv12
    port map (
            O => \N__35776\,
            I => g_4
        );

    \I__5592\ : Odrv12
    port map (
            O => \N__35773\,
            I => g_4
        );

    \I__5591\ : InMux
    port map (
            O => \N__35768\,
            I => \N__35765\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__35765\,
            I => \N__35761\
        );

    \I__5589\ : InMux
    port map (
            O => \N__35764\,
            I => \N__35757\
        );

    \I__5588\ : Span4Mux_h
    port map (
            O => \N__35761\,
            I => \N__35754\
        );

    \I__5587\ : InMux
    port map (
            O => \N__35760\,
            I => \N__35751\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__35757\,
            I => \N__35748\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__35754\,
            I => \N__35745\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__35751\,
            I => \N__35742\
        );

    \I__5583\ : Span4Mux_v
    port map (
            O => \N__35748\,
            I => \N__35739\
        );

    \I__5582\ : Span4Mux_h
    port map (
            O => \N__35745\,
            I => \N__35736\
        );

    \I__5581\ : Span12Mux_v
    port map (
            O => \N__35742\,
            I => \N__35731\
        );

    \I__5580\ : Sp12to4
    port map (
            O => \N__35739\,
            I => \N__35731\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__35736\,
            I => \N__35728\
        );

    \I__5578\ : Odrv12
    port map (
            O => \N__35731\,
            I => g_6
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__35728\,
            I => g_6
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__35723\,
            I => \N__35719\
        );

    \I__5575\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35716\
        );

    \I__5574\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35713\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__35716\,
            I => \N__35709\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35706\
        );

    \I__5571\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35703\
        );

    \I__5570\ : Span4Mux_h
    port map (
            O => \N__35709\,
            I => \N__35700\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__35706\,
            I => \N__35695\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__35703\,
            I => \N__35695\
        );

    \I__5567\ : Span4Mux_v
    port map (
            O => \N__35700\,
            I => \N__35692\
        );

    \I__5566\ : Sp12to4
    port map (
            O => \N__35695\,
            I => \N__35689\
        );

    \I__5565\ : Sp12to4
    port map (
            O => \N__35692\,
            I => \N__35686\
        );

    \I__5564\ : Span12Mux_h
    port map (
            O => \N__35689\,
            I => \N__35683\
        );

    \I__5563\ : Odrv12
    port map (
            O => \N__35686\,
            I => g_10
        );

    \I__5562\ : Odrv12
    port map (
            O => \N__35683\,
            I => g_10
        );

    \I__5561\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__35675\,
            I => \N__35672\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__35672\,
            I => \N__35668\
        );

    \I__5558\ : CascadeMux
    port map (
            O => \N__35671\,
            I => \N__35665\
        );

    \I__5557\ : Span4Mux_h
    port map (
            O => \N__35668\,
            I => \N__35661\
        );

    \I__5556\ : InMux
    port map (
            O => \N__35665\,
            I => \N__35658\
        );

    \I__5555\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35655\
        );

    \I__5554\ : Span4Mux_v
    port map (
            O => \N__35661\,
            I => \N__35652\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__35658\,
            I => \N__35647\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__35655\,
            I => \N__35647\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__35652\,
            I => \N__35644\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__35647\,
            I => \N__35641\
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__35644\,
            I => g_11
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__35641\,
            I => g_11
        );

    \I__5547\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35633\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35628\
        );

    \I__5545\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35625\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__35631\,
            I => \N__35622\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__35628\,
            I => \N__35619\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__35625\,
            I => \N__35616\
        );

    \I__5541\ : InMux
    port map (
            O => \N__35622\,
            I => \N__35613\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__35619\,
            I => \N__35610\
        );

    \I__5539\ : Span4Mux_h
    port map (
            O => \N__35616\,
            I => \N__35605\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__35613\,
            I => \N__35605\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__35610\,
            I => \N__35602\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__35605\,
            I => \N__35599\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__35602\,
            I => f_2
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__35599\,
            I => f_2
        );

    \I__5533\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35591\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__35591\,
            I => \ALU.d_RNIUT8OG4Z0Z_0\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__35588\,
            I => \N__35585\
        );

    \I__5530\ : InMux
    port map (
            O => \N__35585\,
            I => \N__35582\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__35582\,
            I => \N__35579\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__35579\,
            I => \ALU.lshift_3_ns_1_14\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__35576\,
            I => \ALU.N_646_cascade_\
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__35573\,
            I => \ALU.lshift_15_ns_1_14_cascade_\
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__35570\,
            I => \N__35567\
        );

    \I__5524\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35563\
        );

    \I__5523\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35560\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__35563\,
            I => \N__35557\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__35560\,
            I => \N__35554\
        );

    \I__5520\ : Span4Mux_h
    port map (
            O => \N__35557\,
            I => \N__35551\
        );

    \I__5519\ : Span4Mux_v
    port map (
            O => \N__35554\,
            I => \N__35547\
        );

    \I__5518\ : Span4Mux_h
    port map (
            O => \N__35551\,
            I => \N__35544\
        );

    \I__5517\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35541\
        );

    \I__5516\ : Span4Mux_v
    port map (
            O => \N__35547\,
            I => \N__35538\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__35544\,
            I => \N__35533\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__35541\,
            I => \N__35533\
        );

    \I__5513\ : Sp12to4
    port map (
            O => \N__35538\,
            I => \N__35530\
        );

    \I__5512\ : Span4Mux_v
    port map (
            O => \N__35533\,
            I => \N__35527\
        );

    \I__5511\ : Span12Mux_h
    port map (
            O => \N__35530\,
            I => \N__35524\
        );

    \I__5510\ : Span4Mux_h
    port map (
            O => \N__35527\,
            I => \N__35521\
        );

    \I__5509\ : Odrv12
    port map (
            O => \N__35524\,
            I => g_2
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__35521\,
            I => g_2
        );

    \I__5507\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35513\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__35513\,
            I => \N__35510\
        );

    \I__5505\ : Span4Mux_h
    port map (
            O => \N__35510\,
            I => \N__35507\
        );

    \I__5504\ : Odrv4
    port map (
            O => \N__35507\,
            I => \ALU.mult_17_8\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__35504\,
            I => \N__35501\
        );

    \I__5502\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35498\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__35498\,
            I => \ALU.mult_19_8\
        );

    \I__5500\ : InMux
    port map (
            O => \N__35495\,
            I => \ALU.mult_25_c7\
        );

    \I__5499\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35489\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__35489\,
            I => \N__35486\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__35486\,
            I => \N__35483\
        );

    \I__5496\ : Odrv4
    port map (
            O => \N__35483\,
            I => \ALU.mult_17_9\
        );

    \I__5495\ : CascadeMux
    port map (
            O => \N__35480\,
            I => \N__35477\
        );

    \I__5494\ : InMux
    port map (
            O => \N__35477\,
            I => \N__35474\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__35474\,
            I => \ALU.mult_19_9\
        );

    \I__5492\ : InMux
    port map (
            O => \N__35471\,
            I => \ALU.mult_25_c8\
        );

    \I__5491\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__35465\,
            I => \ALU.mult_19_10\
        );

    \I__5489\ : CascadeMux
    port map (
            O => \N__35462\,
            I => \N__35459\
        );

    \I__5488\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35456\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__35456\,
            I => \N__35453\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__35453\,
            I => \N__35450\
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__35450\,
            I => \ALU.mult_17_10\
        );

    \I__5484\ : InMux
    port map (
            O => \N__35447\,
            I => \ALU.mult_25_c9\
        );

    \I__5483\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35441\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__35441\,
            I => \N__35438\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__35438\,
            I => \N__35435\
        );

    \I__5480\ : Odrv4
    port map (
            O => \N__35435\,
            I => \ALU.mult_17_11\
        );

    \I__5479\ : CascadeMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__5478\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__35426\,
            I => \ALU.mult_19_11\
        );

    \I__5476\ : InMux
    port map (
            O => \N__35423\,
            I => \ALU.mult_25_c10\
        );

    \I__5475\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35417\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__35417\,
            I => \N__35414\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__35414\,
            I => \N__35411\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__35411\,
            I => \ALU.mult_17_12\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__35408\,
            I => \N__35405\
        );

    \I__5470\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35402\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__35402\,
            I => \ALU.mult_19_12\
        );

    \I__5468\ : InMux
    port map (
            O => \N__35399\,
            I => \bfn_16_10_0_\
        );

    \I__5467\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35393\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__35393\,
            I => \N__35390\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__35390\,
            I => \N__35387\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__35387\,
            I => \ALU.mult_17_13\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__35384\,
            I => \N__35381\
        );

    \I__5462\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35378\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__35378\,
            I => \ALU.mult_19_13\
        );

    \I__5460\ : InMux
    port map (
            O => \N__35375\,
            I => \ALU.mult_25_c12\
        );

    \I__5459\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35369\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__35366\,
            I => \N__35363\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__35363\,
            I => \ALU.mult_17_14\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__35360\,
            I => \N__35357\
        );

    \I__5454\ : InMux
    port map (
            O => \N__35357\,
            I => \N__35354\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__35354\,
            I => \ALU.mult_19_14\
        );

    \I__5452\ : InMux
    port map (
            O => \N__35351\,
            I => \ALU.mult_25_c13\
        );

    \I__5451\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35345\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__35345\,
            I => \N__35342\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__35342\,
            I => \N__35339\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__35339\,
            I => \ALU.mult_424_c_RNIUVTALZ0Z4\
        );

    \I__5447\ : InMux
    port map (
            O => \N__35336\,
            I => \ALU.mult_25_c14\
        );

    \I__5446\ : CascadeMux
    port map (
            O => \N__35333\,
            I => \PROM.ROMDATA.m2_cascade_\
        );

    \I__5445\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35327\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__35327\,
            I => \ALU.mult_7_6\
        );

    \I__5443\ : CascadeMux
    port map (
            O => \N__35324\,
            I => \N__35321\
        );

    \I__5442\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35318\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__35318\,
            I => \N__35315\
        );

    \I__5440\ : Span4Mux_h
    port map (
            O => \N__35315\,
            I => \N__35312\
        );

    \I__5439\ : Span4Mux_h
    port map (
            O => \N__35312\,
            I => \N__35309\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__35309\,
            I => \ALU.status_18_cry_0_c_RNOZ0\
        );

    \I__5437\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35303\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__35303\,
            I => \N__35300\
        );

    \I__5435\ : Odrv4
    port map (
            O => \N__35300\,
            I => \ALU.mult_5_4\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__35297\,
            I => \N__35294\
        );

    \I__5433\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35291\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__35291\,
            I => \N__35288\
        );

    \I__5431\ : Span4Mux_h
    port map (
            O => \N__35288\,
            I => \N__35285\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__35285\,
            I => \ALU.mult_17_4\
        );

    \I__5429\ : InMux
    port map (
            O => \N__35282\,
            I => \N__35279\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__35279\,
            I => \N__35276\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__35276\,
            I => \N__35273\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__35273\,
            I => \N__35270\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__35270\,
            I => \ALU.mult_391_c_RNIEC73TZ0Z4\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__35267\,
            I => \N__35264\
        );

    \I__5423\ : InMux
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35258\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__35258\,
            I => \N__35255\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__35255\,
            I => \ALU.mult_17_5\
        );

    \I__5419\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35249\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__35249\,
            I => \ALU.mult_5\
        );

    \I__5417\ : InMux
    port map (
            O => \N__35246\,
            I => \ALU.mult_25_c4\
        );

    \I__5416\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35240\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__35240\,
            I => \ALU.mult_173_c_RNIO8AOZ0Z16\
        );

    \I__5414\ : CascadeMux
    port map (
            O => \N__35237\,
            I => \N__35233\
        );

    \I__5413\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35230\
        );

    \I__5412\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35227\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__35230\,
            I => \N__35222\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__35227\,
            I => \N__35222\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__35222\,
            I => \N__35219\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__35219\,
            I => \ALU.mult_17_6\
        );

    \I__5407\ : InMux
    port map (
            O => \N__35216\,
            I => \ALU.mult_25_c5\
        );

    \I__5406\ : InMux
    port map (
            O => \N__35213\,
            I => \N__35210\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__35210\,
            I => \ALU.mult_19_7\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__35207\,
            I => \N__35204\
        );

    \I__5403\ : InMux
    port map (
            O => \N__35204\,
            I => \N__35201\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__35201\,
            I => \N__35198\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__35198\,
            I => \N__35195\
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__35195\,
            I => \ALU.mult_17_7\
        );

    \I__5399\ : InMux
    port map (
            O => \N__35192\,
            I => \ALU.mult_25_c6\
        );

    \I__5398\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35186\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__35186\,
            I => \N__35183\
        );

    \I__5396\ : Span4Mux_h
    port map (
            O => \N__35183\,
            I => \N__35179\
        );

    \I__5395\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35176\
        );

    \I__5394\ : Odrv4
    port map (
            O => \N__35179\,
            I => \CONTROL.N_350_1\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__35176\,
            I => \CONTROL.N_350_1\
        );

    \I__5392\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35168\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__35168\,
            I => \N__35165\
        );

    \I__5390\ : Span4Mux_h
    port map (
            O => \N__35165\,
            I => \N__35162\
        );

    \I__5389\ : Span4Mux_v
    port map (
            O => \N__35162\,
            I => \N__35159\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__35159\,
            I => \CONTROL.N_345\
        );

    \I__5387\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35153\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__35153\,
            I => \N__35150\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__35150\,
            I => \N__35147\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__35147\,
            I => \N__35144\
        );

    \I__5383\ : Odrv4
    port map (
            O => \N__35144\,
            I => \CONTROL.N_346\
        );

    \I__5382\ : InMux
    port map (
            O => \N__35141\,
            I => \N__35138\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__35138\,
            I => \N__35135\
        );

    \I__5380\ : Span4Mux_v
    port map (
            O => \N__35135\,
            I => \N__35131\
        );

    \I__5379\ : InMux
    port map (
            O => \N__35134\,
            I => \N__35128\
        );

    \I__5378\ : Span4Mux_h
    port map (
            O => \N__35131\,
            I => \N__35125\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__35128\,
            I => \CONTROL.N_255\
        );

    \I__5376\ : Odrv4
    port map (
            O => \N__35125\,
            I => \CONTROL.N_255\
        );

    \I__5375\ : CascadeMux
    port map (
            O => \N__35120\,
            I => \CONTROL.N_345_cascade_\
        );

    \I__5374\ : IoInMux
    port map (
            O => \N__35117\,
            I => \N__35114\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__35114\,
            I => \N__35109\
        );

    \I__5372\ : IoInMux
    port map (
            O => \N__35113\,
            I => \N__35106\
        );

    \I__5371\ : IoInMux
    port map (
            O => \N__35112\,
            I => \N__35103\
        );

    \I__5370\ : IoSpan4Mux
    port map (
            O => \N__35109\,
            I => \N__35090\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__35106\,
            I => \N__35090\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__35103\,
            I => \N__35090\
        );

    \I__5367\ : IoInMux
    port map (
            O => \N__35102\,
            I => \N__35087\
        );

    \I__5366\ : IoInMux
    port map (
            O => \N__35101\,
            I => \N__35084\
        );

    \I__5365\ : IoInMux
    port map (
            O => \N__35100\,
            I => \N__35081\
        );

    \I__5364\ : IoInMux
    port map (
            O => \N__35099\,
            I => \N__35078\
        );

    \I__5363\ : IoInMux
    port map (
            O => \N__35098\,
            I => \N__35075\
        );

    \I__5362\ : IoInMux
    port map (
            O => \N__35097\,
            I => \N__35072\
        );

    \I__5361\ : IoSpan4Mux
    port map (
            O => \N__35090\,
            I => \N__35056\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__35087\,
            I => \N__35056\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__35084\,
            I => \N__35056\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__35081\,
            I => \N__35056\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__35078\,
            I => \N__35056\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__35075\,
            I => \N__35056\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__35072\,
            I => \N__35056\
        );

    \I__5354\ : IoInMux
    port map (
            O => \N__35071\,
            I => \N__35053\
        );

    \I__5353\ : IoSpan4Mux
    port map (
            O => \N__35056\,
            I => \N__35045\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__35053\,
            I => \N__35045\
        );

    \I__5351\ : IoInMux
    port map (
            O => \N__35052\,
            I => \N__35042\
        );

    \I__5350\ : IoInMux
    port map (
            O => \N__35051\,
            I => \N__35039\
        );

    \I__5349\ : IoInMux
    port map (
            O => \N__35050\,
            I => \N__35036\
        );

    \I__5348\ : IoSpan4Mux
    port map (
            O => \N__35045\,
            I => \N__35027\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__35042\,
            I => \N__35027\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__35039\,
            I => \N__35027\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__35036\,
            I => \N__35027\
        );

    \I__5344\ : IoSpan4Mux
    port map (
            O => \N__35027\,
            I => \N__35022\
        );

    \I__5343\ : IoInMux
    port map (
            O => \N__35026\,
            I => \N__35019\
        );

    \I__5342\ : IoInMux
    port map (
            O => \N__35025\,
            I => \N__35016\
        );

    \I__5341\ : Span4Mux_s0_h
    port map (
            O => \N__35022\,
            I => \N__35013\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__35019\,
            I => \N__35008\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__35016\,
            I => \N__35008\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__35013\,
            I => \N__35002\
        );

    \I__5337\ : IoSpan4Mux
    port map (
            O => \N__35008\,
            I => \N__35002\
        );

    \I__5336\ : IoInMux
    port map (
            O => \N__35007\,
            I => \N__34999\
        );

    \I__5335\ : Span4Mux_s0_h
    port map (
            O => \N__35002\,
            I => \N__34996\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__34999\,
            I => \N__34991\
        );

    \I__5333\ : Sp12to4
    port map (
            O => \N__34996\,
            I => \N__34991\
        );

    \I__5332\ : Span12Mux_s8_h
    port map (
            O => \N__34991\,
            I => \N__34986\
        );

    \I__5331\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34981\
        );

    \I__5330\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34981\
        );

    \I__5329\ : Span12Mux_v
    port map (
            O => \N__34986\,
            I => \N__34978\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__34981\,
            I => \N__34975\
        );

    \I__5327\ : Odrv12
    port map (
            O => \N__34978\,
            I => \ramWrite\
        );

    \I__5326\ : Odrv12
    port map (
            O => \N__34975\,
            I => \ramWrite\
        );

    \I__5325\ : CEMux
    port map (
            O => \N__34970\,
            I => \N__34967\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__34967\,
            I => \N__34961\
        );

    \I__5323\ : CEMux
    port map (
            O => \N__34966\,
            I => \N__34958\
        );

    \I__5322\ : CEMux
    port map (
            O => \N__34965\,
            I => \N__34955\
        );

    \I__5321\ : CEMux
    port map (
            O => \N__34964\,
            I => \N__34951\
        );

    \I__5320\ : Span4Mux_h
    port map (
            O => \N__34961\,
            I => \N__34946\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__34958\,
            I => \N__34946\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__34955\,
            I => \N__34943\
        );

    \I__5317\ : CEMux
    port map (
            O => \N__34954\,
            I => \N__34940\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__34951\,
            I => \N__34937\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__34946\,
            I => \N__34930\
        );

    \I__5314\ : Span4Mux_v
    port map (
            O => \N__34943\,
            I => \N__34930\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__34940\,
            I => \N__34930\
        );

    \I__5312\ : Span4Mux_h
    port map (
            O => \N__34937\,
            I => \N__34927\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__34930\,
            I => \N__34924\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__34927\,
            I => \CONTROL.un1_busState114_1_0Z0Z_0\
        );

    \I__5309\ : Odrv4
    port map (
            O => \N__34924\,
            I => \CONTROL.un1_busState114_1_0Z0Z_0\
        );

    \I__5308\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34916\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__34916\,
            I => \N__34913\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__34913\,
            I => \N__34910\
        );

    \I__5305\ : Span4Mux_h
    port map (
            O => \N__34910\,
            I => \N__34907\
        );

    \I__5304\ : Span4Mux_v
    port map (
            O => \N__34907\,
            I => \N__34903\
        );

    \I__5303\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34900\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__34903\,
            I => \CONTROL.ctrlOut_10\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__34900\,
            I => \CONTROL.ctrlOut_10\
        );

    \I__5300\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34892\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__34892\,
            I => \N__34889\
        );

    \I__5298\ : Odrv4
    port map (
            O => \N__34889\,
            I => \CONTROL.dout_reto_10\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__34886\,
            I => \PROM.ROMDATA.m1_cascade_\
        );

    \I__5296\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34880\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__34880\,
            I => \CONTROL.N_339\
        );

    \I__5294\ : CascadeMux
    port map (
            O => \N__34877\,
            I => \CONTROL.N_219_cascade_\
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__34874\,
            I => \CONTROL.m28_0_120_i_i_a2_0_0_cascade_\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__34871\,
            I => \CONTROL.busState_1_RNO_1Z0Z_1_cascade_\
        );

    \I__5291\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34865\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__34865\,
            I => \N__34862\
        );

    \I__5289\ : Span4Mux_h
    port map (
            O => \N__34862\,
            I => \N__34859\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__34859\,
            I => \CONTROL.busState_1_RNO_0Z0Z_1\
        );

    \I__5287\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34853\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34850\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__34850\,
            I => \CONTROL.g0_3_i_1_1\
        );

    \I__5284\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34844\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__34844\,
            I => \N__34841\
        );

    \I__5282\ : Span4Mux_v
    port map (
            O => \N__34841\,
            I => \N__34838\
        );

    \I__5281\ : Span4Mux_h
    port map (
            O => \N__34838\,
            I => \N__34835\
        );

    \I__5280\ : Sp12to4
    port map (
            O => \N__34835\,
            I => \N__34832\
        );

    \I__5279\ : Odrv12
    port map (
            O => \N__34832\,
            I => \gpuOut_c_2\
        );

    \I__5278\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34826\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__34826\,
            I => \CONTROL.N_163\
        );

    \I__5276\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34820\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__34820\,
            I => \CONTROL.g0_3_i_2_1\
        );

    \I__5274\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34811\
        );

    \I__5273\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34811\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__34811\,
            I => \CONTROL.un1_addrstackptr_c3_0\
        );

    \I__5271\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34802\
        );

    \I__5270\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34802\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__34802\,
            I => \N__34799\
        );

    \I__5268\ : Span4Mux_h
    port map (
            O => \N__34799\,
            I => \N__34796\
        );

    \I__5267\ : Span4Mux_v
    port map (
            O => \N__34796\,
            I => \N__34792\
        );

    \I__5266\ : CascadeMux
    port map (
            O => \N__34795\,
            I => \N__34789\
        );

    \I__5265\ : Span4Mux_v
    port map (
            O => \N__34792\,
            I => \N__34786\
        );

    \I__5264\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34783\
        );

    \I__5263\ : Odrv4
    port map (
            O => \N__34786\,
            I => \CONTROL.addrstack_1_3\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__34783\,
            I => \CONTROL.addrstack_1_3\
        );

    \I__5261\ : InMux
    port map (
            O => \N__34778\,
            I => \N__34775\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__34775\,
            I => \CONTROL.N_5\
        );

    \I__5259\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34765\
        );

    \I__5258\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34762\
        );

    \I__5257\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34757\
        );

    \I__5256\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34757\
        );

    \I__5255\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34754\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34750\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34743\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__34757\,
            I => \N__34743\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34743\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__34753\,
            I => \N__34740\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__34750\,
            I => \N__34736\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__34743\,
            I => \N__34733\
        );

    \I__5247\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34728\
        );

    \I__5246\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34728\
        );

    \I__5245\ : Span4Mux_h
    port map (
            O => \N__34736\,
            I => \N__34725\
        );

    \I__5244\ : Sp12to4
    port map (
            O => \N__34733\,
            I => \N__34722\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__34728\,
            I => \CONTROL.addrstackptrZ0Z_3\
        );

    \I__5242\ : Odrv4
    port map (
            O => \N__34725\,
            I => \CONTROL.addrstackptrZ0Z_3\
        );

    \I__5241\ : Odrv12
    port map (
            O => \N__34722\,
            I => \CONTROL.addrstackptrZ0Z_3\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__34715\,
            I => \CONTROL.N_83_0_cascade_\
        );

    \I__5239\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__34709\,
            I => \CONTROL.m28_0_120_i_i_4\
        );

    \I__5237\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34703\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__34703\,
            I => \CONTROL.N_75_0\
        );

    \I__5235\ : CascadeMux
    port map (
            O => \N__34700\,
            I => \CONTROL.N_75_0_cascade_\
        );

    \I__5234\ : InMux
    port map (
            O => \N__34697\,
            I => \N__34694\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__34694\,
            I => \N__34691\
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__34691\,
            I => \CONTROL.m38_i_2\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__34688\,
            I => \ALU.c_RNIJMOB4_0Z0Z_1_cascade_\
        );

    \I__5230\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34682\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__34682\,
            I => \N__34678\
        );

    \I__5228\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34675\
        );

    \I__5227\ : Sp12to4
    port map (
            O => \N__34678\,
            I => \N__34670\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__34675\,
            I => \N__34670\
        );

    \I__5225\ : Odrv12
    port map (
            O => \N__34670\,
            I => \ALU.d_RNID42JAZ0Z_1\
        );

    \I__5224\ : InMux
    port map (
            O => \N__34667\,
            I => \N__34664\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__34664\,
            I => \ALU.operand2_6_ns_1_1\
        );

    \I__5222\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34658\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__34658\,
            I => \ALU.N_1246\
        );

    \I__5220\ : CascadeMux
    port map (
            O => \N__34655\,
            I => \ALU.operand2_3_ns_1_1_cascade_\
        );

    \I__5219\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34649\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__34649\,
            I => \ALU.N_1198\
        );

    \I__5217\ : InMux
    port map (
            O => \N__34646\,
            I => \N__34640\
        );

    \I__5216\ : InMux
    port map (
            O => \N__34645\,
            I => \N__34640\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__34640\,
            I => \ALU.combOperand2_d_bmZ0Z_1\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__34637\,
            I => \ALU.N_1198_cascade_\
        );

    \I__5213\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34631\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__34631\,
            I => \ALU.c_RNIJMOB4Z0Z_1\
        );

    \I__5211\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34625\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__34625\,
            I => \CONTROL.g0_3_i_a7_2_1\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__34622\,
            I => \CONTROL.N_5_cascade_\
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__34619\,
            I => \N__34616\
        );

    \I__5207\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34613\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__34613\,
            I => \N__34610\
        );

    \I__5205\ : Span4Mux_v
    port map (
            O => \N__34610\,
            I => \N__34607\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__34607\,
            I => \N__34604\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__34604\,
            I => \CONTROL.addrstackptr_8_3\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__34601\,
            I => \ALU.dout_3_ns_1_3_cascade_\
        );

    \I__5201\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34595\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__34595\,
            I => \ALU.N_1136\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__34592\,
            I => \ALU.N_1088_cascade_\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__34589\,
            I => \aluOut_3_cascade_\
        );

    \I__5197\ : InMux
    port map (
            O => \N__34586\,
            I => \N__34583\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__34583\,
            I => \N__34580\
        );

    \I__5195\ : Span4Mux_h
    port map (
            O => \N__34580\,
            I => \N__34577\
        );

    \I__5194\ : Span4Mux_v
    port map (
            O => \N__34577\,
            I => \N__34574\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__34574\,
            I => \busState_1_RNIH16V3_2\
        );

    \I__5192\ : CascadeMux
    port map (
            O => \N__34571\,
            I => \ALU.dout_3_ns_1_13_cascade_\
        );

    \I__5191\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34562\
        );

    \I__5190\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34562\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__34562\,
            I => \N__34553\
        );

    \I__5188\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34548\
        );

    \I__5187\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34548\
        );

    \I__5186\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34543\
        );

    \I__5185\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34543\
        );

    \I__5184\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34537\
        );

    \I__5183\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34537\
        );

    \I__5182\ : Span4Mux_h
    port map (
            O => \N__34553\,
            I => \N__34534\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__34548\,
            I => \N__34531\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__34543\,
            I => \N__34528\
        );

    \I__5179\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34525\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__34537\,
            I => \N__34518\
        );

    \I__5177\ : Span4Mux_v
    port map (
            O => \N__34534\,
            I => \N__34518\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__34531\,
            I => \N__34518\
        );

    \I__5175\ : Odrv4
    port map (
            O => \N__34528\,
            I => \aluOperand1_2_rep2\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__34525\,
            I => \aluOperand1_2_rep2\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__34518\,
            I => \aluOperand1_2_rep2\
        );

    \I__5172\ : CascadeMux
    port map (
            O => \N__34511\,
            I => \ALU.dout_6_ns_1_13_cascade_\
        );

    \I__5171\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34505\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__34505\,
            I => \ALU.N_1098\
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__34502\,
            I => \ALU.N_1146_cascade_\
        );

    \I__5168\ : InMux
    port map (
            O => \N__34499\,
            I => \N__34496\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__34496\,
            I => \N__34493\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__34493\,
            I => \CONTROL.N_190\
        );

    \I__5165\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34487\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__34487\,
            I => \N__34484\
        );

    \I__5163\ : Span4Mux_h
    port map (
            O => \N__34484\,
            I => \N__34478\
        );

    \I__5162\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34475\
        );

    \I__5161\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34472\
        );

    \I__5160\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34469\
        );

    \I__5159\ : Odrv4
    port map (
            O => \N__34478\,
            I => \CONTROL.bus_7_a1_1_8\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__34475\,
            I => \CONTROL.bus_7_a1_1_8\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__34472\,
            I => \CONTROL.bus_7_a1_1_8\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__34469\,
            I => \CONTROL.bus_7_a1_1_8\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__34460\,
            I => \aluOut_13_cascade_\
        );

    \I__5154\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34451\
        );

    \I__5153\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34451\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__34451\,
            I => \N__34448\
        );

    \I__5151\ : Span4Mux_h
    port map (
            O => \N__34448\,
            I => \N__34445\
        );

    \I__5150\ : Odrv4
    port map (
            O => \N__34445\,
            I => \CONTROL.bus_0_13\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__34442\,
            I => \PROM.ROMDATA.m238_am_1_cascade_\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__34439\,
            I => \PROM.ROMDATA.m238_am_cascade_\
        );

    \I__5147\ : CascadeMux
    port map (
            O => \N__34436\,
            I => \PROM.ROMDATA.m244_ns_1_cascade_\
        );

    \I__5146\ : CascadeMux
    port map (
            O => \N__34433\,
            I => \N__34429\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__34432\,
            I => \N__34424\
        );

    \I__5144\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34421\
        );

    \I__5143\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34414\
        );

    \I__5142\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34414\
        );

    \I__5141\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34414\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__34421\,
            I => \PROM.ROMDATA.m244_ns_1\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__34414\,
            I => \PROM.ROMDATA.m244_ns_1\
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__34409\,
            I => \ALU.dout_6_ns_1_3_cascade_\
        );

    \I__5137\ : CascadeMux
    port map (
            O => \N__34406\,
            I => \aluOut_9_cascade_\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__34403\,
            I => \N__34400\
        );

    \I__5135\ : InMux
    port map (
            O => \N__34400\,
            I => \N__34396\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__34399\,
            I => \N__34393\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__34396\,
            I => \N__34389\
        );

    \I__5132\ : InMux
    port map (
            O => \N__34393\,
            I => \N__34386\
        );

    \I__5131\ : InMux
    port map (
            O => \N__34392\,
            I => \N__34383\
        );

    \I__5130\ : Span4Mux_h
    port map (
            O => \N__34389\,
            I => \N__34380\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__34386\,
            I => \N__34377\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__34383\,
            I => \N__34374\
        );

    \I__5127\ : Span4Mux_v
    port map (
            O => \N__34380\,
            I => \N__34371\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__34377\,
            I => \N__34366\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__34374\,
            I => \N__34366\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__34371\,
            I => \N__34363\
        );

    \I__5123\ : Span4Mux_v
    port map (
            O => \N__34366\,
            I => \N__34360\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__34363\,
            I => h_2
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__34360\,
            I => h_2
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__34355\,
            I => \ALU.dout_6_ns_1_2_cascade_\
        );

    \I__5119\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34345\
        );

    \I__5117\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34342\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__34345\,
            I => \N__34337\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34337\
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__34337\,
            I => \ALU.aZ0Z_2\
        );

    \I__5113\ : CascadeMux
    port map (
            O => \N__34334\,
            I => \N__34330\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__34333\,
            I => \N__34327\
        );

    \I__5111\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34324\
        );

    \I__5110\ : InMux
    port map (
            O => \N__34327\,
            I => \N__34321\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__34324\,
            I => \N__34318\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__34321\,
            I => \N__34315\
        );

    \I__5107\ : Odrv12
    port map (
            O => \N__34318\,
            I => \ALU.eZ0Z_2\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__34315\,
            I => \ALU.eZ0Z_2\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__34310\,
            I => \ALU.dout_3_ns_1_2_cascade_\
        );

    \I__5104\ : CascadeMux
    port map (
            O => \N__34307\,
            I => \ALU.N_1087_cascade_\
        );

    \I__5103\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34301\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__34301\,
            I => \ALU.N_1135\
        );

    \I__5101\ : InMux
    port map (
            O => \N__34298\,
            I => \N__34294\
        );

    \I__5100\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34291\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__34294\,
            I => \ALU_N_1086\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__34291\,
            I => \ALU_N_1086\
        );

    \I__5097\ : InMux
    port map (
            O => \N__34286\,
            I => \N__34283\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__34283\,
            I => \CONTROL.operand1_ne_RNIBQE03_0Z0Z_0\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__34280\,
            I => \ALU.addsub_cry_1_c_RNIJP8KZ0Z37_cascade_\
        );

    \I__5094\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34274\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__34274\,
            I => \ALU.addsub_cry_1_c_RNIJP8KZ0Z37\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__34271\,
            I => \ALU.addsub_cry_1_c_RNIICPECZ0Z7_cascade_\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__34268\,
            I => \ALU.dout_3_ns_1_9_cascade_\
        );

    \I__5090\ : CascadeMux
    port map (
            O => \N__34265\,
            I => \ALU.dout_6_ns_1_9_cascade_\
        );

    \I__5089\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34259\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__34259\,
            I => \ALU.N_1094\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__34256\,
            I => \ALU.N_1142_cascade_\
        );

    \I__5086\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34250\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__34250\,
            I => \ALU.mult_388_c_RNIBULDPZ0Z3\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__34247\,
            I => \ALU.mult_388_c_RNIEAAJHZ0Z7_cascade_\
        );

    \I__5083\ : IoInMux
    port map (
            O => \N__34244\,
            I => \N__34238\
        );

    \I__5082\ : IoInMux
    port map (
            O => \N__34243\,
            I => \N__34235\
        );

    \I__5081\ : InMux
    port map (
            O => \N__34242\,
            I => \N__34230\
        );

    \I__5080\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34230\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__34238\,
            I => \N__34227\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__34235\,
            I => \N__34224\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34221\
        );

    \I__5076\ : Span12Mux_s6_h
    port map (
            O => \N__34227\,
            I => \N__34218\
        );

    \I__5075\ : IoSpan4Mux
    port map (
            O => \N__34224\,
            I => \N__34215\
        );

    \I__5074\ : Span4Mux_v
    port map (
            O => \N__34221\,
            I => \N__34212\
        );

    \I__5073\ : Span12Mux_h
    port map (
            O => \N__34218\,
            I => \N__34209\
        );

    \I__5072\ : Span4Mux_s2_h
    port map (
            O => \N__34215\,
            I => \N__34206\
        );

    \I__5071\ : Span4Mux_v
    port map (
            O => \N__34212\,
            I => \N__34203\
        );

    \I__5070\ : Span12Mux_v
    port map (
            O => \N__34209\,
            I => \N__34200\
        );

    \I__5069\ : Sp12to4
    port map (
            O => \N__34206\,
            I => \N__34197\
        );

    \I__5068\ : Span4Mux_h
    port map (
            O => \N__34203\,
            I => \N__34194\
        );

    \I__5067\ : Odrv12
    port map (
            O => \N__34200\,
            I => bus_3
        );

    \I__5066\ : Odrv12
    port map (
            O => \N__34197\,
            I => bus_3
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__34194\,
            I => bus_3
        );

    \I__5064\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34184\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__34184\,
            I => \ALU.mult_388_c_RNIEAAJHZ0Z7\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__34181\,
            I => \ALU.mult_388_c_RNIPGN6QZ0Z7_cascade_\
        );

    \I__5061\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34174\
        );

    \I__5060\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34171\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__34174\,
            I => \N__34168\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__34171\,
            I => \N__34165\
        );

    \I__5057\ : Span4Mux_h
    port map (
            O => \N__34168\,
            I => \N__34160\
        );

    \I__5056\ : Span4Mux_v
    port map (
            O => \N__34165\,
            I => \N__34160\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__34160\,
            I => \ALU.a_15_d_sZ0Z_5\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__34157\,
            I => \N__34154\
        );

    \I__5053\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34151\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34148\
        );

    \I__5051\ : Span4Mux_v
    port map (
            O => \N__34148\,
            I => \N__34145\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__34145\,
            I => \ALU.mult_2\
        );

    \I__5049\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34139\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__34139\,
            I => \N__34136\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__34136\,
            I => \ALU.log_1_2\
        );

    \I__5046\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34129\
        );

    \I__5045\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34126\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__34129\,
            I => \ALU.a_15_d_sZ0Z_3\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__34126\,
            I => \ALU.a_15_d_sZ0Z_3\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__34121\,
            I => \ALU.addsub_cry_1_c_RNI8FKPLZ0Z3_cascade_\
        );

    \I__5041\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34115\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__34115\,
            I => \ALU.mult_5_c_RNI6ET5DZ0Z3\
        );

    \I__5039\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34109\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__34109\,
            I => \N__34106\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__34106\,
            I => \N__34103\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__34103\,
            I => \ALU.mult_3_3\
        );

    \I__5035\ : InMux
    port map (
            O => \N__34100\,
            I => \N__34096\
        );

    \I__5034\ : InMux
    port map (
            O => \N__34099\,
            I => \N__34092\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__34096\,
            I => \N__34089\
        );

    \I__5032\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34086\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34083\
        );

    \I__5030\ : Sp12to4
    port map (
            O => \N__34089\,
            I => \N__34078\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__34086\,
            I => \N__34078\
        );

    \I__5028\ : Span4Mux_h
    port map (
            O => \N__34083\,
            I => \N__34075\
        );

    \I__5027\ : Span12Mux_h
    port map (
            O => \N__34078\,
            I => \N__34072\
        );

    \I__5026\ : Odrv4
    port map (
            O => \N__34075\,
            I => \busState_1_RNIBS0U1_2\
        );

    \I__5025\ : Odrv12
    port map (
            O => \N__34072\,
            I => \busState_1_RNIBS0U1_2\
        );

    \I__5024\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34063\
        );

    \I__5023\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34060\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__34063\,
            I => \N__34055\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__34060\,
            I => \N__34055\
        );

    \I__5020\ : Span4Mux_h
    port map (
            O => \N__34055\,
            I => \N__34052\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__34052\,
            I => \operand1_ne_RNIR8FK7_0\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__34049\,
            I => \ALU.status_19_0_cascade_\
        );

    \I__5017\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34043\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__5015\ : Span4Mux_h
    port map (
            O => \N__34040\,
            I => \N__34037\
        );

    \I__5014\ : Odrv4
    port map (
            O => \N__34037\,
            I => \ALU.mult_95_c_RNOZ0\
        );

    \I__5013\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34031\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34028\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__34028\,
            I => \N__34025\
        );

    \I__5010\ : Odrv4
    port map (
            O => \N__34025\,
            I => \ALU.mult_3\
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__34022\,
            I => \ALU.addsub_cry_2_c_RNIUFTGNZ0Z3_cascade_\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__34019\,
            I => \ALU.mult_486_c_RNIPJD0IZ0Z5_cascade_\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__34016\,
            I => \N__34013\
        );

    \I__5006\ : InMux
    port map (
            O => \N__34013\,
            I => \N__34008\
        );

    \I__5005\ : InMux
    port map (
            O => \N__34012\,
            I => \N__34005\
        );

    \I__5004\ : InMux
    port map (
            O => \N__34011\,
            I => \N__34002\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__33997\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__34005\,
            I => \N__33997\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__34002\,
            I => \N__33994\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__33997\,
            I => \N__33990\
        );

    \I__4999\ : Span12Mux_v
    port map (
            O => \N__33994\,
            I => \N__33987\
        );

    \I__4998\ : InMux
    port map (
            O => \N__33993\,
            I => \N__33984\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__33990\,
            I => \ALU.combOperand2_0_5\
        );

    \I__4996\ : Odrv12
    port map (
            O => \N__33987\,
            I => \ALU.combOperand2_0_5\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__33984\,
            I => \ALU.combOperand2_0_5\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__33977\,
            I => \N__33974\
        );

    \I__4993\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33971\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__33971\,
            I => \N__33968\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__33968\,
            I => \ALU.d_RNICGRJGZ0Z_1\
        );

    \I__4990\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33962\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__33962\,
            I => \ALU.addsub_cry_4_c_RNI2RZ0Z6596\
        );

    \I__4988\ : CascadeMux
    port map (
            O => \N__33959\,
            I => \N__33956\
        );

    \I__4987\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33953\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__33953\,
            I => \N__33950\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__33950\,
            I => \ALU.d_RNIBVMTLZ0Z_5\
        );

    \I__4984\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33944\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__33944\,
            I => \N__33941\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__33941\,
            I => \N__33938\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__33938\,
            I => \ALU.d_RNIVMDLOZ0Z_5\
        );

    \I__4980\ : InMux
    port map (
            O => \N__33935\,
            I => \ALU.mult_19_c8\
        );

    \I__4979\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33929\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__33929\,
            I => \N__33926\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__33926\,
            I => \ALU.mult_7_10\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__33923\,
            I => \N__33920\
        );

    \I__4975\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33917\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__33917\,
            I => \ALU.mult_5_10\
        );

    \I__4973\ : InMux
    port map (
            O => \N__33914\,
            I => \ALU.mult_19_c9\
        );

    \I__4972\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33908\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__33908\,
            I => \N__33905\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__33905\,
            I => \ALU.mult_7_11\
        );

    \I__4969\ : CascadeMux
    port map (
            O => \N__33902\,
            I => \N__33899\
        );

    \I__4968\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33896\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__33896\,
            I => \N__33893\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__33893\,
            I => \ALU.mult_5_11\
        );

    \I__4965\ : InMux
    port map (
            O => \N__33890\,
            I => \ALU.mult_19_c10\
        );

    \I__4964\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33884\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__33884\,
            I => \ALU.mult_5_12\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__33881\,
            I => \N__33878\
        );

    \I__4961\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33875\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__33875\,
            I => \N__33872\
        );

    \I__4959\ : Odrv12
    port map (
            O => \N__33872\,
            I => \ALU.mult_7_12\
        );

    \I__4958\ : InMux
    port map (
            O => \N__33869\,
            I => \ALU.mult_19_c11\
        );

    \I__4957\ : InMux
    port map (
            O => \N__33866\,
            I => \N__33863\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__33863\,
            I => \ALU.mult_5_13\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__33860\,
            I => \N__33857\
        );

    \I__4954\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33854\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__33854\,
            I => \N__33851\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__33851\,
            I => \N__33848\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__33848\,
            I => \ALU.mult_7_13\
        );

    \I__4950\ : InMux
    port map (
            O => \N__33845\,
            I => \ALU.mult_19_c12\
        );

    \I__4949\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33839\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__33839\,
            I => \ALU.mult_5_14\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__33836\,
            I => \N__33833\
        );

    \I__4946\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33830\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__33830\,
            I => \N__33827\
        );

    \I__4944\ : Span4Mux_h
    port map (
            O => \N__33827\,
            I => \N__33824\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__33824\,
            I => \ALU.mult_7_14\
        );

    \I__4942\ : InMux
    port map (
            O => \N__33821\,
            I => \bfn_15_10_0_\
        );

    \I__4941\ : InMux
    port map (
            O => \N__33818\,
            I => \ALU.mult_19_c14\
        );

    \I__4940\ : CascadeMux
    port map (
            O => \N__33815\,
            I => \N__33812\
        );

    \I__4939\ : InMux
    port map (
            O => \N__33812\,
            I => \N__33809\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__33809\,
            I => \ALU.mult_19_c14_THRU_CO\
        );

    \I__4937\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33803\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__33800\,
            I => \ALU.mult_3_2\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__33797\,
            I => \N__33794\
        );

    \I__4933\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33791\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__33791\,
            I => \N__33788\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__4930\ : Sp12to4
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__4929\ : Span12Mux_v
    port map (
            O => \N__33782\,
            I => \N__33779\
        );

    \I__4928\ : Span12Mux_v
    port map (
            O => \N__33779\,
            I => \N__33776\
        );

    \I__4927\ : Odrv12
    port map (
            O => \N__33776\,
            I => \CONTROL.addrstack_1_i\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__33773\,
            I => \N__33770\
        );

    \I__4925\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33767\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__33767\,
            I => \ALU.d_RNII2KJ41Z0Z_4\
        );

    \I__4923\ : IoInMux
    port map (
            O => \N__33764\,
            I => \N__33760\
        );

    \I__4922\ : IoInMux
    port map (
            O => \N__33763\,
            I => \N__33757\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__33760\,
            I => \N__33754\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__33757\,
            I => \N__33751\
        );

    \I__4919\ : Span4Mux_s3_h
    port map (
            O => \N__33754\,
            I => \N__33748\
        );

    \I__4918\ : Span4Mux_s3_h
    port map (
            O => \N__33751\,
            I => \N__33745\
        );

    \I__4917\ : Span4Mux_v
    port map (
            O => \N__33748\,
            I => \N__33741\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__33745\,
            I => \N__33738\
        );

    \I__4915\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33735\
        );

    \I__4914\ : Sp12to4
    port map (
            O => \N__33741\,
            I => \N__33732\
        );

    \I__4913\ : Sp12to4
    port map (
            O => \N__33738\,
            I => \N__33729\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33726\
        );

    \I__4911\ : Span12Mux_h
    port map (
            O => \N__33732\,
            I => \N__33721\
        );

    \I__4910\ : Span12Mux_v
    port map (
            O => \N__33729\,
            I => \N__33721\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__33726\,
            I => \N__33718\
        );

    \I__4908\ : Odrv12
    port map (
            O => \N__33721\,
            I => bus_4
        );

    \I__4907\ : Odrv4
    port map (
            O => \N__33718\,
            I => bus_4
        );

    \I__4906\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33710\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__33710\,
            I => \ALU.mult_173_c_RNOZ0\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__33707\,
            I => \N__33704\
        );

    \I__4903\ : InMux
    port map (
            O => \N__33704\,
            I => \N__33701\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__33701\,
            I => \ALU.mult_5_6\
        );

    \I__4901\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33695\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__33695\,
            I => \N__33692\
        );

    \I__4899\ : Odrv12
    port map (
            O => \N__33692\,
            I => \ALU.mult_7_7\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__33689\,
            I => \N__33686\
        );

    \I__4897\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33683\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__33683\,
            I => \ALU.mult_5_7\
        );

    \I__4895\ : InMux
    port map (
            O => \N__33680\,
            I => \ALU.mult_19_c6\
        );

    \I__4894\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__33674\,
            I => \N__33671\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__33668\,
            I => \ALU.mult_7_8\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__33665\,
            I => \N__33662\
        );

    \I__4889\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33659\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__33659\,
            I => \ALU.mult_5_8\
        );

    \I__4887\ : InMux
    port map (
            O => \N__33656\,
            I => \ALU.mult_19_c7\
        );

    \I__4886\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33650\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33647\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__33647\,
            I => \ALU.mult_7_9\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__33644\,
            I => \N__33641\
        );

    \I__4882\ : InMux
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__33638\,
            I => \ALU.mult_5_9\
        );

    \I__4880\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33632\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__33626\,
            I => \N__33623\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__33623\,
            I => \CONTROL.tempCounterZ0Z_0\
        );

    \I__4875\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33617\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__33617\,
            I => \N__33614\
        );

    \I__4873\ : Sp12to4
    port map (
            O => \N__33614\,
            I => \N__33611\
        );

    \I__4872\ : Span12Mux_h
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__4871\ : Odrv12
    port map (
            O => \N__33608\,
            I => \CONTROL.tempCounterZ0Z_5\
        );

    \I__4870\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33602\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__33602\,
            I => \N__33599\
        );

    \I__4868\ : Span4Mux_h
    port map (
            O => \N__33599\,
            I => \N__33596\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__33596\,
            I => \N__33593\
        );

    \I__4866\ : Sp12to4
    port map (
            O => \N__33593\,
            I => \N__33590\
        );

    \I__4865\ : Odrv12
    port map (
            O => \N__33590\,
            I => \CONTROL.tempCounterZ0Z_3\
        );

    \I__4864\ : InMux
    port map (
            O => \N__33587\,
            I => \N__33583\
        );

    \I__4863\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33580\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__33583\,
            I => \N__33577\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33572\
        );

    \I__4860\ : Span4Mux_h
    port map (
            O => \N__33577\,
            I => \N__33572\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__33572\,
            I => \CONTROL.programCounter_1_8\
        );

    \I__4858\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33566\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__33566\,
            I => \N__33563\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__33563\,
            I => \N__33560\
        );

    \I__4855\ : Span4Mux_h
    port map (
            O => \N__33560\,
            I => \N__33557\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__33557\,
            I => \CONTROL.tempCounterZ0Z_8\
        );

    \I__4853\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33551\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__33551\,
            I => \N__33548\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__33548\,
            I => \N__33545\
        );

    \I__4850\ : Span4Mux_h
    port map (
            O => \N__33545\,
            I => \N__33542\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__33542\,
            I => \CONTROL.tempCounterZ0Z_4\
        );

    \I__4848\ : InMux
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__33536\,
            I => \N__33533\
        );

    \I__4846\ : Span4Mux_h
    port map (
            O => \N__33533\,
            I => \N__33530\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__33530\,
            I => \N__33527\
        );

    \I__4844\ : Odrv4
    port map (
            O => \N__33527\,
            I => \CONTROL.tempCounterZ0Z_1\
        );

    \I__4843\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33521\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__33521\,
            I => \N__33518\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__33518\,
            I => \N__33515\
        );

    \I__4840\ : Span4Mux_h
    port map (
            O => \N__33515\,
            I => \N__33512\
        );

    \I__4839\ : Odrv4
    port map (
            O => \N__33512\,
            I => \CONTROL.tempCounterZ0Z_7\
        );

    \I__4838\ : InMux
    port map (
            O => \N__33509\,
            I => \N__33506\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__33506\,
            I => \N__33503\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__33503\,
            I => \N__33500\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__33500\,
            I => \CONTROL.tempCounterZ0Z_12\
        );

    \I__4834\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33494\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__33494\,
            I => \N__33491\
        );

    \I__4832\ : Span4Mux_v
    port map (
            O => \N__33491\,
            I => \N__33488\
        );

    \I__4831\ : Span4Mux_h
    port map (
            O => \N__33488\,
            I => \N__33485\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__33485\,
            I => \CONTROL.tempCounterZ0Z_2\
        );

    \I__4829\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33479\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__33479\,
            I => \N__33476\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__33476\,
            I => \CONTROL.N_430\
        );

    \I__4826\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33470\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__33470\,
            I => \N__33467\
        );

    \I__4824\ : Span4Mux_h
    port map (
            O => \N__33467\,
            I => \N__33464\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__33464\,
            I => \CONTROL.un1_busState98_1_1_0Z0Z_0\
        );

    \I__4822\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33458\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__33458\,
            I => \N__33454\
        );

    \I__4820\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33451\
        );

    \I__4819\ : Span4Mux_h
    port map (
            O => \N__33454\,
            I => \N__33448\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__33451\,
            I => \N__33445\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__33448\,
            I => \CONTROL.programCounter_1_15\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__33445\,
            I => \CONTROL.programCounter_1_15\
        );

    \I__4815\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33437\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__33437\,
            I => \CONTROL.programCounter_1_reto_15\
        );

    \I__4813\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33430\
        );

    \I__4812\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33427\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__33430\,
            I => \CONTROL.ctrlOut_15\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__33427\,
            I => \CONTROL.ctrlOut_15\
        );

    \I__4809\ : InMux
    port map (
            O => \N__33422\,
            I => \N__33419\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__33419\,
            I => \CONTROL.dout_reto_15\
        );

    \I__4807\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33413\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__33413\,
            I => \N__33410\
        );

    \I__4805\ : Span4Mux_v
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__4804\ : Span4Mux_h
    port map (
            O => \N__33407\,
            I => \N__33404\
        );

    \I__4803\ : Odrv4
    port map (
            O => \N__33404\,
            I => \PROM.ROMDATA.m465_am\
        );

    \I__4802\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33398\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__33398\,
            I => \N__33395\
        );

    \I__4800\ : Span4Mux_h
    port map (
            O => \N__33395\,
            I => \N__33392\
        );

    \I__4799\ : Span4Mux_v
    port map (
            O => \N__33392\,
            I => \N__33388\
        );

    \I__4798\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33385\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__33388\,
            I => \CONTROL.ctrlOut_7\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__33385\,
            I => \CONTROL.ctrlOut_7\
        );

    \I__4795\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33377\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__33377\,
            I => \CONTROL.N_180\
        );

    \I__4793\ : InMux
    port map (
            O => \N__33374\,
            I => \N__33371\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__33371\,
            I => \N__33368\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__33368\,
            I => \N__33365\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__33365\,
            I => \N__33362\
        );

    \I__4789\ : Span4Mux_v
    port map (
            O => \N__33362\,
            I => \N__33359\
        );

    \I__4788\ : Span4Mux_h
    port map (
            O => \N__33359\,
            I => \N__33356\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__33356\,
            I => \gpuOut_c_3\
        );

    \I__4786\ : CascadeMux
    port map (
            O => \N__33353\,
            I => \N__33350\
        );

    \I__4785\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33347\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__33347\,
            I => \N_164\
        );

    \I__4783\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33338\
        );

    \I__4782\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33338\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__33338\,
            I => \N__33335\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__33335\,
            I => \N__33332\
        );

    \I__4779\ : Span4Mux_v
    port map (
            O => \N__33332\,
            I => \N__33329\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__33329\,
            I => \N__33326\
        );

    \I__4777\ : IoSpan4Mux
    port map (
            O => \N__33326\,
            I => \N__33323\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__33323\,
            I => \D3_in_c\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__33320\,
            I => \N_164_cascade_\
        );

    \I__4774\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33314\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__33314\,
            I => \N__33310\
        );

    \I__4772\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33307\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__33310\,
            I => \N__33301\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__33307\,
            I => \N__33301\
        );

    \I__4769\ : InMux
    port map (
            O => \N__33306\,
            I => \N__33298\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__33301\,
            I => \controlWord_16\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__33298\,
            I => \controlWord_16\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__33293\,
            I => \N__33290\
        );

    \I__4765\ : CascadeBuf
    port map (
            O => \N__33290\,
            I => \N__33287\
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__33287\,
            I => \N__33284\
        );

    \I__4763\ : CascadeBuf
    port map (
            O => \N__33284\,
            I => \N__33281\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__33281\,
            I => \N__33278\
        );

    \I__4761\ : CascadeBuf
    port map (
            O => \N__33278\,
            I => \N__33275\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__4759\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__33269\,
            I => \N__33266\
        );

    \I__4757\ : Span4Mux_h
    port map (
            O => \N__33266\,
            I => \N__33263\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__33263\,
            I => \N__33260\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__33260\,
            I => \CONTROL_romAddReg_7_0\
        );

    \I__4754\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33254\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33251\
        );

    \I__4752\ : Span4Mux_h
    port map (
            O => \N__33251\,
            I => \N__33248\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__33248\,
            I => \N__33244\
        );

    \I__4750\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33241\
        );

    \I__4749\ : Odrv4
    port map (
            O => \N__33244\,
            I => \controlWord_17\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__33241\,
            I => \controlWord_17\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__33236\,
            I => \controlWord_17_cascade_\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__33233\,
            I => \N__33230\
        );

    \I__4745\ : CascadeBuf
    port map (
            O => \N__33230\,
            I => \N__33227\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__33227\,
            I => \N__33224\
        );

    \I__4743\ : CascadeBuf
    port map (
            O => \N__33224\,
            I => \N__33221\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__33221\,
            I => \N__33218\
        );

    \I__4741\ : CascadeBuf
    port map (
            O => \N__33218\,
            I => \N__33215\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__33215\,
            I => \N__33212\
        );

    \I__4739\ : InMux
    port map (
            O => \N__33212\,
            I => \N__33209\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__4737\ : Span12Mux_s10_v
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__4736\ : Odrv12
    port map (
            O => \N__33203\,
            I => \CONTROL_romAddReg_7_1\
        );

    \I__4735\ : InMux
    port map (
            O => \N__33200\,
            I => \N__33197\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__33197\,
            I => \N__33194\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__33194\,
            I => \CONTROL.N_169\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__33191\,
            I => \N__33188\
        );

    \I__4731\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33185\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__33185\,
            I => \N__33182\
        );

    \I__4729\ : Span4Mux_v
    port map (
            O => \N__33182\,
            I => \N__33179\
        );

    \I__4728\ : Span4Mux_v
    port map (
            O => \N__33179\,
            I => \N__33176\
        );

    \I__4727\ : Sp12to4
    port map (
            O => \N__33176\,
            I => \N__33173\
        );

    \I__4726\ : Span12Mux_h
    port map (
            O => \N__33173\,
            I => \N__33170\
        );

    \I__4725\ : Odrv12
    port map (
            O => \N__33170\,
            I => \D8_in_c\
        );

    \I__4724\ : InMux
    port map (
            O => \N__33167\,
            I => \N__33163\
        );

    \I__4723\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33160\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__33163\,
            I => \N__33157\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__33160\,
            I => \N__33154\
        );

    \I__4720\ : Span4Mux_v
    port map (
            O => \N__33157\,
            I => \N__33151\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__33154\,
            I => \N__33148\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__33151\,
            I => \CONTROL.N_185\
        );

    \I__4717\ : Odrv4
    port map (
            O => \N__33148\,
            I => \CONTROL.N_185\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__33143\,
            I => \N__33140\
        );

    \I__4715\ : InMux
    port map (
            O => \N__33140\,
            I => \N__33136\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__33139\,
            I => \N__33133\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__33136\,
            I => \N__33130\
        );

    \I__4712\ : InMux
    port map (
            O => \N__33133\,
            I => \N__33127\
        );

    \I__4711\ : Span4Mux_v
    port map (
            O => \N__33130\,
            I => \N__33124\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__33127\,
            I => \N__33121\
        );

    \I__4709\ : Span4Mux_v
    port map (
            O => \N__33124\,
            I => \N__33116\
        );

    \I__4708\ : Span4Mux_v
    port map (
            O => \N__33121\,
            I => \N__33116\
        );

    \I__4707\ : Span4Mux_h
    port map (
            O => \N__33116\,
            I => \N__33113\
        );

    \I__4706\ : Span4Mux_h
    port map (
            O => \N__33113\,
            I => \N__33110\
        );

    \I__4705\ : Sp12to4
    port map (
            O => \N__33110\,
            I => \N__33107\
        );

    \I__4704\ : Span12Mux_v
    port map (
            O => \N__33107\,
            I => \N__33104\
        );

    \I__4703\ : Odrv12
    port map (
            O => \N__33104\,
            I => \D4_in_c\
        );

    \I__4702\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33098\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__33098\,
            I => \N__33095\
        );

    \I__4700\ : Span12Mux_h
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__4699\ : Span12Mux_v
    port map (
            O => \N__33092\,
            I => \N__33089\
        );

    \I__4698\ : Odrv12
    port map (
            O => \N__33089\,
            I => \CONTROL.busState_1_RNIU83C1_0Z0Z_2\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__33086\,
            I => \N__33083\
        );

    \I__4696\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33080\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__33080\,
            I => \N__33077\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__33077\,
            I => \N__33074\
        );

    \I__4693\ : Sp12to4
    port map (
            O => \N__33074\,
            I => \N__33071\
        );

    \I__4692\ : Span12Mux_h
    port map (
            O => \N__33071\,
            I => \N__33068\
        );

    \I__4691\ : Odrv12
    port map (
            O => \N__33068\,
            I => \D2_in_c\
        );

    \I__4690\ : InMux
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__33059\
        );

    \I__4688\ : Span4Mux_v
    port map (
            O => \N__33059\,
            I => \N__33054\
        );

    \I__4687\ : InMux
    port map (
            O => \N__33058\,
            I => \N__33051\
        );

    \I__4686\ : CascadeMux
    port map (
            O => \N__33057\,
            I => \N__33048\
        );

    \I__4685\ : Span4Mux_v
    port map (
            O => \N__33054\,
            I => \N__33043\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33043\
        );

    \I__4683\ : InMux
    port map (
            O => \N__33048\,
            I => \N__33040\
        );

    \I__4682\ : Span4Mux_h
    port map (
            O => \N__33043\,
            I => \N__33037\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__33040\,
            I => \N_228_0\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__33037\,
            I => \N_228_0\
        );

    \I__4679\ : InMux
    port map (
            O => \N__33032\,
            I => \N__33029\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__33029\,
            I => \N__33026\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__33026\,
            I => \N__33023\
        );

    \I__4676\ : Sp12to4
    port map (
            O => \N__33023\,
            I => \N__33020\
        );

    \I__4675\ : Odrv12
    port map (
            O => \N__33020\,
            I => \CONTROL.busState_1_RNILAEH1Z0Z_2\
        );

    \I__4674\ : InMux
    port map (
            O => \N__33017\,
            I => \N__33014\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__33014\,
            I => \N__33011\
        );

    \I__4672\ : Span4Mux_v
    port map (
            O => \N__33011\,
            I => \N__33008\
        );

    \I__4671\ : Span4Mux_v
    port map (
            O => \N__33008\,
            I => \N__33005\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__33005\,
            I => \N__33002\
        );

    \I__4669\ : Span4Mux_h
    port map (
            O => \N__33002\,
            I => \N__32999\
        );

    \I__4668\ : IoSpan4Mux
    port map (
            O => \N__32999\,
            I => \N__32996\
        );

    \I__4667\ : Odrv4
    port map (
            O => \N__32996\,
            I => \gpuOut_c_1\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__32993\,
            I => \N__32990\
        );

    \I__4665\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32987\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__32987\,
            I => \N_162\
        );

    \I__4663\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32978\
        );

    \I__4662\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32978\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32975\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__32975\,
            I => \N__32972\
        );

    \I__4659\ : Span4Mux_h
    port map (
            O => \N__32972\,
            I => \N__32969\
        );

    \I__4658\ : Sp12to4
    port map (
            O => \N__32969\,
            I => \N__32966\
        );

    \I__4657\ : Odrv12
    port map (
            O => \N__32966\,
            I => \D1_in_c\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__32963\,
            I => \N_162_cascade_\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__32960\,
            I => \ALU.operand2_3_ns_1_2_cascade_\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__32957\,
            I => \ALU.N_1199_cascade_\
        );

    \I__4653\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32951\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__32951\,
            I => \ALU.N_1199\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__32948\,
            I => \ALU.c_RNIJ1JO4_0Z0Z_2_cascade_\
        );

    \I__4650\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32942\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__32942\,
            I => \ALU.c_RNIJ1JO4Z0Z_2\
        );

    \I__4648\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32930\
        );

    \I__4647\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32930\
        );

    \I__4646\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32930\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__32930\,
            I => \N__32927\
        );

    \I__4644\ : Odrv12
    port map (
            O => \N__32927\,
            I => \ALU.d_RNIARKGBZ0Z_2\
        );

    \I__4643\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32921\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__32921\,
            I => \ALU.operand2_6_ns_1_2\
        );

    \I__4641\ : InMux
    port map (
            O => \N__32918\,
            I => \N__32915\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__32915\,
            I => \ALU.N_1247\
        );

    \I__4639\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32906\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__32906\,
            I => \N__32903\
        );

    \I__4636\ : Span4Mux_v
    port map (
            O => \N__32903\,
            I => \N__32900\
        );

    \I__4635\ : Sp12to4
    port map (
            O => \N__32900\,
            I => \N__32897\
        );

    \I__4634\ : Span12Mux_h
    port map (
            O => \N__32897\,
            I => \N__32894\
        );

    \I__4633\ : Odrv12
    port map (
            O => \N__32894\,
            I => \gpuOut_c_13\
        );

    \I__4632\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32888\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__4630\ : Span4Mux_h
    port map (
            O => \N__32885\,
            I => \N__32882\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__32882\,
            I => \N__32879\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__32879\,
            I => \N__32876\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__32876\,
            I => \N__32873\
        );

    \I__4626\ : Span4Mux_h
    port map (
            O => \N__32873\,
            I => \N__32870\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__32870\,
            I => \D13_in_c\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__32867\,
            I => \CONTROL.N_174_cascade_\
        );

    \I__4623\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32861\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__32861\,
            I => \N__32858\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__32858\,
            I => \N__32855\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__32855\,
            I => \N__32852\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__32852\,
            I => \ALU.d_RNIHD7AOZ0Z_7\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__32849\,
            I => \CONTROL.operand1_ne_RNIHKCU2Z0Z_0_cascade_\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__32846\,
            I => \N__32842\
        );

    \I__4616\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32837\
        );

    \I__4615\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32837\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32834\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__32834\,
            I => \operand1_ne_RNIDN8E7_0\
        );

    \I__4612\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32828\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__32828\,
            I => \ALU.dout_6_ns_1_0\
        );

    \I__4610\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32816\
        );

    \I__4609\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32816\
        );

    \I__4608\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32811\
        );

    \I__4607\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32811\
        );

    \I__4606\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32806\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32801\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__32811\,
            I => \N__32801\
        );

    \I__4603\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32796\
        );

    \I__4602\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32796\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__32806\,
            I => \aluOperand1_2_rep1\
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__32801\,
            I => \aluOperand1_2_rep1\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__32796\,
            I => \aluOperand1_2_rep1\
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__32789\,
            I => \ALU.dout_3_ns_1_0_cascade_\
        );

    \I__4597\ : CascadeMux
    port map (
            O => \N__32786\,
            I => \ALU_N_1085_cascade_\
        );

    \I__4596\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32780\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__32780\,
            I => \CONTROL.operand1_ne_RNIHKCU2_0Z0Z_0\
        );

    \I__4594\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32771\
        );

    \I__4593\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32771\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__32771\,
            I => \ALU_N_1133\
        );

    \I__4591\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32762\
        );

    \I__4590\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32762\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__32762\,
            I => \ALU_N_1085\
        );

    \I__4588\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32753\
        );

    \I__4587\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32753\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__32750\,
            I => \busState_1_RNI9P5V3_2\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__32747\,
            I => \ALU.dout_3_ns_1_1_cascade_\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__32744\,
            I => \ALU_N_1086_cascade_\
        );

    \I__4582\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__32738\,
            I => \ALU_N_1134\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__32735\,
            I => \ALU.dout_6_ns_1_6_cascade_\
        );

    \I__4579\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__32729\,
            I => \N__32725\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__32728\,
            I => \N__32722\
        );

    \I__4576\ : Span4Mux_h
    port map (
            O => \N__32725\,
            I => \N__32719\
        );

    \I__4575\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32716\
        );

    \I__4574\ : Sp12to4
    port map (
            O => \N__32719\,
            I => \N__32713\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__32716\,
            I => \ALU.eZ0Z_6\
        );

    \I__4572\ : Odrv12
    port map (
            O => \N__32713\,
            I => \ALU.eZ0Z_6\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__32708\,
            I => \ALU.dout_3_ns_1_6_cascade_\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__32705\,
            I => \ALU.N_1091_cascade_\
        );

    \I__4569\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32699\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__32699\,
            I => \ALU.N_1139\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__32696\,
            I => \aluOut_6_cascade_\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__4565\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32684\
        );

    \I__4564\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32684\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__32681\,
            I => \N__32678\
        );

    \I__4561\ : Odrv4
    port map (
            O => \N__32678\,
            I => \ALU.d_RNIR3N75Z0Z_6\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__32675\,
            I => \ALU.dout_6_ns_1_1_cascade_\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__32672\,
            I => \ALU_N_1134_cascade_\
        );

    \I__4558\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32666\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__32666\,
            I => \CONTROL.operand1_ne_RNIBQE03Z0Z_0\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__32663\,
            I => \N__32659\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__32662\,
            I => \N__32656\
        );

    \I__4554\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32653\
        );

    \I__4553\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32650\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32645\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__32650\,
            I => \N__32645\
        );

    \I__4550\ : Span4Mux_v
    port map (
            O => \N__32645\,
            I => \N__32642\
        );

    \I__4549\ : Span4Mux_h
    port map (
            O => \N__32642\,
            I => \N__32639\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__32639\,
            I => \ALU.eZ0Z_4\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__32636\,
            I => \N__32632\
        );

    \I__4546\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32629\
        );

    \I__4545\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32626\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__32629\,
            I => \N__32623\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32620\
        );

    \I__4542\ : Span4Mux_v
    port map (
            O => \N__32623\,
            I => \N__32617\
        );

    \I__4541\ : Span4Mux_v
    port map (
            O => \N__32620\,
            I => \N__32614\
        );

    \I__4540\ : Sp12to4
    port map (
            O => \N__32617\,
            I => \N__32609\
        );

    \I__4539\ : Sp12to4
    port map (
            O => \N__32614\,
            I => \N__32609\
        );

    \I__4538\ : Odrv12
    port map (
            O => \N__32609\,
            I => \ALU.eZ0Z_10\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__32606\,
            I => \N__32603\
        );

    \I__4536\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32600\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__32600\,
            I => \N__32596\
        );

    \I__4534\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32593\
        );

    \I__4533\ : Span4Mux_v
    port map (
            O => \N__32596\,
            I => \N__32590\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__32593\,
            I => \N__32587\
        );

    \I__4531\ : Span4Mux_h
    port map (
            O => \N__32590\,
            I => \N__32584\
        );

    \I__4530\ : Span12Mux_v
    port map (
            O => \N__32587\,
            I => \N__32581\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__32584\,
            I => \N__32578\
        );

    \I__4528\ : Odrv12
    port map (
            O => \N__32581\,
            I => \ALU.eZ0Z_11\
        );

    \I__4527\ : Odrv4
    port map (
            O => \N__32578\,
            I => \ALU.eZ0Z_11\
        );

    \I__4526\ : IoInMux
    port map (
            O => \N__32573\,
            I => \N__32570\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32564\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__32569\,
            I => \N__32559\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__32568\,
            I => \N__32555\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__32567\,
            I => \N__32551\
        );

    \I__4521\ : IoSpan4Mux
    port map (
            O => \N__32564\,
            I => \N__32548\
        );

    \I__4520\ : SRMux
    port map (
            O => \N__32563\,
            I => \N__32545\
        );

    \I__4519\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32531\
        );

    \I__4518\ : InMux
    port map (
            O => \N__32559\,
            I => \N__32531\
        );

    \I__4517\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32531\
        );

    \I__4516\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32531\
        );

    \I__4515\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32531\
        );

    \I__4514\ : InMux
    port map (
            O => \N__32551\,
            I => \N__32531\
        );

    \I__4513\ : Span4Mux_s3_v
    port map (
            O => \N__32548\,
            I => \N__32527\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32524\
        );

    \I__4511\ : SRMux
    port map (
            O => \N__32544\,
            I => \N__32521\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__32531\,
            I => \N__32518\
        );

    \I__4509\ : SRMux
    port map (
            O => \N__32530\,
            I => \N__32515\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__32527\,
            I => \N__32502\
        );

    \I__4507\ : Span4Mux_v
    port map (
            O => \N__32524\,
            I => \N__32502\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__32521\,
            I => \N__32502\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__32518\,
            I => \N__32502\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N__32502\
        );

    \I__4503\ : SRMux
    port map (
            O => \N__32514\,
            I => \N__32499\
        );

    \I__4502\ : SRMux
    port map (
            O => \N__32513\,
            I => \N__32496\
        );

    \I__4501\ : Span4Mux_v
    port map (
            O => \N__32502\,
            I => \N__32486\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__32499\,
            I => \N__32486\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__32496\,
            I => \N__32486\
        );

    \I__4498\ : SRMux
    port map (
            O => \N__32495\,
            I => \N__32483\
        );

    \I__4497\ : IoInMux
    port map (
            O => \N__32494\,
            I => \N__32476\
        );

    \I__4496\ : IoInMux
    port map (
            O => \N__32493\,
            I => \N__32473\
        );

    \I__4495\ : Span4Mux_v
    port map (
            O => \N__32486\,
            I => \N__32468\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__32483\,
            I => \N__32468\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__32482\,
            I => \N__32465\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__32481\,
            I => \N__32461\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__32480\,
            I => \N__32458\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__32479\,
            I => \N__32453\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__32476\,
            I => \N__32448\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32448\
        );

    \I__4487\ : Span4Mux_v
    port map (
            O => \N__32468\,
            I => \N__32445\
        );

    \I__4486\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32442\
        );

    \I__4485\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32429\
        );

    \I__4484\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32429\
        );

    \I__4483\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32429\
        );

    \I__4482\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32429\
        );

    \I__4481\ : InMux
    port map (
            O => \N__32456\,
            I => \N__32429\
        );

    \I__4480\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32429\
        );

    \I__4479\ : Span4Mux_s3_h
    port map (
            O => \N__32448\,
            I => \N__32424\
        );

    \I__4478\ : Span4Mux_v
    port map (
            O => \N__32445\,
            I => \N__32424\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__32442\,
            I => \N__32417\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__32429\,
            I => \N__32417\
        );

    \I__4475\ : Sp12to4
    port map (
            O => \N__32424\,
            I => \N__32417\
        );

    \I__4474\ : Span12Mux_h
    port map (
            O => \N__32417\,
            I => \N__32414\
        );

    \I__4473\ : Odrv12
    port map (
            O => \N__32414\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__32411\,
            I => \N__32408\
        );

    \I__4471\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32405\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__32405\,
            I => \ALU.d_RNI290AE1Z0Z_0\
        );

    \I__4469\ : InMux
    port map (
            O => \N__32402\,
            I => \N__32399\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__32399\,
            I => \ALU.d_RNI5MTIOZ0Z_1\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__32396\,
            I => \busState_1_RNICT0U1_2_cascade_\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__32393\,
            I => \N__32389\
        );

    \I__4465\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32384\
        );

    \I__4464\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32384\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__32384\,
            I => \busState_1_RNICT0U1_2\
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__32381\,
            I => \N_227_0_cascade_\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__32378\,
            I => \N__32375\
        );

    \I__4460\ : InMux
    port map (
            O => \N__32375\,
            I => \N__32372\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__32372\,
            I => \N__32369\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__32369\,
            I => \N__32366\
        );

    \I__4457\ : Span4Mux_h
    port map (
            O => \N__32366\,
            I => \N__32363\
        );

    \I__4456\ : Span4Mux_h
    port map (
            O => \N__32363\,
            I => \N__32360\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__32360\,
            I => \ALU.status_18_cry_2_c_RNOZ0\
        );

    \I__4454\ : CascadeMux
    port map (
            O => \N__32357\,
            I => \N__32354\
        );

    \I__4453\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32351\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__32351\,
            I => \DROM_ROMDATA_dintern_2ro\
        );

    \I__4451\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32342\
        );

    \I__4450\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32342\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__32342\,
            I => \N__32339\
        );

    \I__4448\ : Span4Mux_h
    port map (
            O => \N__32339\,
            I => \N__32336\
        );

    \I__4447\ : Span4Mux_v
    port map (
            O => \N__32336\,
            I => \N__32333\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__32333\,
            I => \DROM.ROMDATA.dintern_0_0_NEW_2\
        );

    \I__4445\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32327\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__32327\,
            I => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_2\
        );

    \I__4443\ : CEMux
    port map (
            O => \N__32324\,
            I => \N__32315\
        );

    \I__4442\ : CEMux
    port map (
            O => \N__32323\,
            I => \N__32312\
        );

    \I__4441\ : InMux
    port map (
            O => \N__32322\,
            I => \N__32309\
        );

    \I__4440\ : CEMux
    port map (
            O => \N__32321\,
            I => \N__32304\
        );

    \I__4439\ : CEMux
    port map (
            O => \N__32320\,
            I => \N__32296\
        );

    \I__4438\ : CEMux
    port map (
            O => \N__32319\,
            I => \N__32290\
        );

    \I__4437\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32290\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__32315\,
            I => \N__32287\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__32312\,
            I => \N__32282\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__32309\,
            I => \N__32282\
        );

    \I__4433\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32277\
        );

    \I__4432\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32277\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__32304\,
            I => \N__32274\
        );

    \I__4430\ : InMux
    port map (
            O => \N__32303\,
            I => \N__32265\
        );

    \I__4429\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32265\
        );

    \I__4428\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32265\
        );

    \I__4427\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32265\
        );

    \I__4426\ : CEMux
    port map (
            O => \N__32299\,
            I => \N__32257\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32254\
        );

    \I__4424\ : InMux
    port map (
            O => \N__32295\,
            I => \N__32251\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__32290\,
            I => \N__32248\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__32287\,
            I => \N__32243\
        );

    \I__4421\ : Span4Mux_h
    port map (
            O => \N__32282\,
            I => \N__32240\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__32277\,
            I => \N__32237\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__32274\,
            I => \N__32232\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32232\
        );

    \I__4417\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32221\
        );

    \I__4416\ : InMux
    port map (
            O => \N__32263\,
            I => \N__32221\
        );

    \I__4415\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32221\
        );

    \I__4414\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32221\
        );

    \I__4413\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32221\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__32257\,
            I => \N__32212\
        );

    \I__4411\ : Span4Mux_v
    port map (
            O => \N__32254\,
            I => \N__32212\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__32251\,
            I => \N__32212\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__32248\,
            I => \N__32212\
        );

    \I__4408\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32207\
        );

    \I__4407\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32207\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__32243\,
            I => \N__32200\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__32240\,
            I => \N__32200\
        );

    \I__4404\ : Span4Mux_h
    port map (
            O => \N__32237\,
            I => \N__32200\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__32232\,
            I => \DROM.ROMDATA.dintern_0_0_sr_enZ0\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__32221\,
            I => \DROM.ROMDATA.dintern_0_0_sr_enZ0\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__32212\,
            I => \DROM.ROMDATA.dintern_0_0_sr_enZ0\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__32207\,
            I => \DROM.ROMDATA.dintern_0_0_sr_enZ0\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__32200\,
            I => \DROM.ROMDATA.dintern_0_0_sr_enZ0\
        );

    \I__4398\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32186\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__32186\,
            I => \ALU.mult_1_12\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__32183\,
            I => \N__32180\
        );

    \I__4395\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32177\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__32177\,
            I => \N__32174\
        );

    \I__4393\ : Span4Mux_v
    port map (
            O => \N__32174\,
            I => \N__32171\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__32171\,
            I => \ALU.mult_3_12\
        );

    \I__4391\ : InMux
    port map (
            O => \N__32168\,
            I => \ALU.mult_17_c11\
        );

    \I__4390\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32162\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__32162\,
            I => \ALU.mult_1_13\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__32159\,
            I => \N__32156\
        );

    \I__4387\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32153\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__32153\,
            I => \N__32150\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__32147\,
            I => \ALU.mult_3_13\
        );

    \I__4383\ : InMux
    port map (
            O => \N__32144\,
            I => \ALU.mult_17_c12\
        );

    \I__4382\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32138\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__32138\,
            I => \ALU.mult_1_14\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__4379\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32129\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__32129\,
            I => \N__32126\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__32126\,
            I => \N__32123\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__32123\,
            I => \ALU.mult_3_14\
        );

    \I__4375\ : InMux
    port map (
            O => \N__32120\,
            I => \ALU.mult_17_c13\
        );

    \I__4374\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__32114\,
            I => \N__32111\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__32111\,
            I => \ALU.mult_227_c_RNIBPRVZ0Z92\
        );

    \I__4371\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32105\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__32105\,
            I => \ALU.mult_83_c_RNIKEU6BZ0Z2\
        );

    \I__4369\ : InMux
    port map (
            O => \N__32102\,
            I => \ALU.mult_17_c14\
        );

    \I__4368\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32096\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__32096\,
            I => \ALU.d_RNIHU6RLZ0Z_1\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__32093\,
            I => \N__32090\
        );

    \I__4365\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32087\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__32087\,
            I => \N__32084\
        );

    \I__4363\ : Span4Mux_h
    port map (
            O => \N__32084\,
            I => \N__32081\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__32081\,
            I => \ALU.d_RNI2E4JE1Z0Z_4\
        );

    \I__4361\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32075\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__32075\,
            I => \N__32072\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__32072\,
            I => \N__32069\
        );

    \I__4358\ : Span4Mux_v
    port map (
            O => \N__32069\,
            I => \N__32066\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__32066\,
            I => \ALU.N_860\
        );

    \I__4356\ : InMux
    port map (
            O => \N__32063\,
            I => \N__32060\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__32060\,
            I => \ALU.mult_5_c_RNOZ0\
        );

    \I__4354\ : InMux
    port map (
            O => \N__32057\,
            I => \N__32054\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__32054\,
            I => \N__32051\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__32051\,
            I => \N__32048\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__32048\,
            I => \ALU.mult_3_4\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__32045\,
            I => \N__32042\
        );

    \I__4349\ : InMux
    port map (
            O => \N__32042\,
            I => \N__32039\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__32039\,
            I => \ALU.mult_1_4\
        );

    \I__4347\ : InMux
    port map (
            O => \N__32036\,
            I => \ALU.mult_17_c3\
        );

    \I__4346\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32030\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__32030\,
            I => \ALU.mult_1_5\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__32027\,
            I => \N__32024\
        );

    \I__4343\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32021\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__32021\,
            I => \N__32018\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__32018\,
            I => \N__32015\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__32015\,
            I => \ALU.mult_3_5\
        );

    \I__4339\ : InMux
    port map (
            O => \N__32012\,
            I => \ALU.mult_17_c4\
        );

    \I__4338\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32006\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__32006\,
            I => \N__32003\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__32003\,
            I => \ALU.mult_1_6\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__32000\,
            I => \N__31997\
        );

    \I__4334\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31994\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__31994\,
            I => \N__31991\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__31991\,
            I => \N__31988\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__31988\,
            I => \ALU.mult_3_6\
        );

    \I__4330\ : InMux
    port map (
            O => \N__31985\,
            I => \ALU.mult_17_c5\
        );

    \I__4329\ : InMux
    port map (
            O => \N__31982\,
            I => \N__31979\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__31979\,
            I => \ALU.mult_1_7\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__31976\,
            I => \N__31973\
        );

    \I__4326\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31970\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__31970\,
            I => \N__31967\
        );

    \I__4324\ : Span4Mux_h
    port map (
            O => \N__31967\,
            I => \N__31964\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__31964\,
            I => \ALU.mult_3_7\
        );

    \I__4322\ : InMux
    port map (
            O => \N__31961\,
            I => \ALU.mult_17_c6\
        );

    \I__4321\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31955\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__31955\,
            I => \ALU.mult_1_8\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__31952\,
            I => \N__31949\
        );

    \I__4318\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31946\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__31946\,
            I => \N__31943\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__31943\,
            I => \N__31940\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__31940\,
            I => \ALU.mult_3_8\
        );

    \I__4314\ : InMux
    port map (
            O => \N__31937\,
            I => \ALU.mult_17_c7\
        );

    \I__4313\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31931\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__31931\,
            I => \N__31928\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__31928\,
            I => \ALU.mult_1_9\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__31925\,
            I => \N__31922\
        );

    \I__4309\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31919\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__31919\,
            I => \N__31916\
        );

    \I__4307\ : Span4Mux_h
    port map (
            O => \N__31916\,
            I => \N__31913\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__31913\,
            I => \ALU.mult_3_9\
        );

    \I__4305\ : InMux
    port map (
            O => \N__31910\,
            I => \ALU.mult_17_c8\
        );

    \I__4304\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31904\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__31904\,
            I => \N__31901\
        );

    \I__4302\ : Odrv12
    port map (
            O => \N__31901\,
            I => \ALU.mult_3_10\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__31898\,
            I => \N__31895\
        );

    \I__4300\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31892\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__31892\,
            I => \ALU.mult_1_10\
        );

    \I__4298\ : InMux
    port map (
            O => \N__31889\,
            I => \bfn_14_11_0_\
        );

    \I__4297\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31883\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__31883\,
            I => \ALU.mult_1_11\
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__31880\,
            I => \N__31877\
        );

    \I__4294\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31874\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__31874\,
            I => \N__31871\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__31871\,
            I => \N__31868\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__31868\,
            I => \ALU.mult_3_11\
        );

    \I__4290\ : InMux
    port map (
            O => \N__31865\,
            I => \ALU.mult_17_c10\
        );

    \I__4289\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31859\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__31859\,
            I => \N__31856\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__31856\,
            I => \N__31853\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__31853\,
            I => \ALU.d_RNIB5POHZ0Z_5\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__31850\,
            I => \N__31847\
        );

    \I__4284\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31844\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__31844\,
            I => \N__31841\
        );

    \I__4282\ : Odrv12
    port map (
            O => \N__31841\,
            I => \ALU.d_RNIPNF141Z0Z_4\
        );

    \I__4281\ : InMux
    port map (
            O => \N__31838\,
            I => \bfn_14_9_0_\
        );

    \I__4280\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31832\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31829\
        );

    \I__4278\ : Odrv12
    port map (
            O => \N__31829\,
            I => \ALU.d_RNI88K161Z0Z_4\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__31826\,
            I => \N__31823\
        );

    \I__4276\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31820\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31817\
        );

    \I__4274\ : Span4Mux_v
    port map (
            O => \N__31817\,
            I => \N__31814\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__31814\,
            I => \ALU.d_RNIMQM8IZ0Z_5\
        );

    \I__4272\ : InMux
    port map (
            O => \N__31811\,
            I => \ALU.mult_5_c13\
        );

    \I__4271\ : InMux
    port map (
            O => \N__31808\,
            I => \N__31805\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__31805\,
            I => \ALU.mult_7_c14_THRU_CO\
        );

    \I__4269\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31799\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__31799\,
            I => \N__31796\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__31796\,
            I => \N__31793\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__31793\,
            I => \N__31790\
        );

    \I__4265\ : Odrv4
    port map (
            O => \N__31790\,
            I => \ALU.d_RNIKDVI51Z0Z_4\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__31787\,
            I => \N__31784\
        );

    \I__4263\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31781\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__31781\,
            I => \N__31778\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__31778\,
            I => \N__31775\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__31775\,
            I => \N__31772\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__31772\,
            I => \ALU.d_RNIRU9M31Z0Z_6\
        );

    \I__4258\ : InMux
    port map (
            O => \N__31769\,
            I => \ALU.mult_5_c14\
        );

    \I__4257\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31763\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__31763\,
            I => \N__31760\
        );

    \I__4255\ : Span4Mux_h
    port map (
            O => \N__31760\,
            I => \N__31757\
        );

    \I__4254\ : Span4Mux_h
    port map (
            O => \N__31757\,
            I => \N__31752\
        );

    \I__4253\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31747\
        );

    \I__4252\ : InMux
    port map (
            O => \N__31755\,
            I => \N__31747\
        );

    \I__4251\ : Sp12to4
    port map (
            O => \N__31752\,
            I => \N__31744\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__31747\,
            I => \N__31741\
        );

    \I__4249\ : Span12Mux_v
    port map (
            O => \N__31744\,
            I => \N__31738\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__31741\,
            I => \N__31735\
        );

    \I__4247\ : Odrv12
    port map (
            O => \N__31738\,
            I => bus_0_12
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__31735\,
            I => bus_0_12
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__31730\,
            I => \N__31727\
        );

    \I__4244\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31724\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__31724\,
            I => \ALU.mult_239_c_RNOZ0Z_0\
        );

    \I__4242\ : InMux
    port map (
            O => \N__31721\,
            I => \N__31718\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__31718\,
            I => \ALU.mult_239_c_RNOZ0\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__31715\,
            I => \N__31711\
        );

    \I__4239\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31706\
        );

    \I__4238\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31706\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__31706\,
            I => \N__31703\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__31703\,
            I => \ALU.mult_1_2\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__31700\,
            I => \N__31697\
        );

    \I__4234\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31694\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__31694\,
            I => \ALU.mult_1_3\
        );

    \I__4232\ : InMux
    port map (
            O => \N__31691\,
            I => \ALU.mult_17_c2\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__31688\,
            I => \N__31685\
        );

    \I__4230\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31682\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__31682\,
            I => \ALU.mult_173_c_RNOZ0Z_0\
        );

    \I__4228\ : InMux
    port map (
            O => \N__31679\,
            I => \ALU.mult_5_c5\
        );

    \I__4227\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31673\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31670\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__31670\,
            I => \ALU.d_RNIFGNR61Z0Z_4\
        );

    \I__4224\ : InMux
    port map (
            O => \N__31667\,
            I => \ALU.mult_5_c6\
        );

    \I__4223\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31661\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__31661\,
            I => \ALU.d_RNICP0UGZ0Z_5\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__31658\,
            I => \N__31655\
        );

    \I__4220\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31652\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__31652\,
            I => \ALU.d_RNI6CL331Z0Z_4\
        );

    \I__4218\ : InMux
    port map (
            O => \N__31649\,
            I => \ALU.mult_5_c7\
        );

    \I__4217\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31643\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__31643\,
            I => \N__31640\
        );

    \I__4215\ : Span4Mux_h
    port map (
            O => \N__31640\,
            I => \N__31637\
        );

    \I__4214\ : Odrv4
    port map (
            O => \N__31637\,
            I => \ALU.d_RNI2RK5IZ0Z_5\
        );

    \I__4213\ : InMux
    port map (
            O => \N__31634\,
            I => \ALU.mult_5_c8\
        );

    \I__4212\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31628\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__31628\,
            I => \N__31625\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__31622\,
            I => \ALU.d_RNIOFVDIZ0Z_5\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__31619\,
            I => \N__31616\
        );

    \I__4207\ : InMux
    port map (
            O => \N__31616\,
            I => \N__31613\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__31613\,
            I => \N__31610\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__31610\,
            I => \ALU.d_RNI5SIF41Z0Z_4\
        );

    \I__4204\ : InMux
    port map (
            O => \N__31607\,
            I => \ALU.mult_5_c9\
        );

    \I__4203\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31601\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__31601\,
            I => \N__31598\
        );

    \I__4201\ : Span4Mux_h
    port map (
            O => \N__31598\,
            I => \N__31595\
        );

    \I__4200\ : Span4Mux_h
    port map (
            O => \N__31595\,
            I => \N__31592\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__31592\,
            I => \ALU.d_RNILKJ1IZ0Z_5\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__31589\,
            I => \N__31586\
        );

    \I__4197\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31583\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__31583\,
            I => \N__31580\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__31577\,
            I => \ALU.d_RNIJTUN21Z0Z_4\
        );

    \I__4193\ : InMux
    port map (
            O => \N__31574\,
            I => \ALU.mult_5_c10\
        );

    \I__4192\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31568\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31565\
        );

    \I__4190\ : Span4Mux_v
    port map (
            O => \N__31565\,
            I => \N__31562\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__31562\,
            I => \ALU.d_RNI6HBMGZ0Z_5\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__31559\,
            I => \N__31556\
        );

    \I__4187\ : InMux
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__31550\,
            I => \N__31547\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__31547\,
            I => \ALU.d_RNI9E4F21Z0Z_4\
        );

    \I__4183\ : InMux
    port map (
            O => \N__31544\,
            I => \ALU.mult_5_c11\
        );

    \I__4182\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31538\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__31538\,
            I => \CONTROL.g1_0\
        );

    \I__4180\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31532\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__31532\,
            I => \N__31528\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__31531\,
            I => \N__31525\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__31528\,
            I => \N__31521\
        );

    \I__4176\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31518\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__31524\,
            I => \N__31515\
        );

    \I__4174\ : Span4Mux_h
    port map (
            O => \N__31521\,
            I => \N__31512\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__31518\,
            I => \N__31509\
        );

    \I__4172\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31506\
        );

    \I__4171\ : Odrv4
    port map (
            O => \N__31512\,
            I => \CONTROL.addrstack_1_1\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__31509\,
            I => \CONTROL.addrstack_1_1\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__31506\,
            I => \CONTROL.addrstack_1_1\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__31499\,
            I => \CONTROL.g1_0_cascade_\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__31496\,
            I => \CONTROL.g0_1_i_a6Z0Z_4_cascade_\
        );

    \I__4166\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31489\
        );

    \I__4165\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31486\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__31489\,
            I => \CONTROL.N_9\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__31486\,
            I => \CONTROL.N_9\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__31481\,
            I => \N__31478\
        );

    \I__4161\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31475\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__31475\,
            I => \N__31472\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__31472\,
            I => \N__31469\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__31469\,
            I => \CONTROL.g0_0_1\
        );

    \I__4157\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31463\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__31463\,
            I => \N__31459\
        );

    \I__4155\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31456\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__31459\,
            I => \N__31451\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__31456\,
            I => \N__31451\
        );

    \I__4152\ : Span4Mux_v
    port map (
            O => \N__31451\,
            I => \N__31448\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__31448\,
            I => \CONTROL.N_366\
        );

    \I__4150\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31441\
        );

    \I__4149\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31438\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__31441\,
            I => \CONTROL.g0_1_i_3\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__31438\,
            I => \CONTROL.g0_1_i_3\
        );

    \I__4146\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31430\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__31430\,
            I => \N__31427\
        );

    \I__4144\ : Odrv12
    port map (
            O => \N__31427\,
            I => \CONTROL.addrstack_15\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__31424\,
            I => \N__31421\
        );

    \I__4142\ : InMux
    port map (
            O => \N__31421\,
            I => \N__31418\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__31418\,
            I => \N__31415\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__31415\,
            I => \CONTROL.addrstack_reto_15\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__31412\,
            I => \N__31408\
        );

    \I__4138\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31405\
        );

    \I__4137\ : InMux
    port map (
            O => \N__31408\,
            I => \N__31401\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__31405\,
            I => \N__31398\
        );

    \I__4135\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31395\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31390\
        );

    \I__4133\ : Span4Mux_h
    port map (
            O => \N__31398\,
            I => \N__31390\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__31395\,
            I => \N__31387\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__31390\,
            I => \N__31384\
        );

    \I__4130\ : Span12Mux_v
    port map (
            O => \N__31387\,
            I => \N__31381\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__31384\,
            I => \controlWord_30\
        );

    \I__4128\ : Odrv12
    port map (
            O => \N__31381\,
            I => \controlWord_30\
        );

    \I__4127\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31373\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31370\
        );

    \I__4125\ : Odrv12
    port map (
            O => \N__31370\,
            I => \PROM.ROMDATA.m471_ns\
        );

    \I__4124\ : InMux
    port map (
            O => \N__31367\,
            I => \N__31364\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__31364\,
            I => \N__31361\
        );

    \I__4122\ : Span4Mux_v
    port map (
            O => \N__31361\,
            I => \N__31358\
        );

    \I__4121\ : Span4Mux_v
    port map (
            O => \N__31358\,
            I => \N__31355\
        );

    \I__4120\ : Sp12to4
    port map (
            O => \N__31355\,
            I => \N__31352\
        );

    \I__4119\ : Span12Mux_h
    port map (
            O => \N__31352\,
            I => \N__31349\
        );

    \I__4118\ : Odrv12
    port map (
            O => \N__31349\,
            I => \gpuOut_c_8\
        );

    \I__4117\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31342\
        );

    \I__4116\ : InMux
    port map (
            O => \N__31345\,
            I => \N__31339\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__31342\,
            I => \CONTROL.ctrlOut_8\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__31339\,
            I => \CONTROL.ctrlOut_8\
        );

    \I__4113\ : IoInMux
    port map (
            O => \N__31334\,
            I => \N__31331\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__31331\,
            I => \N__31328\
        );

    \I__4111\ : IoSpan4Mux
    port map (
            O => \N__31328\,
            I => \N__31325\
        );

    \I__4110\ : Sp12to4
    port map (
            O => \N__31325\,
            I => \N__31322\
        );

    \I__4109\ : Span12Mux_s7_h
    port map (
            O => \N__31322\,
            I => \N__31319\
        );

    \I__4108\ : Span12Mux_v
    port map (
            O => \N__31319\,
            I => \N__31316\
        );

    \I__4107\ : Span12Mux_h
    port map (
            O => \N__31316\,
            I => \N__31313\
        );

    \I__4106\ : Odrv12
    port map (
            O => \N__31313\,
            I => \A0_c\
        );

    \I__4105\ : IoInMux
    port map (
            O => \N__31310\,
            I => \N__31307\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__31307\,
            I => \N__31304\
        );

    \I__4103\ : IoSpan4Mux
    port map (
            O => \N__31304\,
            I => \N__31301\
        );

    \I__4102\ : Span4Mux_s2_h
    port map (
            O => \N__31301\,
            I => \N__31298\
        );

    \I__4101\ : Span4Mux_h
    port map (
            O => \N__31298\,
            I => \N__31295\
        );

    \I__4100\ : Sp12to4
    port map (
            O => \N__31295\,
            I => \N__31291\
        );

    \I__4099\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31288\
        );

    \I__4098\ : Span12Mux_h
    port map (
            O => \N__31291\,
            I => \N__31285\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31282\
        );

    \I__4096\ : Odrv12
    port map (
            O => \N__31285\,
            I => \A1_c\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__31282\,
            I => \A1_c\
        );

    \I__4094\ : InMux
    port map (
            O => \N__31277\,
            I => \N__31272\
        );

    \I__4093\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31269\
        );

    \I__4092\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31266\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__31272\,
            I => \N__31263\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31260\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__31266\,
            I => \N__31257\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__31263\,
            I => \N__31254\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__31260\,
            I => \N__31251\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__31257\,
            I => \N__31246\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__31254\,
            I => \N__31246\
        );

    \I__4084\ : Span4Mux_h
    port map (
            O => \N__31251\,
            I => \N__31243\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__31246\,
            I => \controlWord_26\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__31243\,
            I => \controlWord_26\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__31238\,
            I => \N__31235\
        );

    \I__4080\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31230\
        );

    \I__4079\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31227\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__31233\,
            I => \N__31224\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__31230\,
            I => \N__31221\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31218\
        );

    \I__4075\ : InMux
    port map (
            O => \N__31224\,
            I => \N__31215\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__31221\,
            I => \N__31212\
        );

    \I__4073\ : Span12Mux_v
    port map (
            O => \N__31218\,
            I => \N__31207\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__31215\,
            I => \N__31207\
        );

    \I__4071\ : Odrv4
    port map (
            O => \N__31212\,
            I => \controlWord_27\
        );

    \I__4070\ : Odrv12
    port map (
            O => \N__31207\,
            I => \controlWord_27\
        );

    \I__4069\ : IoInMux
    port map (
            O => \N__31202\,
            I => \N__31199\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__31199\,
            I => \N__31196\
        );

    \I__4067\ : Span12Mux_s9_v
    port map (
            O => \N__31196\,
            I => \N__31193\
        );

    \I__4066\ : Span12Mux_h
    port map (
            O => \N__31193\,
            I => \N__31189\
        );

    \I__4065\ : InMux
    port map (
            O => \N__31192\,
            I => \N__31186\
        );

    \I__4064\ : Odrv12
    port map (
            O => \N__31189\,
            I => \A10_c\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__31186\,
            I => \A10_c\
        );

    \I__4062\ : IoInMux
    port map (
            O => \N__31181\,
            I => \N__31178\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__31178\,
            I => \N__31175\
        );

    \I__4060\ : IoSpan4Mux
    port map (
            O => \N__31175\,
            I => \N__31172\
        );

    \I__4059\ : Sp12to4
    port map (
            O => \N__31172\,
            I => \N__31169\
        );

    \I__4058\ : Span12Mux_s7_h
    port map (
            O => \N__31169\,
            I => \N__31165\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__31168\,
            I => \N__31162\
        );

    \I__4056\ : Span12Mux_h
    port map (
            O => \N__31165\,
            I => \N__31159\
        );

    \I__4055\ : InMux
    port map (
            O => \N__31162\,
            I => \N__31156\
        );

    \I__4054\ : Odrv12
    port map (
            O => \N__31159\,
            I => \A11_c\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__31156\,
            I => \A11_c\
        );

    \I__4052\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31148\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__31148\,
            I => \N__31145\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__31145\,
            I => \N__31142\
        );

    \I__4049\ : Sp12to4
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__4048\ : Odrv12
    port map (
            O => \N__31139\,
            I => \RAM.un1_WR_105_0Z0Z_9\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__31136\,
            I => \N__31133\
        );

    \I__4046\ : InMux
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__31130\,
            I => \N__31127\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__31127\,
            I => \N__31124\
        );

    \I__4043\ : Span4Mux_v
    port map (
            O => \N__31124\,
            I => \N__31120\
        );

    \I__4042\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31117\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__31120\,
            I => \controlWord_25\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__31117\,
            I => \controlWord_25\
        );

    \I__4039\ : IoInMux
    port map (
            O => \N__31112\,
            I => \N__31109\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__31109\,
            I => \N__31106\
        );

    \I__4037\ : Span4Mux_s3_v
    port map (
            O => \N__31106\,
            I => \N__31103\
        );

    \I__4036\ : Span4Mux_h
    port map (
            O => \N__31103\,
            I => \N__31100\
        );

    \I__4035\ : Sp12to4
    port map (
            O => \N__31100\,
            I => \N__31097\
        );

    \I__4034\ : Span12Mux_h
    port map (
            O => \N__31097\,
            I => \N__31093\
        );

    \I__4033\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__4032\ : Odrv12
    port map (
            O => \N__31093\,
            I => \A9_c\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__31090\,
            I => \A9_c\
        );

    \I__4030\ : CascadeMux
    port map (
            O => \N__31085\,
            I => \N__31081\
        );

    \I__4029\ : InMux
    port map (
            O => \N__31084\,
            I => \N__31078\
        );

    \I__4028\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31075\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__31078\,
            I => \N__31072\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__31075\,
            I => \N__31069\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__31072\,
            I => \N__31066\
        );

    \I__4024\ : Span4Mux_v
    port map (
            O => \N__31069\,
            I => \N__31063\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__31066\,
            I => \controlWord_24\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__31063\,
            I => \controlWord_24\
        );

    \I__4021\ : IoInMux
    port map (
            O => \N__31058\,
            I => \N__31055\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__31055\,
            I => \N__31052\
        );

    \I__4019\ : Span4Mux_s3_h
    port map (
            O => \N__31052\,
            I => \N__31049\
        );

    \I__4018\ : Span4Mux_h
    port map (
            O => \N__31049\,
            I => \N__31046\
        );

    \I__4017\ : Span4Mux_h
    port map (
            O => \N__31046\,
            I => \N__31043\
        );

    \I__4016\ : Span4Mux_h
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__31040\,
            I => \N__31036\
        );

    \I__4014\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31033\
        );

    \I__4013\ : Odrv4
    port map (
            O => \N__31036\,
            I => \A8_c\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__31033\,
            I => \A8_c\
        );

    \I__4011\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__31025\,
            I => \N__31022\
        );

    \I__4009\ : Span4Mux_h
    port map (
            O => \N__31022\,
            I => \N__31019\
        );

    \I__4008\ : Span4Mux_v
    port map (
            O => \N__31019\,
            I => \N__31016\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__31016\,
            I => \N__31013\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__31013\,
            I => \gpuOut_c_0\
        );

    \I__4005\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31007\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__4003\ : Span12Mux_v
    port map (
            O => \N__31004\,
            I => \N__31001\
        );

    \I__4002\ : Odrv12
    port map (
            O => \N__31001\,
            I => \D0_in_c\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__30998\,
            I => \CONTROL.N_161_cascade_\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__30995\,
            I => \N__30989\
        );

    \I__3999\ : InMux
    port map (
            O => \N__30994\,
            I => \N__30984\
        );

    \I__3998\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30984\
        );

    \I__3997\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30979\
        );

    \I__3996\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30979\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30976\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__30979\,
            I => \N__30973\
        );

    \I__3993\ : Span4Mux_h
    port map (
            O => \N__30976\,
            I => \N__30970\
        );

    \I__3992\ : Span4Mux_h
    port map (
            O => \N__30973\,
            I => \N__30967\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__30970\,
            I => \PROM.ROMDATA.m520\
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__30967\,
            I => \PROM.ROMDATA.m520\
        );

    \I__3989\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30959\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__30959\,
            I => \N__30956\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__30956\,
            I => \N__30953\
        );

    \I__3986\ : Span4Mux_v
    port map (
            O => \N__30953\,
            I => \N__30950\
        );

    \I__3985\ : Sp12to4
    port map (
            O => \N__30950\,
            I => \N__30947\
        );

    \I__3984\ : Span12Mux_h
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__3983\ : Odrv12
    port map (
            O => \N__30944\,
            I => \gpuOut_c_15\
        );

    \I__3982\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30938\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__30938\,
            I => \N_176\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__30935\,
            I => \N__30931\
        );

    \I__3979\ : InMux
    port map (
            O => \N__30934\,
            I => \N__30928\
        );

    \I__3978\ : InMux
    port map (
            O => \N__30931\,
            I => \N__30925\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__30928\,
            I => \N__30922\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30919\
        );

    \I__3975\ : Span4Mux_h
    port map (
            O => \N__30922\,
            I => \N__30916\
        );

    \I__3974\ : Span4Mux_v
    port map (
            O => \N__30919\,
            I => \N__30913\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__30916\,
            I => \N__30910\
        );

    \I__3972\ : Span4Mux_v
    port map (
            O => \N__30913\,
            I => \N__30907\
        );

    \I__3971\ : Span4Mux_v
    port map (
            O => \N__30910\,
            I => \N__30904\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__30907\,
            I => \N__30901\
        );

    \I__3969\ : Span4Mux_h
    port map (
            O => \N__30904\,
            I => \N__30898\
        );

    \I__3968\ : IoSpan4Mux
    port map (
            O => \N__30901\,
            I => \N__30895\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__30898\,
            I => \D15_in_c\
        );

    \I__3966\ : Odrv4
    port map (
            O => \N__30895\,
            I => \D15_in_c\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__30890\,
            I => \N_176_cascade_\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__30887\,
            I => \CONTROL.N_89_cascade_\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__30884\,
            I => \CONTROL.aluReadBus_1_sqmuxa_0_a2_0Z0Z_0_cascade_\
        );

    \I__3962\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30872\
        );

    \I__3961\ : InMux
    port map (
            O => \N__30880\,
            I => \N__30872\
        );

    \I__3960\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30872\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__30872\,
            I => \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_0\
        );

    \I__3958\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30866\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30863\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__30863\,
            I => \N__30860\
        );

    \I__3955\ : Sp12to4
    port map (
            O => \N__30860\,
            I => \N__30857\
        );

    \I__3954\ : Odrv12
    port map (
            O => \N__30857\,
            I => \gpuOut_c_10\
        );

    \I__3953\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30851\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__30851\,
            I => \N__30848\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__30848\,
            I => \N__30845\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__30845\,
            I => \N__30842\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__30842\,
            I => \N__30839\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__30839\,
            I => \D10_in_c\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__30836\,
            I => \CONTROL.N_171_cascade_\
        );

    \I__3946\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30830\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__30830\,
            I => \N__30827\
        );

    \I__3944\ : Span4Mux_v
    port map (
            O => \N__30827\,
            I => \N__30824\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__30824\,
            I => \CONTROL.N_187\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__30821\,
            I => \CONTROL.un1_busState12_2_i_a2_0_1_tz_0_cascade_\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__30818\,
            I => \CONTROL.N_244_cascade_\
        );

    \I__3940\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30812\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__30812\,
            I => \CONTROL.un1_busState14_1_i_o2_0\
        );

    \I__3938\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30806\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__30806\,
            I => \N__30803\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__30803\,
            I => \CONTROL.aluReadBus_r_1\
        );

    \I__3935\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30797\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__30797\,
            I => \CONTROL.un1_busState14_1_i_a2_1_iZ0Z_1\
        );

    \I__3933\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30784\
        );

    \I__3932\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30784\
        );

    \I__3931\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30781\
        );

    \I__3930\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30778\
        );

    \I__3929\ : InMux
    port map (
            O => \N__30790\,
            I => \N__30773\
        );

    \I__3928\ : InMux
    port map (
            O => \N__30789\,
            I => \N__30773\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__30784\,
            I => \N__30770\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__30781\,
            I => \CONTROL.N_244\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__30778\,
            I => \CONTROL.N_244\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__30773\,
            I => \CONTROL.N_244\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__30770\,
            I => \CONTROL.N_244\
        );

    \I__3922\ : CEMux
    port map (
            O => \N__30761\,
            I => \N__30756\
        );

    \I__3921\ : CEMux
    port map (
            O => \N__30760\,
            I => \N__30753\
        );

    \I__3920\ : CEMux
    port map (
            O => \N__30759\,
            I => \N__30749\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30746\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__30753\,
            I => \N__30743\
        );

    \I__3917\ : CEMux
    port map (
            O => \N__30752\,
            I => \N__30740\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__30749\,
            I => \N__30736\
        );

    \I__3915\ : Span4Mux_v
    port map (
            O => \N__30746\,
            I => \N__30729\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__30743\,
            I => \N__30729\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__30740\,
            I => \N__30729\
        );

    \I__3912\ : CEMux
    port map (
            O => \N__30739\,
            I => \N__30726\
        );

    \I__3911\ : Span4Mux_v
    port map (
            O => \N__30736\,
            I => \N__30723\
        );

    \I__3910\ : Span4Mux_h
    port map (
            O => \N__30729\,
            I => \N__30720\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__30726\,
            I => \N__30717\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__30723\,
            I => \N__30714\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__30720\,
            I => \CONTROL.N_58\
        );

    \I__3906\ : Odrv12
    port map (
            O => \N__30717\,
            I => \CONTROL.N_58\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__30714\,
            I => \CONTROL.N_58\
        );

    \I__3904\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30704\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__30704\,
            I => \CONTROL.N_89\
        );

    \I__3902\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30698\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__30698\,
            I => \N__30695\
        );

    \I__3900\ : Span4Mux_v
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__3899\ : Span4Mux_v
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__3898\ : Span4Mux_v
    port map (
            O => \N__30689\,
            I => \N__30686\
        );

    \I__3897\ : IoSpan4Mux
    port map (
            O => \N__30686\,
            I => \N__30683\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__30683\,
            I => \D11_in_c\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__30680\,
            I => \CONTROL.N_172_cascade_\
        );

    \I__3894\ : InMux
    port map (
            O => \N__30677\,
            I => \N__30674\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__30671\,
            I => \N_188\
        );

    \I__3891\ : InMux
    port map (
            O => \N__30668\,
            I => \N__30665\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30661\
        );

    \I__3889\ : InMux
    port map (
            O => \N__30664\,
            I => \N__30658\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__30661\,
            I => \N_204\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__30658\,
            I => \N_204\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__30653\,
            I => \N_188_cascade_\
        );

    \I__3885\ : InMux
    port map (
            O => \N__30650\,
            I => \N__30647\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__30644\,
            I => \N__30640\
        );

    \I__3882\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30637\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__30640\,
            I => \CONTROL.ctrlOut_11\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__30637\,
            I => \CONTROL.ctrlOut_11\
        );

    \I__3879\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30629\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__30629\,
            I => \N__30626\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__30626\,
            I => \N__30623\
        );

    \I__3876\ : Span4Mux_v
    port map (
            O => \N__30623\,
            I => \N__30620\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__30620\,
            I => \N__30617\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__30617\,
            I => \N__30614\
        );

    \I__3873\ : Odrv4
    port map (
            O => \N__30614\,
            I => \gpuOut_c_12\
        );

    \I__3872\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30608\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__30608\,
            I => \N__30605\
        );

    \I__3870\ : Span4Mux_v
    port map (
            O => \N__30605\,
            I => \N__30602\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__30602\,
            I => \N__30599\
        );

    \I__3868\ : Span4Mux_v
    port map (
            O => \N__30599\,
            I => \N__30596\
        );

    \I__3867\ : Span4Mux_h
    port map (
            O => \N__30596\,
            I => \N__30593\
        );

    \I__3866\ : Odrv4
    port map (
            O => \N__30593\,
            I => \D12_in_c\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__30590\,
            I => \CONTROL.N_173_cascade_\
        );

    \I__3864\ : InMux
    port map (
            O => \N__30587\,
            I => \N__30584\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__30584\,
            I => \CONTROL.N_189\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__30581\,
            I => \CONTROL.un1_busState14_1_i_o2_0_cascade_\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__30578\,
            I => \CONTROL.busState_1_RNIRA1I6Z0Z_2_cascade_\
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__30575\,
            I => \N__30572\
        );

    \I__3859\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30569\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__30569\,
            I => \N__30566\
        );

    \I__3857\ : Span4Mux_v
    port map (
            O => \N__30566\,
            I => \N__30563\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__30563\,
            I => \ALU.d_RNI8VHNHZ0Z_1\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__30560\,
            I => \ALU.dout_3_ns_1_12_cascade_\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__30557\,
            I => \ALU.dout_6_ns_1_12_cascade_\
        );

    \I__3853\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30551\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__30551\,
            I => \ALU.N_1097\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__30548\,
            I => \ALU.N_1145_cascade_\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__30545\,
            I => \aluOut_12_cascade_\
        );

    \I__3849\ : InMux
    port map (
            O => \N__30542\,
            I => \N__30536\
        );

    \I__3848\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30536\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__30536\,
            I => \N__30533\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__30533\,
            I => \N__30530\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__30530\,
            I => \CONTROL.bus_0_12\
        );

    \I__3844\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30524\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__3842\ : Span4Mux_h
    port map (
            O => \N__30521\,
            I => \N__30518\
        );

    \I__3841\ : Span4Mux_v
    port map (
            O => \N__30518\,
            I => \N__30515\
        );

    \I__3840\ : Span4Mux_v
    port map (
            O => \N__30515\,
            I => \N__30512\
        );

    \I__3839\ : Span4Mux_v
    port map (
            O => \N__30512\,
            I => \N__30509\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__30509\,
            I => \N__30506\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__30506\,
            I => \gpuOut_c_11\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__30503\,
            I => \N__30500\
        );

    \I__3835\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30497\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__30497\,
            I => \N__30494\
        );

    \I__3833\ : Odrv12
    port map (
            O => \N__30494\,
            I => \ALU.mult_5_c_RNOZ0Z_0\
        );

    \I__3832\ : InMux
    port map (
            O => \N__30491\,
            I => \N__30485\
        );

    \I__3831\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30485\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__30485\,
            I => \N__30482\
        );

    \I__3829\ : Span4Mux_h
    port map (
            O => \N__30482\,
            I => \N__30479\
        );

    \I__3828\ : Span4Mux_h
    port map (
            O => \N__30479\,
            I => \N__30476\
        );

    \I__3827\ : Odrv4
    port map (
            O => \N__30476\,
            I => \DROM.ROMDATA.dintern_0_0_NEW_0\
        );

    \I__3826\ : InMux
    port map (
            O => \N__30473\,
            I => \N__30470\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__30470\,
            I => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_0\
        );

    \I__3824\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30464\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__30464\,
            I => \N__30461\
        );

    \I__3822\ : Span12Mux_v
    port map (
            O => \N__30461\,
            I => \N__30458\
        );

    \I__3821\ : Span12Mux_h
    port map (
            O => \N__30458\,
            I => \N__30455\
        );

    \I__3820\ : Odrv12
    port map (
            O => \N__30455\,
            I => \gpuOut_c_14\
        );

    \I__3819\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30449\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__30449\,
            I => \N__30446\
        );

    \I__3817\ : Span12Mux_h
    port map (
            O => \N__30446\,
            I => \N__30442\
        );

    \I__3816\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30439\
        );

    \I__3815\ : Odrv12
    port map (
            O => \N__30442\,
            I => \CONTROL.ctrlOut_14\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__30439\,
            I => \CONTROL.ctrlOut_14\
        );

    \I__3813\ : InMux
    port map (
            O => \N__30434\,
            I => \N__30431\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__30431\,
            I => \N__30428\
        );

    \I__3811\ : Span4Mux_h
    port map (
            O => \N__30428\,
            I => \N__30425\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__30425\,
            I => \N__30422\
        );

    \I__3809\ : Sp12to4
    port map (
            O => \N__30422\,
            I => \N__30419\
        );

    \I__3808\ : Span12Mux_v
    port map (
            O => \N__30419\,
            I => \N__30416\
        );

    \I__3807\ : Odrv12
    port map (
            O => \N__30416\,
            I => \D14_in_c\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__30413\,
            I => \CONTROL.N_175_cascade_\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__30410\,
            I => \N_191_cascade_\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__30407\,
            I => \N__30403\
        );

    \I__3803\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30400\
        );

    \I__3802\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30397\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__30400\,
            I => \N__30394\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30391\
        );

    \I__3799\ : Span4Mux_h
    port map (
            O => \N__30394\,
            I => \N__30388\
        );

    \I__3798\ : Span4Mux_h
    port map (
            O => \N__30391\,
            I => \N__30383\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__30388\,
            I => \N__30383\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__30380\,
            I => \CONTROL_addrstack_reto_11\
        );

    \I__3794\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30374\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__30374\,
            I => \N__30370\
        );

    \I__3792\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30367\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__30370\,
            I => \N__30364\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__30367\,
            I => \N__30361\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__30364\,
            I => \N__30358\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__30361\,
            I => \N__30355\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__30358\,
            I => \N_426\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__30355\,
            I => \N_426\
        );

    \I__3785\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30347\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30343\
        );

    \I__3783\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30340\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__30343\,
            I => \N__30335\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__30340\,
            I => \N__30335\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__30335\,
            I => \N__30332\
        );

    \I__3779\ : Span4Mux_h
    port map (
            O => \N__30332\,
            I => \N__30329\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__30329\,
            I => \progRomAddress_11\
        );

    \I__3777\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30323\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__30323\,
            I => \N__30320\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__30320\,
            I => \N__30317\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__30317\,
            I => \ALU.d_RNILJMRC1_0Z0Z_8\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__30314\,
            I => \ALU.combOperand2_1Z0Z_0_cascade_\
        );

    \I__3772\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30308\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__3770\ : Span4Mux_v
    port map (
            O => \N__30305\,
            I => \N__30302\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__30302\,
            I => dintern_adflt_3_x
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__30299\,
            I => \DROM_ROMDATA_dintern_0ro_cascade_\
        );

    \I__3767\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30293\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30290\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__30290\,
            I => \N__30287\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__30287\,
            I => \CONTROL.bus_6_a0_sx_0\
        );

    \I__3763\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30281\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__30281\,
            I => \ALU.mult_3_c14_THRU_CO\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__30278\,
            I => \N__30275\
        );

    \I__3760\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__30269\,
            I => \N__30266\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__30266\,
            I => \ALU.d_RNI3D2O61Z0Z_2\
        );

    \I__3756\ : InMux
    port map (
            O => \N__30263\,
            I => \ALU.mult_1_c14\
        );

    \I__3755\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__30257\,
            I => \ALU.d_RNI83GO51Z0Z_0\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__30254\,
            I => \N__30251\
        );

    \I__3752\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30248\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__30248\,
            I => \ALU.d_RNIPIBO31Z0Z_0\
        );

    \I__3750\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30242\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__30242\,
            I => \N__30239\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__30239\,
            I => \ALU.d_RNIIHC6LZ0Z_3\
        );

    \I__3747\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30233\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__30233\,
            I => \ALU.d_RNITH0K51Z0Z_0\
        );

    \I__3745\ : InMux
    port map (
            O => \N__30230\,
            I => \N__30227\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__30227\,
            I => \N__30224\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__30224\,
            I => \ALU.d_RNI0H41KZ0Z_1\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__30221\,
            I => \N__30218\
        );

    \I__3741\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30215\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__30215\,
            I => \ALU.d_RNIETL861Z0Z_0\
        );

    \I__3739\ : InMux
    port map (
            O => \N__30212\,
            I => \N__30209\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__30209\,
            I => \ALU.d_RNI8FM541Z0Z_0\
        );

    \I__3737\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30203\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__30203\,
            I => \N__30200\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__30200\,
            I => \ALU.d_RNIGIF4D1Z0Z_2\
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__30197\,
            I => \N__30194\
        );

    \I__3733\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30191\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__30191\,
            I => \N__30188\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__30188\,
            I => \ALU.d_RNIRJ3VHZ0Z_1\
        );

    \I__3730\ : InMux
    port map (
            O => \N__30185\,
            I => \ALU.mult_1_c6\
        );

    \I__3729\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30179\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__30179\,
            I => \N__30176\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__30176\,
            I => \N__30173\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__30173\,
            I => \ALU.d_RNI990621Z0Z_0\
        );

    \I__3725\ : InMux
    port map (
            O => \N__30170\,
            I => \ALU.mult_1_c7\
        );

    \I__3724\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__30164\,
            I => \ALU.d_RNIH49MHZ0Z_1\
        );

    \I__3722\ : InMux
    port map (
            O => \N__30161\,
            I => \bfn_13_12_0_\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__30158\,
            I => \N__30155\
        );

    \I__3720\ : InMux
    port map (
            O => \N__30155\,
            I => \N__30152\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__30152\,
            I => \N__30149\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__30149\,
            I => \ALU.d_RNISP66IZ0Z_1\
        );

    \I__3717\ : InMux
    port map (
            O => \N__30146\,
            I => \ALU.mult_1_c9\
        );

    \I__3716\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30137\
        );

    \I__3714\ : Span4Mux_h
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__30134\,
            I => \ALU.d_RNI0LDMJZ0Z_1\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__30131\,
            I => \N__30128\
        );

    \I__3711\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30125\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__30125\,
            I => \ALU.d_RNIK8R951Z0Z_0\
        );

    \I__3709\ : InMux
    port map (
            O => \N__30122\,
            I => \ALU.mult_1_c10\
        );

    \I__3708\ : InMux
    port map (
            O => \N__30119\,
            I => \ALU.mult_1_c11\
        );

    \I__3707\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30113\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__30113\,
            I => \N__30110\
        );

    \I__3705\ : Span4Mux_v
    port map (
            O => \N__30110\,
            I => \N__30107\
        );

    \I__3704\ : Odrv4
    port map (
            O => \N__30107\,
            I => \ALU.d_RNI9UI0KZ0Z_1\
        );

    \I__3703\ : InMux
    port map (
            O => \N__30104\,
            I => \ALU.mult_1_c12\
        );

    \I__3702\ : InMux
    port map (
            O => \N__30101\,
            I => \ALU.mult_1_c13\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__30098\,
            I => \N__30095\
        );

    \I__3700\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30092\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__30092\,
            I => \N__30089\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__30089\,
            I => \ALU.d_RNIA6P2IZ0Z_7\
        );

    \I__3697\ : InMux
    port map (
            O => \N__30086\,
            I => \ALU.mult_1_c1\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__30083\,
            I => \N__30080\
        );

    \I__3695\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30077\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__30077\,
            I => \ALU.d_RNIFBJI61Z0Z_0\
        );

    \I__3693\ : InMux
    port map (
            O => \N__30074\,
            I => \ALU.mult_1_c2\
        );

    \I__3692\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30068\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__30068\,
            I => \ALU.d_RNIIOGRGZ0Z_1\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__30065\,
            I => \N__30062\
        );

    \I__3689\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30059\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__30059\,
            I => \N__30056\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__30056\,
            I => \N__30053\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__30053\,
            I => \ALU.d_RNI67HQ21Z0Z_0\
        );

    \I__3685\ : InMux
    port map (
            O => \N__30050\,
            I => \ALU.mult_1_c3\
        );

    \I__3684\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__30044\,
            I => \N__30041\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__30041\,
            I => \N__30038\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__30038\,
            I => \ALU.d_RNI8Q43IZ0Z_1\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30032\
        );

    \I__3679\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__30029\,
            I => \N__30026\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__30026\,
            I => \ALU.d_RNIITFA41Z0Z_0\
        );

    \I__3676\ : InMux
    port map (
            O => \N__30023\,
            I => \ALU.mult_1_c4\
        );

    \I__3675\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30017\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__30017\,
            I => \N__30014\
        );

    \I__3673\ : Span4Mux_h
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__30011\,
            I => \ALU.d_RNI5NE641Z0Z_0\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__30008\,
            I => \N__30005\
        );

    \I__3670\ : InMux
    port map (
            O => \N__30005\,
            I => \N__30002\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__3668\ : Odrv12
    port map (
            O => \N__29999\,
            I => \ALU.d_RNIUEFBIZ0Z_1\
        );

    \I__3667\ : InMux
    port map (
            O => \N__29996\,
            I => \ALU.mult_1_c5\
        );

    \I__3666\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29990\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__29990\,
            I => \ALU.d_RNIUFQIGZ0Z_7\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__3663\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__29981\,
            I => \N__29978\
        );

    \I__3661\ : Span4Mux_v
    port map (
            O => \N__29978\,
            I => \N__29975\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__3659\ : Odrv4
    port map (
            O => \N__29972\,
            I => \ALU.d_RNI8JFO21Z0Z_6\
        );

    \I__3658\ : InMux
    port map (
            O => \N__29969\,
            I => \ALU.mult_7_c9\
        );

    \I__3657\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29963\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__29963\,
            I => \N__29960\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__29960\,
            I => \N__29957\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__29957\,
            I => \N__29954\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__29954\,
            I => \ALU.d_RNIKHEQHZ0Z_7\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__29951\,
            I => \N__29948\
        );

    \I__3651\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__29945\,
            I => \N__29942\
        );

    \I__3649\ : Span4Mux_v
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__3648\ : Sp12to4
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__3647\ : Odrv12
    port map (
            O => \N__29936\,
            I => \ALU.d_RNIK9E841Z0Z_6\
        );

    \I__3646\ : InMux
    port map (
            O => \N__29933\,
            I => \ALU.mult_7_c10\
        );

    \I__3645\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29927\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__29927\,
            I => \N__29924\
        );

    \I__3643\ : Span4Mux_v
    port map (
            O => \N__29924\,
            I => \N__29921\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__29921\,
            I => \N__29918\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__29918\,
            I => \ALU.d_RNI73D441Z0Z_6\
        );

    \I__3640\ : InMux
    port map (
            O => \N__29915\,
            I => \ALU.mult_7_c11\
        );

    \I__3639\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29909\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__29909\,
            I => \N__29906\
        );

    \I__3637\ : Span4Mux_v
    port map (
            O => \N__29906\,
            I => \N__29903\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__29903\,
            I => \ALU.d_RNI7BDMHZ0Z_7\
        );

    \I__3635\ : InMux
    port map (
            O => \N__29900\,
            I => \ALU.mult_7_c12\
        );

    \I__3634\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29894\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__29894\,
            I => \N__29891\
        );

    \I__3632\ : Span4Mux_v
    port map (
            O => \N__29891\,
            I => \N__29888\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__29888\,
            I => \ALU.d_RNIBLU321Z0Z_6\
        );

    \I__3630\ : InMux
    port map (
            O => \N__29885\,
            I => \ALU.mult_7_c13\
        );

    \I__3629\ : InMux
    port map (
            O => \N__29882\,
            I => \bfn_13_10_0_\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__29879\,
            I => \N__29876\
        );

    \I__3627\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29873\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__29873\,
            I => \ALU.d_RNIHNHG61Z0Z_6\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__3624\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29864\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__29864\,
            I => \ALU.d_RNI4LU7E1Z0Z_6\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__29861\,
            I => \ALU.d_RNILJMRC1Z0Z_8_cascade_\
        );

    \I__3621\ : InMux
    port map (
            O => \N__29858\,
            I => \ALU.mult_7_c7\
        );

    \I__3620\ : InMux
    port map (
            O => \N__29855\,
            I => \N__29852\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__29852\,
            I => \ALU.d_RNITLGILZ0Z_7\
        );

    \I__3618\ : InMux
    port map (
            O => \N__29849\,
            I => \ALU.mult_7_c8\
        );

    \I__3617\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__29843\,
            I => \N__29839\
        );

    \I__3615\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29836\
        );

    \I__3614\ : Span4Mux_v
    port map (
            O => \N__29839\,
            I => \N__29833\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__29836\,
            I => \N__29830\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__29833\,
            I => \CONTROL.programCounter_1_10\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__29830\,
            I => \CONTROL.programCounter_1_10\
        );

    \I__3610\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29818\
        );

    \I__3609\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29815\
        );

    \I__3608\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29808\
        );

    \I__3607\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29808\
        );

    \I__3606\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29808\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__29818\,
            I => \CONTROL.programCounter11_reto_rep1\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__29815\,
            I => \CONTROL.programCounter11_reto_rep1\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__29808\,
            I => \CONTROL.programCounter11_reto_rep1\
        );

    \I__3602\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__29798\,
            I => \CONTROL.programCounter_1_reto_10\
        );

    \I__3600\ : InMux
    port map (
            O => \N__29795\,
            I => \N__29792\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__29792\,
            I => \CONTROL.N_425\
        );

    \I__3598\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29786\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__29786\,
            I => \N__29783\
        );

    \I__3596\ : Span4Mux_h
    port map (
            O => \N__29783\,
            I => \N__29780\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__29780\,
            I => \CONTROL.programCounter_1_axb_1\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__3593\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__29771\,
            I => \N__29768\
        );

    \I__3591\ : Odrv12
    port map (
            O => \N__29768\,
            I => \CONTROL.addrstackptr_8_1\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__29765\,
            I => \N__29762\
        );

    \I__3589\ : InMux
    port map (
            O => \N__29762\,
            I => \N__29759\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__29759\,
            I => \N__29756\
        );

    \I__3587\ : Odrv12
    port map (
            O => \N__29756\,
            I => \CONTROL.addrstackptr_RNI19JNL91Z0Z_0\
        );

    \I__3586\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29750\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__29750\,
            I => \CONTROL.dout_reto_9\
        );

    \I__3584\ : CascadeMux
    port map (
            O => \N__29747\,
            I => \N__29744\
        );

    \I__3583\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__29741\,
            I => \N__29737\
        );

    \I__3581\ : InMux
    port map (
            O => \N__29740\,
            I => \N__29734\
        );

    \I__3580\ : Span4Mux_v
    port map (
            O => \N__29737\,
            I => \N__29731\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__29734\,
            I => \progRomAddress_15\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__29731\,
            I => \progRomAddress_15\
        );

    \I__3577\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29723\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29719\
        );

    \I__3575\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29716\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__29719\,
            I => \N__29713\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__29716\,
            I => \CONTROL.programCounter_1_11\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__29713\,
            I => \CONTROL.programCounter_1_11\
        );

    \I__3571\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29704\
        );

    \I__3570\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29701\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29695\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29695\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__29700\,
            I => \N__29692\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__29695\,
            I => \N__29689\
        );

    \I__3565\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29686\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__29689\,
            I => \CONTROL.addrstack_1_4\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__29686\,
            I => \CONTROL.addrstack_1_4\
        );

    \I__3562\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29678\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__29678\,
            I => \CONTROL.N_4_1\
        );

    \I__3560\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29671\
        );

    \I__3559\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29668\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__29671\,
            I => \CONTROL.un1_addrstackptr_c4_0\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__29668\,
            I => \CONTROL.un1_addrstackptr_c4_0\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__3555\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29657\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__29657\,
            I => \N__29654\
        );

    \I__3553\ : Span4Mux_h
    port map (
            O => \N__29654\,
            I => \N__29651\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__29651\,
            I => \CONTROL.addrstackptr_8_4\
        );

    \I__3551\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29644\
        );

    \I__3550\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29641\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__29644\,
            I => \N__29638\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__29641\,
            I => \CONTROL.programCounter_1_14\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__29638\,
            I => \CONTROL.programCounter_1_14\
        );

    \I__3546\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29630\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__29630\,
            I => \CONTROL.programCounter_1_reto_14\
        );

    \I__3544\ : InMux
    port map (
            O => \N__29627\,
            I => \N__29624\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__29624\,
            I => \CONTROL.programCounter_1_reto_11\
        );

    \I__3542\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29618\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__29618\,
            I => \CONTROL.dout_reto_11\
        );

    \I__3540\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29612\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__29612\,
            I => \N__29609\
        );

    \I__3538\ : Span4Mux_h
    port map (
            O => \N__29609\,
            I => \N__29606\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__29606\,
            I => \PROM.ROMDATA.m470_am\
        );

    \I__3536\ : InMux
    port map (
            O => \N__29603\,
            I => \N__29600\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__29600\,
            I => \CONTROL.dout_reto_14\
        );

    \I__3534\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29593\
        );

    \I__3533\ : InMux
    port map (
            O => \N__29596\,
            I => \N__29590\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__29593\,
            I => \N__29587\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__29590\,
            I => \N__29584\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__29587\,
            I => \controlWord_18\
        );

    \I__3529\ : Odrv4
    port map (
            O => \N__29584\,
            I => \controlWord_18\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__29579\,
            I => \controlWord_18_cascade_\
        );

    \I__3527\ : IoInMux
    port map (
            O => \N__29576\,
            I => \N__29573\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__29573\,
            I => \N__29570\
        );

    \I__3525\ : IoSpan4Mux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__3524\ : Span4Mux_s0_h
    port map (
            O => \N__29567\,
            I => \N__29564\
        );

    \I__3523\ : Sp12to4
    port map (
            O => \N__29564\,
            I => \N__29561\
        );

    \I__3522\ : Span12Mux_s8_h
    port map (
            O => \N__29561\,
            I => \N__29558\
        );

    \I__3521\ : Span12Mux_h
    port map (
            O => \N__29558\,
            I => \N__29554\
        );

    \I__3520\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29551\
        );

    \I__3519\ : Odrv12
    port map (
            O => \N__29554\,
            I => \A2_c\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__29551\,
            I => \A2_c\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__29546\,
            I => \CONTROL.g0_3_i_1_0_cascade_\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__29543\,
            I => \CONTROL.N_4_1_cascade_\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__29540\,
            I => \N__29536\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__29539\,
            I => \N__29533\
        );

    \I__3513\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29528\
        );

    \I__3512\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29528\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__29528\,
            I => \N__29525\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__29525\,
            I => \N__29522\
        );

    \I__3509\ : Span4Mux_h
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__29519\,
            I => \CONTROL.N_81_0\
        );

    \I__3507\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29513\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__29513\,
            I => \CONTROL.g0_3_i_a7_2_0\
        );

    \I__3505\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29507\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__29507\,
            I => \CONTROL.N_429\
        );

    \I__3503\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29501\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__29501\,
            I => \CONTROL.dout_reto_8\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__29498\,
            I => \CONTROL.gpuWrite_RNOZ0Z_2_cascade_\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__29495\,
            I => \CONTROL.busState96_cascade_\
        );

    \I__3499\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29489\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__29489\,
            I => \CONTROL.busState96\
        );

    \I__3497\ : InMux
    port map (
            O => \N__29486\,
            I => \N__29483\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__29483\,
            I => \CONTROL.N_66_0\
        );

    \I__3495\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29477\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__29477\,
            I => \CONTROL.gpuWrite_RNOZ0Z_0\
        );

    \I__3493\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29470\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__29473\,
            I => \N__29467\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__29470\,
            I => \N__29464\
        );

    \I__3490\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29461\
        );

    \I__3489\ : Odrv12
    port map (
            O => \N__29464\,
            I => \gpuWrite\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__29461\,
            I => \gpuWrite\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__29456\,
            I => \N__29452\
        );

    \I__3486\ : InMux
    port map (
            O => \N__29455\,
            I => \N__29448\
        );

    \I__3485\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29445\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__29451\,
            I => \N__29442\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__29448\,
            I => \N__29439\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__29445\,
            I => \N__29436\
        );

    \I__3481\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29433\
        );

    \I__3480\ : Span4Mux_v
    port map (
            O => \N__29439\,
            I => \N__29430\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__29436\,
            I => \N__29425\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__29433\,
            I => \N__29425\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__29430\,
            I => \N__29420\
        );

    \I__3476\ : Span4Mux_v
    port map (
            O => \N__29425\,
            I => \N__29420\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__29420\,
            I => \controlWord_21\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__29417\,
            I => \RAM.un1_WR_105_0Z0Z_3_cascade_\
        );

    \I__3473\ : IoInMux
    port map (
            O => \N__29414\,
            I => \N__29411\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__29411\,
            I => \N__29408\
        );

    \I__3471\ : Span4Mux_s2_v
    port map (
            O => \N__29408\,
            I => \N__29405\
        );

    \I__3470\ : Span4Mux_h
    port map (
            O => \N__29405\,
            I => \N__29402\
        );

    \I__3469\ : Sp12to4
    port map (
            O => \N__29402\,
            I => \N__29399\
        );

    \I__3468\ : Span12Mux_h
    port map (
            O => \N__29399\,
            I => \N__29395\
        );

    \I__3467\ : InMux
    port map (
            O => \N__29398\,
            I => \N__29392\
        );

    \I__3466\ : Odrv12
    port map (
            O => \N__29395\,
            I => \A5_c\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__29392\,
            I => \A5_c\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__29387\,
            I => \N__29384\
        );

    \I__3463\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__29381\,
            I => \N__29378\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__29378\,
            I => \N__29375\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__29375\,
            I => \N__29372\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__29372\,
            I => \RAM.un1_WR_105_0Z0Z_11\
        );

    \I__3458\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29365\
        );

    \I__3457\ : InMux
    port map (
            O => \N__29368\,
            I => \N__29362\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__29365\,
            I => \N__29359\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__29362\,
            I => \controlWord_23\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__29359\,
            I => \controlWord_23\
        );

    \I__3453\ : IoInMux
    port map (
            O => \N__29354\,
            I => \N__29351\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__29351\,
            I => \N__29348\
        );

    \I__3451\ : Span12Mux_s8_h
    port map (
            O => \N__29348\,
            I => \N__29345\
        );

    \I__3450\ : Span12Mux_h
    port map (
            O => \N__29345\,
            I => \N__29341\
        );

    \I__3449\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29338\
        );

    \I__3448\ : Odrv12
    port map (
            O => \N__29341\,
            I => \A7_c\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__29338\,
            I => \A7_c\
        );

    \I__3446\ : IoInMux
    port map (
            O => \N__29333\,
            I => \N__29330\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__29330\,
            I => \N__29327\
        );

    \I__3444\ : IoSpan4Mux
    port map (
            O => \N__29327\,
            I => \N__29324\
        );

    \I__3443\ : Span4Mux_s3_h
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__3442\ : Sp12to4
    port map (
            O => \N__29321\,
            I => \N__29318\
        );

    \I__3441\ : Span12Mux_s11_h
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__3440\ : Odrv12
    port map (
            O => \N__29315\,
            I => \gpuAddress_3\
        );

    \I__3439\ : IoInMux
    port map (
            O => \N__29312\,
            I => \N__29309\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__29309\,
            I => \N__29306\
        );

    \I__3437\ : IoSpan4Mux
    port map (
            O => \N__29306\,
            I => \N__29303\
        );

    \I__3436\ : Span4Mux_s0_h
    port map (
            O => \N__29303\,
            I => \N__29300\
        );

    \I__3435\ : Sp12to4
    port map (
            O => \N__29300\,
            I => \N__29297\
        );

    \I__3434\ : Span12Mux_s11_h
    port map (
            O => \N__29297\,
            I => \N__29294\
        );

    \I__3433\ : Span12Mux_v
    port map (
            O => \N__29294\,
            I => \N__29291\
        );

    \I__3432\ : Odrv12
    port map (
            O => \N__29291\,
            I => \gpuAddress_4\
        );

    \I__3431\ : IoInMux
    port map (
            O => \N__29288\,
            I => \N__29285\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29282\
        );

    \I__3429\ : Span4Mux_s0_h
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__3428\ : Span4Mux_h
    port map (
            O => \N__29279\,
            I => \N__29276\
        );

    \I__3427\ : Sp12to4
    port map (
            O => \N__29276\,
            I => \N__29273\
        );

    \I__3426\ : Span12Mux_v
    port map (
            O => \N__29273\,
            I => \N__29270\
        );

    \I__3425\ : Odrv12
    port map (
            O => \N__29270\,
            I => \gpuAddress_5\
        );

    \I__3424\ : IoInMux
    port map (
            O => \N__29267\,
            I => \N__29264\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__29264\,
            I => \N__29261\
        );

    \I__3422\ : Span12Mux_s3_h
    port map (
            O => \N__29261\,
            I => \N__29258\
        );

    \I__3421\ : Span12Mux_v
    port map (
            O => \N__29258\,
            I => \N__29255\
        );

    \I__3420\ : Odrv12
    port map (
            O => \N__29255\,
            I => \gpuAddress_6\
        );

    \I__3419\ : IoInMux
    port map (
            O => \N__29252\,
            I => \N__29249\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__29249\,
            I => \N__29246\
        );

    \I__3417\ : Span12Mux_s2_h
    port map (
            O => \N__29246\,
            I => \N__29243\
        );

    \I__3416\ : Span12Mux_h
    port map (
            O => \N__29243\,
            I => \N__29240\
        );

    \I__3415\ : Span12Mux_v
    port map (
            O => \N__29240\,
            I => \N__29237\
        );

    \I__3414\ : Odrv12
    port map (
            O => \N__29237\,
            I => \gpuAddress_7\
        );

    \I__3413\ : IoInMux
    port map (
            O => \N__29234\,
            I => \N__29231\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29228\
        );

    \I__3411\ : IoSpan4Mux
    port map (
            O => \N__29228\,
            I => \N__29225\
        );

    \I__3410\ : Span4Mux_s2_h
    port map (
            O => \N__29225\,
            I => \N__29222\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__29222\,
            I => \N__29219\
        );

    \I__3408\ : Span4Mux_v
    port map (
            O => \N__29219\,
            I => \N__29216\
        );

    \I__3407\ : Span4Mux_h
    port map (
            O => \N__29216\,
            I => \N__29213\
        );

    \I__3406\ : Span4Mux_h
    port map (
            O => \N__29213\,
            I => \N__29210\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__29210\,
            I => \gpuAddress_8\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__29207\,
            I => \CONTROL.un1_busState119_1_i_0_1_cascade_\
        );

    \I__3403\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29201\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__29201\,
            I => \N__29198\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__29198\,
            I => \N__29195\
        );

    \I__3400\ : Span4Mux_v
    port map (
            O => \N__29195\,
            I => \N__29192\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__29192\,
            I => \N__29189\
        );

    \I__3398\ : IoSpan4Mux
    port map (
            O => \N__29189\,
            I => \N__29186\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__29186\,
            I => \gpuOut_c_7\
        );

    \I__3396\ : InMux
    port map (
            O => \N__29183\,
            I => \N__29180\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__29180\,
            I => \N_168\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__29177\,
            I => \N_168_cascade_\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__29174\,
            I => \N__29170\
        );

    \I__3392\ : InMux
    port map (
            O => \N__29173\,
            I => \N__29165\
        );

    \I__3391\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29165\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__29165\,
            I => \N__29162\
        );

    \I__3389\ : Span4Mux_v
    port map (
            O => \N__29162\,
            I => \N__29159\
        );

    \I__3388\ : Span4Mux_v
    port map (
            O => \N__29159\,
            I => \N__29156\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__3386\ : Span4Mux_v
    port map (
            O => \N__29153\,
            I => \N__29150\
        );

    \I__3385\ : IoSpan4Mux
    port map (
            O => \N__29150\,
            I => \N__29147\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__29147\,
            I => \D7_in_c\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__29144\,
            I => \CONTROL.bus_7_ns_1_7_cascade_\
        );

    \I__3382\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29135\
        );

    \I__3381\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29135\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__29135\,
            I => \N__29132\
        );

    \I__3379\ : Span4Mux_v
    port map (
            O => \N__29132\,
            I => \N__29129\
        );

    \I__3378\ : Span4Mux_h
    port map (
            O => \N__29129\,
            I => \N__29126\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__29126\,
            I => \PROM_ROMDATA_dintern_23ro\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__29123\,
            I => \CONTROL.bus_7_a1_1_8_cascade_\
        );

    \I__3375\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29117\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__29117\,
            I => \N__29114\
        );

    \I__3373\ : Span4Mux_v
    port map (
            O => \N__29114\,
            I => \N__29111\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__29111\,
            I => \CONTROL.bus_sx_8\
        );

    \I__3371\ : IoInMux
    port map (
            O => \N__29108\,
            I => \N__29105\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29102\
        );

    \I__3369\ : Span4Mux_s3_h
    port map (
            O => \N__29102\,
            I => \N__29099\
        );

    \I__3368\ : Span4Mux_h
    port map (
            O => \N__29099\,
            I => \N__29096\
        );

    \I__3367\ : Sp12to4
    port map (
            O => \N__29096\,
            I => \N__29093\
        );

    \I__3366\ : Span12Mux_v
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__3365\ : Odrv12
    port map (
            O => \N__29090\,
            I => \gpuAddress_2\
        );

    \I__3364\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29084\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__29084\,
            I => \ALU.c_RNI3MHFZ0Z_11\
        );

    \I__3362\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29078\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__29078\,
            I => \ALU.dout_3_ns_1_11\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__29075\,
            I => \ALU.dout_3_ns_1_10_cascade_\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__29072\,
            I => \ALU.dout_6_ns_1_10_cascade_\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__29069\,
            I => \ALU.N_1143_cascade_\
        );

    \I__3357\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29063\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__29063\,
            I => \ALU.N_1095\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__29060\,
            I => \aluOut_10_cascade_\
        );

    \I__3354\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29053\
        );

    \I__3353\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29050\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__29053\,
            I => \N__29047\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__29050\,
            I => \N__29044\
        );

    \I__3350\ : Span4Mux_v
    port map (
            O => \N__29047\,
            I => \N__29041\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__29044\,
            I => \N__29038\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__29041\,
            I => \CONTROL.bus_0_10\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__29038\,
            I => \CONTROL.bus_0_10\
        );

    \I__3346\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29030\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__29030\,
            I => \ALU_N_1141\
        );

    \I__3344\ : InMux
    port map (
            O => \N__29027\,
            I => \N__29023\
        );

    \I__3343\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29020\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__29023\,
            I => \ALU_N_1093\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__29020\,
            I => \ALU_N_1093\
        );

    \I__3340\ : InMux
    port map (
            O => \N__29015\,
            I => \N__29012\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__29012\,
            I => \ALU.N_1144\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__29009\,
            I => \ALU.N_1096_cascade_\
        );

    \I__3337\ : InMux
    port map (
            O => \N__29006\,
            I => \N__29003\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__29003\,
            I => \N__29000\
        );

    \I__3335\ : Span4Mux_h
    port map (
            O => \N__29000\,
            I => \N__28997\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__28997\,
            I => \DROM_ROMDATA_dintern_11ro\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__28994\,
            I => \aluOut_11_cascade_\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__28991\,
            I => \ALU.operand2_7_ns_1_11_cascade_\
        );

    \I__3331\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28985\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28982\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__28982\,
            I => \ALU.b_RNI2TJC1Z0Z_11\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__28979\,
            I => \ALU.operand2_11_cascade_\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__28976\,
            I => \ALU.d_RNIMR627Z0Z_11_cascade_\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__28973\,
            I => \N__28970\
        );

    \I__3325\ : InMux
    port map (
            O => \N__28970\,
            I => \N__28967\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__28967\,
            I => \ALU.a_RNIV5PUZ0Z_11\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__28964\,
            I => \N__28961\
        );

    \I__3322\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28958\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__28958\,
            I => \N__28955\
        );

    \I__3320\ : Odrv12
    port map (
            O => \N__28955\,
            I => \ALU.d_RNI9IN2HZ0Z_3\
        );

    \I__3319\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28949\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__28949\,
            I => \N__28946\
        );

    \I__3317\ : Span4Mux_v
    port map (
            O => \N__28946\,
            I => \N__28943\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__28943\,
            I => \ALU.a_RNI2N741Z0Z_12\
        );

    \I__3315\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28937\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__28937\,
            I => \N__28934\
        );

    \I__3313\ : Span4Mux_v
    port map (
            O => \N__28934\,
            I => \N__28930\
        );

    \I__3312\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28927\
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__28930\,
            I => \ALU.d_RNIJRM75Z0Z_5\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__28927\,
            I => \ALU.d_RNIJRM75Z0Z_5\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__28922\,
            I => \N__28917\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__28921\,
            I => \N__28914\
        );

    \I__3307\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28911\
        );

    \I__3306\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28908\
        );

    \I__3305\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28905\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28902\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__28908\,
            I => \N__28899\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28896\
        );

    \I__3301\ : Span4Mux_h
    port map (
            O => \N__28902\,
            I => \N__28891\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__28899\,
            I => \N__28891\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__28896\,
            I => \N__28888\
        );

    \I__3298\ : Span4Mux_v
    port map (
            O => \N__28891\,
            I => \N__28885\
        );

    \I__3297\ : Span4Mux_v
    port map (
            O => \N__28888\,
            I => \N__28882\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__28885\,
            I => \DROM_ROMDATA_dintern_5ro\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__28882\,
            I => \DROM_ROMDATA_dintern_5ro\
        );

    \I__3294\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28873\
        );

    \I__3293\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28870\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28867\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28864\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__28867\,
            I => \ALU.d_RNIC0VE6Z0Z_5\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__28864\,
            I => \ALU.d_RNIC0VE6Z0Z_5\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__28859\,
            I => \N__28856\
        );

    \I__3287\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__28853\,
            I => \N__28850\
        );

    \I__3285\ : Odrv12
    port map (
            O => \N__28850\,
            I => \ALU.d_RNI693UNZ0Z_3\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__3283\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28838\
        );

    \I__3281\ : Odrv12
    port map (
            O => \N__28838\,
            I => \ALU.mult_95_c_RNOZ0Z_0\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__28835\,
            I => \ALU.dout_6_ns_1_11_cascade_\
        );

    \I__3279\ : InMux
    port map (
            O => \N__28832\,
            I => \ALU.mult_3_c14\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__28829\,
            I => \N__28826\
        );

    \I__3277\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28823\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__28823\,
            I => \ALU.d_RNI2IA441Z0Z_2\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__28820\,
            I => \N__28817\
        );

    \I__3274\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28814\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28811\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__28811\,
            I => \ALU.d_RNI7SQI21Z0Z_2\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__28808\,
            I => \N__28805\
        );

    \I__3270\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28802\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__3268\ : Odrv12
    port map (
            O => \N__28799\,
            I => \ALU.d_RNID31VFZ0Z_3\
        );

    \I__3267\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28793\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__28793\,
            I => \ALU.d_RNIBRFE41Z0Z_2\
        );

    \I__3265\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28787\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__28787\,
            I => \ALU.d_RNI9DAEHZ0Z_3\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__28784\,
            I => \N__28781\
        );

    \I__3262\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28778\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N__28775\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__28775\,
            I => \ALU.d_RNI07V431Z0Z_2\
        );

    \I__3259\ : InMux
    port map (
            O => \N__28772\,
            I => \ALU.mult_3_c6\
        );

    \I__3258\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__28766\,
            I => \ALU.d_RNIJ0U031Z0Z_2\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__28763\,
            I => \N__28760\
        );

    \I__3255\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28757\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__28757\,
            I => \ALU.d_RNIV1LMHZ0Z_3\
        );

    \I__3253\ : InMux
    port map (
            O => \N__28754\,
            I => \ALU.mult_3_c7\
        );

    \I__3252\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__28748\,
            I => \ALU.d_RNIS69AHZ0Z_3\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__28745\,
            I => \N__28742\
        );

    \I__3249\ : InMux
    port map (
            O => \N__28742\,
            I => \N__28739\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__28739\,
            I => \ALU.d_RNI12A911Z0Z_2\
        );

    \I__3247\ : InMux
    port map (
            O => \N__28736\,
            I => \ALU.mult_3_c8\
        );

    \I__3246\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28730\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__28730\,
            I => \ALU.d_RNINIF011Z0Z_2\
        );

    \I__3244\ : InMux
    port map (
            O => \N__28727\,
            I => \ALU.mult_3_c9\
        );

    \I__3243\ : InMux
    port map (
            O => \N__28724\,
            I => \N__28721\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28718\
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__28718\,
            I => \ALU.d_RNIINE1HZ0Z_3\
        );

    \I__3240\ : InMux
    port map (
            O => \N__28715\,
            I => \bfn_12_12_0_\
        );

    \I__3239\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28709\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__28709\,
            I => \N__28706\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__28706\,
            I => \N__28703\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__28703\,
            I => \ALU.d_RNIMCVI41Z0Z_2\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__28700\,
            I => \N__28697\
        );

    \I__3234\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28694\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__28694\,
            I => \N__28691\
        );

    \I__3232\ : Span4Mux_v
    port map (
            O => \N__28691\,
            I => \N__28688\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__28688\,
            I => \ALU.d_RNITCCHHZ0Z_3\
        );

    \I__3230\ : InMux
    port map (
            O => \N__28685\,
            I => \ALU.mult_3_c11\
        );

    \I__3229\ : InMux
    port map (
            O => \N__28682\,
            I => \N__28679\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__28679\,
            I => \N__28676\
        );

    \I__3227\ : Span4Mux_h
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__28673\,
            I => \N__28670\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__28670\,
            I => \ALU.d_RNI18J1JZ0Z_3\
        );

    \I__3224\ : InMux
    port map (
            O => \N__28667\,
            I => \ALU.mult_3_c12\
        );

    \I__3223\ : InMux
    port map (
            O => \N__28664\,
            I => \ALU.mult_3_c13\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__28661\,
            I => \ALU.status_19_2_cascade_\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__28658\,
            I => \N__28655\
        );

    \I__3220\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28652\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__28652\,
            I => \N__28649\
        );

    \I__3218\ : Span4Mux_h
    port map (
            O => \N__28649\,
            I => \N__28646\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__28646\,
            I => \N__28643\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__28643\,
            I => \romOut_4\
        );

    \I__3215\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28637\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__28637\,
            I => \N__28634\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__28634\,
            I => \CONTROL.busState_1_RNI7U266Z0Z_2\
        );

    \I__3212\ : InMux
    port map (
            O => \N__28631\,
            I => \ALU.mult_3_c3\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__28628\,
            I => \N__28625\
        );

    \I__3210\ : InMux
    port map (
            O => \N__28625\,
            I => \N__28622\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__28622\,
            I => \ALU.d_RNITK2D51Z0Z_2\
        );

    \I__3208\ : InMux
    port map (
            O => \N__28619\,
            I => \ALU.mult_3_c4\
        );

    \I__3207\ : InMux
    port map (
            O => \N__28616\,
            I => \N__28613\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__28613\,
            I => \ALU.d_RNIJBM6GZ0Z_3\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__28610\,
            I => \N__28607\
        );

    \I__3204\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28604\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__28604\,
            I => \ALU.d_RNIKG0L11Z0Z_2\
        );

    \I__3202\ : InMux
    port map (
            O => \N__28601\,
            I => \ALU.mult_3_c5\
        );

    \I__3201\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28595\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__28595\,
            I => \N__28592\
        );

    \I__3199\ : Span4Mux_v
    port map (
            O => \N__28592\,
            I => \N__28589\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__28589\,
            I => \ALU.status_17_I_1_c_RNOZ0\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__28586\,
            I => \ALU.N_834_cascade_\
        );

    \I__3196\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28580\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28577\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__28577\,
            I => \N__28573\
        );

    \I__3193\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28570\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__28573\,
            I => \N__28567\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__28570\,
            I => \busState_1_RNIDU0U1_2\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__28567\,
            I => \busState_1_RNIDU0U1_2\
        );

    \I__3189\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28559\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__28559\,
            I => \CONTROL.programCounter_1_reto_9\
        );

    \I__3187\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28553\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__28553\,
            I => \CONTROL.addrstack_reto_9\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__28550\,
            I => \CONTROL.N_424_cascade_\
        );

    \I__3184\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28544\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__28544\,
            I => \N__28541\
        );

    \I__3182\ : Odrv12
    port map (
            O => \N__28541\,
            I => \progRomAddress_9\
        );

    \I__3181\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28532\
        );

    \I__3180\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28532\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__28532\,
            I => \CONTROL_addrstack_reto_8\
        );

    \I__3178\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__28526\,
            I => \N_423\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__28523\,
            I => \progRomAddress_9_cascade_\
        );

    \I__3175\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28514\
        );

    \I__3174\ : InMux
    port map (
            O => \N__28519\,
            I => \N__28514\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__28511\,
            I => \N__28508\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__28508\,
            I => \PROM.ROMDATA.dintern_adfltZ0Z_3\
        );

    \I__3170\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28502\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__28502\,
            I => \N__28499\
        );

    \I__3168\ : Odrv12
    port map (
            O => \N__28499\,
            I => \CONTROL.tempCounterZ0Z_10\
        );

    \I__3167\ : InMux
    port map (
            O => \N__28496\,
            I => \N__28492\
        );

    \I__3166\ : InMux
    port map (
            O => \N__28495\,
            I => \N__28489\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28484\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__28489\,
            I => \N__28484\
        );

    \I__3163\ : Odrv12
    port map (
            O => \N__28484\,
            I => \CONTROL.programCounter_1_9\
        );

    \I__3162\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28478\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__28478\,
            I => \N__28475\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__28475\,
            I => \CONTROL.tempCounterZ0Z_9\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__3158\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__28466\,
            I => \ALU.rshift_3_ns_1_2\
        );

    \I__3156\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28460\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__28460\,
            I => \N__28457\
        );

    \I__3154\ : Span4Mux_v
    port map (
            O => \N__28457\,
            I => \N__28454\
        );

    \I__3153\ : Span4Mux_h
    port map (
            O => \N__28454\,
            I => \N__28451\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__28451\,
            I => \CONTROL.addrstack_13\
        );

    \I__3151\ : InMux
    port map (
            O => \N__28448\,
            I => \N__28445\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__28445\,
            I => \CONTROL.addrstack_reto_13\
        );

    \I__3149\ : InMux
    port map (
            O => \N__28442\,
            I => \N__28435\
        );

    \I__3148\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28435\
        );

    \I__3147\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28432\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__28435\,
            I => \N__28429\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__28432\,
            I => \progRomAddress_10\
        );

    \I__3144\ : Odrv12
    port map (
            O => \N__28429\,
            I => \progRomAddress_10\
        );

    \I__3143\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28421\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__28421\,
            I => \CONTROL.addrstack_reto_12\
        );

    \I__3141\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28414\
        );

    \I__3140\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28411\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__28414\,
            I => \N__28408\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__28411\,
            I => \progRomAddress_12\
        );

    \I__3137\ : Odrv12
    port map (
            O => \N__28408\,
            I => \progRomAddress_12\
        );

    \I__3136\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28400\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__28400\,
            I => \N__28397\
        );

    \I__3134\ : Span4Mux_h
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__28394\,
            I => \CONTROL.addrstack_10\
        );

    \I__3132\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28388\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__28388\,
            I => \CONTROL.addrstack_reto_10\
        );

    \I__3130\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28382\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__28382\,
            I => \CONTROL.programCounter_1_reto_8\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__28379\,
            I => \N_423_cascade_\
        );

    \I__3127\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28373\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__28373\,
            I => \N__28370\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__28370\,
            I => \CONTROL.programCounter_1_axb_8\
        );

    \I__3124\ : CEMux
    port map (
            O => \N__28367\,
            I => \N__28364\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__28364\,
            I => \N__28361\
        );

    \I__3122\ : Span4Mux_v
    port map (
            O => \N__28361\,
            I => \N__28358\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__28358\,
            I => \CONTROL.programCounter10\
        );

    \I__3120\ : InMux
    port map (
            O => \N__28355\,
            I => \CONTROL.programCounter_1_cry_11\
        );

    \I__3119\ : InMux
    port map (
            O => \N__28352\,
            I => \CONTROL.programCounter_1_cry_12\
        );

    \I__3118\ : InMux
    port map (
            O => \N__28349\,
            I => \CONTROL.programCounter_1_cry_13\
        );

    \I__3117\ : InMux
    port map (
            O => \N__28346\,
            I => \CONTROL.programCounter_1_cry_14\
        );

    \I__3116\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28339\
        );

    \I__3115\ : InMux
    port map (
            O => \N__28342\,
            I => \N__28336\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__28339\,
            I => \N__28333\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__28336\,
            I => \N__28328\
        );

    \I__3112\ : Span4Mux_h
    port map (
            O => \N__28333\,
            I => \N__28328\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__28328\,
            I => \CONTROL.programCounter_1_13\
        );

    \I__3110\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28322\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__28322\,
            I => \CONTROL.programCounter_1_reto_13\
        );

    \I__3108\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28316\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__28316\,
            I => \CONTROL.dout_reto_13\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__28313\,
            I => \CONTROL.N_428_cascade_\
        );

    \I__3105\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28306\
        );

    \I__3104\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28303\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__28306\,
            I => \N__28300\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__28303\,
            I => \progRomAddress_13\
        );

    \I__3101\ : Odrv12
    port map (
            O => \N__28300\,
            I => \progRomAddress_13\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__3099\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28289\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__28289\,
            I => \CONTROL.addrstack_reto_14\
        );

    \I__3097\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28282\
        );

    \I__3096\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28279\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__28282\,
            I => \N__28276\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__28279\,
            I => \progRomAddress_14\
        );

    \I__3093\ : Odrv12
    port map (
            O => \N__28276\,
            I => \progRomAddress_14\
        );

    \I__3092\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28268\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__3090\ : Span4Mux_v
    port map (
            O => \N__28265\,
            I => \N__28262\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__28262\,
            I => \CONTROL.programCounter_1_axb_3\
        );

    \I__3088\ : InMux
    port map (
            O => \N__28259\,
            I => \CONTROL.programCounter_1_cry_2\
        );

    \I__3087\ : InMux
    port map (
            O => \N__28256\,
            I => \CONTROL.programCounter_1_cry_3\
        );

    \I__3086\ : InMux
    port map (
            O => \N__28253\,
            I => \CONTROL.programCounter_1_cry_4\
        );

    \I__3085\ : InMux
    port map (
            O => \N__28250\,
            I => \CONTROL.programCounter_1_cry_5\
        );

    \I__3084\ : InMux
    port map (
            O => \N__28247\,
            I => \CONTROL.programCounter_1_cry_6\
        );

    \I__3083\ : InMux
    port map (
            O => \N__28244\,
            I => \bfn_11_22_0_\
        );

    \I__3082\ : InMux
    port map (
            O => \N__28241\,
            I => \CONTROL.programCounter_1_cry_8\
        );

    \I__3081\ : InMux
    port map (
            O => \N__28238\,
            I => \CONTROL.programCounter_1_cry_9\
        );

    \I__3080\ : InMux
    port map (
            O => \N__28235\,
            I => \CONTROL.programCounter_1_cry_10\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__28232\,
            I => \controlWord_29_cascade_\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__28229\,
            I => \N__28225\
        );

    \I__3077\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28222\
        );

    \I__3076\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28219\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__28222\,
            I => \N__28216\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__28219\,
            I => \N__28213\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__28216\,
            I => \controlWord_28\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__28213\,
            I => \controlWord_28\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__28208\,
            I => \controlWord_28_cascade_\
        );

    \I__3070\ : IoInMux
    port map (
            O => \N__28205\,
            I => \N__28202\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__28202\,
            I => \N__28199\
        );

    \I__3068\ : IoSpan4Mux
    port map (
            O => \N__28199\,
            I => \N__28196\
        );

    \I__3067\ : Span4Mux_s2_h
    port map (
            O => \N__28196\,
            I => \N__28193\
        );

    \I__3066\ : Sp12to4
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__3065\ : Span12Mux_h
    port map (
            O => \N__28190\,
            I => \N__28187\
        );

    \I__3064\ : Span12Mux_v
    port map (
            O => \N__28187\,
            I => \N__28183\
        );

    \I__3063\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28180\
        );

    \I__3062\ : Odrv12
    port map (
            O => \N__28183\,
            I => \A12_c\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__28180\,
            I => \A12_c\
        );

    \I__3060\ : IoInMux
    port map (
            O => \N__28175\,
            I => \N__28172\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__28172\,
            I => \N__28169\
        );

    \I__3058\ : Span4Mux_s3_v
    port map (
            O => \N__28169\,
            I => \N__28166\
        );

    \I__3057\ : Span4Mux_h
    port map (
            O => \N__28166\,
            I => \N__28163\
        );

    \I__3056\ : Sp12to4
    port map (
            O => \N__28163\,
            I => \N__28160\
        );

    \I__3055\ : Span12Mux_h
    port map (
            O => \N__28160\,
            I => \N__28156\
        );

    \I__3054\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28153\
        );

    \I__3053\ : Odrv12
    port map (
            O => \N__28156\,
            I => \A13_c\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__28153\,
            I => \A13_c\
        );

    \I__3051\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28145\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__28145\,
            I => \N__28142\
        );

    \I__3049\ : Span4Mux_v
    port map (
            O => \N__28142\,
            I => \N__28139\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__28139\,
            I => \RAM.un1_WR_105_0Z0Z_10\
        );

    \I__3047\ : InMux
    port map (
            O => \N__28136\,
            I => \CONTROL.programCounter_1_cry_0\
        );

    \I__3046\ : InMux
    port map (
            O => \N__28133\,
            I => \CONTROL.programCounter_1_cry_1\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__28130\,
            I => \CONTROL.busState_1_e_1_0_cascade_\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__28127\,
            I => \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0_cascade_\
        );

    \I__3043\ : CEMux
    port map (
            O => \N__28124\,
            I => \N__28119\
        );

    \I__3042\ : CEMux
    port map (
            O => \N__28123\,
            I => \N__28116\
        );

    \I__3041\ : CEMux
    port map (
            O => \N__28122\,
            I => \N__28113\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28105\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__28116\,
            I => \N__28105\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__28113\,
            I => \N__28102\
        );

    \I__3037\ : CEMux
    port map (
            O => \N__28112\,
            I => \N__28099\
        );

    \I__3036\ : CEMux
    port map (
            O => \N__28111\,
            I => \N__28096\
        );

    \I__3035\ : CEMux
    port map (
            O => \N__28110\,
            I => \N__28093\
        );

    \I__3034\ : Span4Mux_v
    port map (
            O => \N__28105\,
            I => \N__28086\
        );

    \I__3033\ : Span4Mux_v
    port map (
            O => \N__28102\,
            I => \N__28086\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__28099\,
            I => \N__28086\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__28096\,
            I => \N_29\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__28093\,
            I => \N_29\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__28086\,
            I => \N_29\
        );

    \I__3028\ : InMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__28076\,
            I => \CONTROL.N_352\
        );

    \I__3026\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__28070\,
            I => \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0\
        );

    \I__3024\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28064\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__28064\,
            I => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_3\
        );

    \I__3022\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28058\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__28058\,
            I => \N__28054\
        );

    \I__3020\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28051\
        );

    \I__3019\ : Span4Mux_h
    port map (
            O => \N__28054\,
            I => \N__28048\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__28051\,
            I => \N__28045\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__28048\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_3\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__28045\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_3\
        );

    \I__3015\ : InMux
    port map (
            O => \N__28040\,
            I => \N__28037\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__28037\,
            I => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_0\
        );

    \I__3013\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28030\
        );

    \I__3012\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28027\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__28030\,
            I => \N__28024\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__28027\,
            I => \N__28021\
        );

    \I__3009\ : Span4Mux_h
    port map (
            O => \N__28024\,
            I => \N__28018\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__28021\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_0\
        );

    \I__3007\ : Odrv4
    port map (
            O => \N__28018\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_0\
        );

    \I__3006\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28007\
        );

    \I__3005\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28007\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__28004\,
            I => \N__28000\
        );

    \I__3002\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27997\
        );

    \I__3001\ : Span4Mux_v
    port map (
            O => \N__28000\,
            I => \N__27994\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__27997\,
            I => \DROM_ROMDATA_dintern_4ro\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__27994\,
            I => \DROM_ROMDATA_dintern_4ro\
        );

    \I__2998\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27985\
        );

    \I__2997\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27982\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27979\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__27982\,
            I => \N__27976\
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__27979\,
            I => \controlWord_29\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__27976\,
            I => \controlWord_29\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__27971\,
            I => \ALU.dout_3_ns_1_8_cascade_\
        );

    \I__2991\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__27965\,
            I => \ALU.c_RNIFT2SZ0Z_8\
        );

    \I__2989\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__2987\ : Span4Mux_h
    port map (
            O => \N__27956\,
            I => \N__27950\
        );

    \I__2986\ : InMux
    port map (
            O => \N__27955\,
            I => \N__27943\
        );

    \I__2985\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27943\
        );

    \I__2984\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27943\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__27950\,
            I => \dataRomAddress_10\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__27943\,
            I => \dataRomAddress_10\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__27938\,
            I => \N__27933\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__27937\,
            I => \N__27930\
        );

    \I__2979\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27927\
        );

    \I__2978\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27922\
        );

    \I__2977\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27922\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__27927\,
            I => \dataRomAddress_12\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__27922\,
            I => \dataRomAddress_12\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__27917\,
            I => \PROM.ROMDATA.dintern_adfltZ0Z_4_cascade_\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__27914\,
            I => \PROM.ROMDATA.dintern_12dflt_0Z0Z_1_cascade_\
        );

    \I__2972\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27908\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__27908\,
            I => \PROM.ROMDATA.dintern_adfltZ0Z_4\
        );

    \I__2970\ : InMux
    port map (
            O => \N__27905\,
            I => \N__27902\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__27902\,
            I => \N__27899\
        );

    \I__2968\ : Span12Mux_v
    port map (
            O => \N__27899\,
            I => \N__27893\
        );

    \I__2967\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27890\
        );

    \I__2966\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27885\
        );

    \I__2965\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27885\
        );

    \I__2964\ : Odrv12
    port map (
            O => \N__27893\,
            I => \dataRomAddress_11\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__27890\,
            I => \dataRomAddress_11\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__27885\,
            I => \dataRomAddress_11\
        );

    \I__2961\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27875\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__27875\,
            I => \ALU.c_RNIAMVQZ0Z_6\
        );

    \I__2959\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27869\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__27869\,
            I => \ALU.d_RNIDV8EZ0Z_6\
        );

    \I__2957\ : InMux
    port map (
            O => \N__27866\,
            I => \N__27863\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__27863\,
            I => \ALU.c_RNI230LZ0Z_10\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__27860\,
            I => \ALU.a_RNIUI741Z0Z_10_cascade_\
        );

    \I__2954\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27854\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__27854\,
            I => \ALU.operand2_7_ns_1_10\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__27851\,
            I => \ALU.dout_6_ns_1_8_cascade_\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__27848\,
            I => \ALU_N_1141_cascade_\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__27845\,
            I => \CONTROL.bus_0_sx_8_cascade_\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__27842\,
            I => \N__27839\
        );

    \I__2948\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27836\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__27836\,
            I => \N__27832\
        );

    \I__2946\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27829\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__27832\,
            I => \CONTROL_bus_0_8\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__27829\,
            I => \CONTROL_bus_0_8\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__27824\,
            I => \ALU.status_19_8_cascade_\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__27821\,
            I => \ALU.operand2_7_ns_1_6_cascade_\
        );

    \I__2941\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__27815\,
            I => \ALU.operand2_6\
        );

    \I__2939\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27809\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__27809\,
            I => \ALU.b_RNI9JSPZ0Z_6\
        );

    \I__2937\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27803\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__27803\,
            I => \ALU.e_RNI6AJMZ0Z_6\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__27800\,
            I => \ALU.operand2_7_ns_1_4_cascade_\
        );

    \I__2934\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27794\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__27794\,
            I => \ALU.operand2_4\
        );

    \I__2932\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27788\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__27788\,
            I => \ALU.c_RNI6IVQZ0Z_4\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__27785\,
            I => \ALU.dout_6_ns_1_4_cascade_\
        );

    \I__2929\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27778\
        );

    \I__2928\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27775\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__27778\,
            I => \ALU.aZ0Z_4\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__27775\,
            I => \ALU.aZ0Z_4\
        );

    \I__2925\ : CascadeMux
    port map (
            O => \N__27770\,
            I => \ALU.dout_3_ns_1_4_cascade_\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__27767\,
            I => \ALU.N_1089_cascade_\
        );

    \I__2923\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27761\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__27761\,
            I => \ALU.N_1137\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__27758\,
            I => \aluOut_4_cascade_\
        );

    \I__2920\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27749\
        );

    \I__2919\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27749\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__27749\,
            I => \ALU.d_RNIBJM75Z0Z_4\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__27746\,
            I => \ALU.addsub_cry_3_c_RNIGCKVJZ0Z5_cascade_\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__27743\,
            I => \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9_cascade_\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__27740\,
            I => \ALU.e_RNI26JMZ0Z_4_cascade_\
        );

    \I__2914\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27734\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__27734\,
            I => \N__27731\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__27731\,
            I => \N__27728\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__27728\,
            I => \CONTROL.tempCounterZ0Z_11\
        );

    \I__2910\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27722\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__27722\,
            I => \N__27719\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__27719\,
            I => \N__27716\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__27716\,
            I => \CONTROL.tempCounterZ0Z_15\
        );

    \I__2906\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27710\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27707\
        );

    \I__2904\ : Span4Mux_v
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__27704\,
            I => \CONTROL.tempCounterZ0Z_14\
        );

    \I__2902\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__27698\,
            I => \N__27695\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__27695\,
            I => \CONTROL.addrstack_8\
        );

    \I__2899\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27689\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__27689\,
            I => \N__27686\
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__27686\,
            I => \CONTROL.addrstack_9\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__27683\,
            I => \N__27680\
        );

    \I__2895\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27677\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__27677\,
            I => \N__27674\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__27674\,
            I => \ALU.status_17_I_9_c_RNOZ0\
        );

    \I__2892\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27668\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__27668\,
            I => \CONTROL.g0_3_iZ0Z_1\
        );

    \I__2890\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27662\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__27662\,
            I => \CONTROL.g0_3_i_a7Z0Z_2\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__27659\,
            I => \N__27656\
        );

    \I__2887\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27653\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__27653\,
            I => \N__27650\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__27650\,
            I => \CONTROL.g0_0_2\
        );

    \I__2884\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27644\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__27644\,
            I => \N__27641\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__27641\,
            I => \N__27638\
        );

    \I__2881\ : Span4Mux_h
    port map (
            O => \N__27638\,
            I => \N__27635\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__27635\,
            I => \CONTROL.addrstack_12\
        );

    \I__2879\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27629\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__27629\,
            I => \N__27626\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__27626\,
            I => \N__27623\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__27623\,
            I => \CONTROL.addrstack_11\
        );

    \I__2875\ : InMux
    port map (
            O => \N__27620\,
            I => \N__27617\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__27617\,
            I => \N__27614\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__27611\,
            I => \CONTROL.addrstack_7\
        );

    \I__2871\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__27605\,
            I => \N__27602\
        );

    \I__2869\ : Span4Mux_h
    port map (
            O => \N__27602\,
            I => \N__27599\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__27599\,
            I => \CONTROL.addrstack_14\
        );

    \I__2867\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27593\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__27593\,
            I => \N__27590\
        );

    \I__2865\ : Span4Mux_v
    port map (
            O => \N__27590\,
            I => \N__27587\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__27587\,
            I => \N__27584\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__27584\,
            I => \N__27581\
        );

    \I__2862\ : Sp12to4
    port map (
            O => \N__27581\,
            I => \N__27578\
        );

    \I__2861\ : Odrv12
    port map (
            O => \N__27578\,
            I => \D6_in_c\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__27575\,
            I => \CONTROL.N_167_cascade_\
        );

    \I__2859\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27568\
        );

    \I__2858\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27565\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__27568\,
            I => \N__27562\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N_183\
        );

    \I__2855\ : Odrv12
    port map (
            O => \N__27562\,
            I => \N_183\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__27557\,
            I => \CONTROL.addrstackptr_N_8_mux_1_0_cascade_\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__2852\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27548\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__27542\,
            I => \CONTROL.addrstackptr_N_6_0_1_i\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__27539\,
            I => \CONTROL.g0_3_i_2_cascade_\
        );

    \I__2847\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__27533\,
            I => \CONTROL.N_4_0\
        );

    \I__2845\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27523\
        );

    \I__2844\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27523\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__27528\,
            I => \N__27520\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__27523\,
            I => \N__27517\
        );

    \I__2841\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__27517\,
            I => \CONTROL.addrstack_1_5\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__27514\,
            I => \CONTROL.addrstack_1_5\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__27509\,
            I => \CONTROL.N_4_0_cascade_\
        );

    \I__2837\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27503\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__27503\,
            I => \CONTROL.addrstackptr_N_8_mux_1_0\
        );

    \I__2835\ : InMux
    port map (
            O => \N__27500\,
            I => \N__27495\
        );

    \I__2834\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27488\
        );

    \I__2833\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27488\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27485\
        );

    \I__2831\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27480\
        );

    \I__2830\ : InMux
    port map (
            O => \N__27493\,
            I => \N__27480\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__27488\,
            I => \N__27477\
        );

    \I__2828\ : Span4Mux_h
    port map (
            O => \N__27485\,
            I => \N__27474\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__27480\,
            I => \CONTROL.addrstackptrZ0Z_5\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__27477\,
            I => \CONTROL.addrstackptrZ0Z_5\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__27474\,
            I => \CONTROL.addrstackptrZ0Z_5\
        );

    \I__2824\ : InMux
    port map (
            O => \N__27467\,
            I => \N__27463\
        );

    \I__2823\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27460\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__27463\,
            I => \N__27457\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__27460\,
            I => \N__27454\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__27457\,
            I => \N__27451\
        );

    \I__2819\ : Span4Mux_h
    port map (
            O => \N__27454\,
            I => \N__27448\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__27451\,
            I => \DROM.ROMDATA.dintern_0_2_NEW_1\
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__27448\,
            I => \DROM.ROMDATA.dintern_0_2_NEW_1\
        );

    \I__2816\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27440\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__27440\,
            I => \N__27437\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__27437\,
            I => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_1\
        );

    \I__2813\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27430\
        );

    \I__2812\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27427\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27424\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__27427\,
            I => \N__27421\
        );

    \I__2809\ : Span4Mux_h
    port map (
            O => \N__27424\,
            I => \N__27418\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__27421\,
            I => \N__27415\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__27418\,
            I => \DROM.ROMDATA.dintern_0_2_NEW_2\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__27415\,
            I => \DROM.ROMDATA.dintern_0_2_NEW_2\
        );

    \I__2805\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__27407\,
            I => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_2\
        );

    \I__2803\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__27401\,
            I => \N__27397\
        );

    \I__2801\ : InMux
    port map (
            O => \N__27400\,
            I => \N__27394\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__27397\,
            I => \N__27391\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__27394\,
            I => \N__27388\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__27391\,
            I => \DROM.ROMDATA.dintern_0_2_NEW_3\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__27388\,
            I => \DROM.ROMDATA.dintern_0_2_NEW_3\
        );

    \I__2796\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27380\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__27380\,
            I => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_3\
        );

    \I__2794\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27373\
        );

    \I__2793\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27370\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__27373\,
            I => \N__27367\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__27370\,
            I => \N__27364\
        );

    \I__2790\ : Span12Mux_v
    port map (
            O => \N__27367\,
            I => \N__27361\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__27364\,
            I => \N__27358\
        );

    \I__2788\ : Odrv12
    port map (
            O => \N__27361\,
            I => \DROM.ROMDATA.dintern_0_3_NEW_0\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__27358\,
            I => \DROM.ROMDATA.dintern_0_3_NEW_0\
        );

    \I__2786\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__27350\,
            I => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_0\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__27347\,
            I => \N__27342\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__27346\,
            I => \N__27339\
        );

    \I__2782\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27334\
        );

    \I__2781\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27334\
        );

    \I__2780\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27331\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__27334\,
            I => \N__27328\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__27331\,
            I => \N__27325\
        );

    \I__2777\ : Span4Mux_h
    port map (
            O => \N__27328\,
            I => \N__27322\
        );

    \I__2776\ : Span4Mux_v
    port map (
            O => \N__27325\,
            I => \N__27317\
        );

    \I__2775\ : Span4Mux_v
    port map (
            O => \N__27322\,
            I => \N__27317\
        );

    \I__2774\ : Odrv4
    port map (
            O => \N__27317\,
            I => \DROM_ROMDATA_dintern_6ro\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__27314\,
            I => \CONTROL.N_199_cascade_\
        );

    \I__2772\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27308\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27305\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__27305\,
            I => \N__27302\
        );

    \I__2769\ : Sp12to4
    port map (
            O => \N__27302\,
            I => \N__27299\
        );

    \I__2768\ : Span12Mux_v
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__2767\ : Odrv12
    port map (
            O => \N__27296\,
            I => \gpuOut_c_6\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__27293\,
            I => \DROM_ROMDATA_dintern_13ro_cascade_\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__27290\,
            I => \N__27287\
        );

    \I__2764\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27278\
        );

    \I__2763\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27278\
        );

    \I__2762\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27271\
        );

    \I__2761\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27271\
        );

    \I__2760\ : InMux
    port map (
            O => \N__27283\,
            I => \N__27271\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__27278\,
            I => \N__27265\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__27271\,
            I => \N__27262\
        );

    \I__2757\ : InMux
    port map (
            O => \N__27270\,
            I => \N__27255\
        );

    \I__2756\ : InMux
    port map (
            O => \N__27269\,
            I => \N__27255\
        );

    \I__2755\ : InMux
    port map (
            O => \N__27268\,
            I => \N__27255\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__27265\,
            I => \CONTROL.bus_7_a0_2_8\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__27262\,
            I => \CONTROL.bus_7_a0_2_8\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__27255\,
            I => \CONTROL.bus_7_a0_2_8\
        );

    \I__2751\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27245\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__27245\,
            I => \DROM_ROMDATA_dintern_13ro\
        );

    \I__2749\ : IoInMux
    port map (
            O => \N__27242\,
            I => \N__27239\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__2747\ : IoSpan4Mux
    port map (
            O => \N__27236\,
            I => \N__27232\
        );

    \I__2746\ : IoInMux
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__2745\ : Span4Mux_s0_h
    port map (
            O => \N__27232\,
            I => \N__27226\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27223\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__27226\,
            I => \N__27220\
        );

    \I__2742\ : IoSpan4Mux
    port map (
            O => \N__27223\,
            I => \N__27217\
        );

    \I__2741\ : Span4Mux_h
    port map (
            O => \N__27220\,
            I => \N__27214\
        );

    \I__2740\ : IoSpan4Mux
    port map (
            O => \N__27217\,
            I => \N__27211\
        );

    \I__2739\ : Sp12to4
    port map (
            O => \N__27214\,
            I => \N__27208\
        );

    \I__2738\ : Span4Mux_s2_h
    port map (
            O => \N__27211\,
            I => \N__27205\
        );

    \I__2737\ : Span12Mux_h
    port map (
            O => \N__27208\,
            I => \N__27202\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__27205\,
            I => \N__27199\
        );

    \I__2735\ : Odrv12
    port map (
            O => \N__27202\,
            I => bus_13
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__27199\,
            I => bus_13
        );

    \I__2733\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27190\
        );

    \I__2732\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27187\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__27190\,
            I => \N__27184\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__27187\,
            I => \DROM_ROMDATA_dintern_10ro\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__27184\,
            I => \DROM_ROMDATA_dintern_10ro\
        );

    \I__2728\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27175\
        );

    \I__2727\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27172\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__27175\,
            I => \N__27169\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__27172\,
            I => \N__27166\
        );

    \I__2724\ : Span4Mux_h
    port map (
            O => \N__27169\,
            I => \N__27163\
        );

    \I__2723\ : Span4Mux_h
    port map (
            O => \N__27166\,
            I => \N__27160\
        );

    \I__2722\ : Odrv4
    port map (
            O => \N__27163\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_1\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__27160\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_1\
        );

    \I__2720\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27152\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__27152\,
            I => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_1\
        );

    \I__2718\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27146\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__27146\,
            I => \N__27142\
        );

    \I__2716\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27139\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__27142\,
            I => \N__27136\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__27139\,
            I => \N__27133\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__27136\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_2\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__27133\,
            I => \DROM.ROMDATA.dintern_0_1_NEW_2\
        );

    \I__2711\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27125\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__27125\,
            I => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_2\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__27122\,
            I => \DROM.ROMDATA.dintern_adfltZ0Z_3_cascade_\
        );

    \I__2708\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__27116\,
            I => \DROM.ROMDATA.dintern_adflt_sxZ0\
        );

    \I__2706\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27104\
        );

    \I__2705\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27104\
        );

    \I__2704\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27104\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__27104\,
            I => \dataRomAddress_13\
        );

    \I__2702\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27092\
        );

    \I__2701\ : InMux
    port map (
            O => \N__27100\,
            I => \N__27092\
        );

    \I__2700\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27092\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__27092\,
            I => \dataRomAddress_14\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__27089\,
            I => \N__27084\
        );

    \I__2697\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27077\
        );

    \I__2696\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27077\
        );

    \I__2695\ : InMux
    port map (
            O => \N__27084\,
            I => \N__27077\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__27077\,
            I => \dataRomAddress_15\
        );

    \I__2693\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27071\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__27071\,
            I => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_1\
        );

    \I__2691\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27064\
        );

    \I__2690\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27061\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__27064\,
            I => \N__27058\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__27061\,
            I => \N__27055\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__27058\,
            I => \N__27050\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__27055\,
            I => \N__27050\
        );

    \I__2685\ : Span4Mux_v
    port map (
            O => \N__27050\,
            I => \N__27047\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__27047\,
            I => \DROM.ROMDATA.dintern_0_3_NEW_1\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__27044\,
            I => \N__27041\
        );

    \I__2682\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27035\
        );

    \I__2680\ : Sp12to4
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__2679\ : Odrv12
    port map (
            O => \N__27032\,
            I => \ALU.status_18_cry_3_c_RNOZ0\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__27029\,
            I => \N_228_0_cascade_\
        );

    \I__2677\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__27023\,
            I => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_3\
        );

    \I__2675\ : InMux
    port map (
            O => \N__27020\,
            I => \N__27014\
        );

    \I__2674\ : InMux
    port map (
            O => \N__27019\,
            I => \N__27014\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__27014\,
            I => \N__27011\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__27011\,
            I => \DROM.ROMDATA.dintern_0_0_NEW_3\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__27008\,
            I => \DROM_ROMDATA_dintern_3ro_cascade_\
        );

    \I__2670\ : InMux
    port map (
            O => \N__27005\,
            I => \N__27002\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__27002\,
            I => \DROM_ROMDATA_dintern_1ro\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__26999\,
            I => \DROM_ROMDATA_dintern_adflt_cascade_\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__26996\,
            I => \N__26993\
        );

    \I__2666\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26990\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26987\
        );

    \I__2664\ : Span4Mux_v
    port map (
            O => \N__26987\,
            I => \N__26984\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__26984\,
            I => \DROM.ROMDATA.dintern_adfltZ0Z_3\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__26981\,
            I => \ALU.operand2_10_cascade_\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__26978\,
            I => \ALU.status_19_9_cascade_\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__26975\,
            I => \ALU.e_RNIBHMNZ0Z_8_cascade_\
        );

    \I__2659\ : InMux
    port map (
            O => \N__26972\,
            I => \N__26969\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__26969\,
            I => \ALU.d_RNIIINJZ0Z_8\
        );

    \I__2657\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26963\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__26963\,
            I => \ALU.operand2_7_ns_1_8\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__26960\,
            I => \ALU.b_RNIE6BVZ0Z_8_cascade_\
        );

    \I__2654\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26954\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26951\
        );

    \I__2652\ : Odrv12
    port map (
            O => \N__26951\,
            I => \ALU.operand2_8\
        );

    \I__2651\ : InMux
    port map (
            O => \N__26948\,
            I => \N__26945\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__26945\,
            I => \busState_1_RNI05PC2_0\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__26942\,
            I => \ALU.operand2_8_cascade_\
        );

    \I__2648\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26936\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__26936\,
            I => \N_182\
        );

    \I__2646\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26927\
        );

    \I__2645\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26927\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__26927\,
            I => \N__26924\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__26924\,
            I => \ALU.combOperand2_0_0_6\
        );

    \I__2642\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26918\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__26918\,
            I => \ALU.b_RNI4VJC1Z0Z_12\
        );

    \I__2640\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26912\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__26912\,
            I => \ALU.d_RNI4BCTZ0Z_10\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__26909\,
            I => \ALU.b_RNI0RJC1Z0Z_10_cascade_\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__26906\,
            I => \N__26902\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__26905\,
            I => \N__26899\
        );

    \I__2635\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26896\
        );

    \I__2634\ : InMux
    port map (
            O => \N__26899\,
            I => \N__26892\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__26896\,
            I => \N__26889\
        );

    \I__2632\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26886\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__26892\,
            I => \N__26883\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__26889\,
            I => \ALU.operand2_10\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__26886\,
            I => \ALU.operand2_10\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__26883\,
            I => \ALU.operand2_10\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__26876\,
            I => \ALU.combOperand2_0_4_cascade_\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__26873\,
            I => \N_181_cascade_\
        );

    \I__2625\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26867\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__26867\,
            I => \ALU.d_RNIVKK66Z0Z_4\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__26864\,
            I => \ALU.d_RNIVKK66Z0Z_4_cascade_\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__26861\,
            I => \N__26858\
        );

    \I__2621\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26854\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__26857\,
            I => \N__26851\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__26854\,
            I => \N__26848\
        );

    \I__2618\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26845\
        );

    \I__2617\ : Span4Mux_h
    port map (
            O => \N__26848\,
            I => \N__26841\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__26845\,
            I => \N__26838\
        );

    \I__2615\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26835\
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__26841\,
            I => \ALU.combOperand2_0_4\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__26838\,
            I => \ALU.combOperand2_0_4\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__26835\,
            I => \ALU.combOperand2_0_4\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__26828\,
            I => \N__26825\
        );

    \I__2610\ : InMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__26822\,
            I => \N__26819\
        );

    \I__2608\ : Sp12to4
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__2607\ : Odrv12
    port map (
            O => \N__26816\,
            I => \ALU.status_17_I_33_c_RNOZ0\
        );

    \I__2606\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26809\
        );

    \I__2605\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26806\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__26809\,
            I => \ALU.combOperand2_0_6\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__26806\,
            I => \ALU.combOperand2_0_6\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__26801\,
            I => \ALU.combOperand2_0_6_cascade_\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__26798\,
            I => \ALU.status_19_5_cascade_\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__26795\,
            I => \ALU.dout_6_ns_1_5_cascade_\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__26792\,
            I => \ALU.N_1138_cascade_\
        );

    \I__2598\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26786\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__26786\,
            I => \ALU.N_1090\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__26783\,
            I => \aluOut_5_cascade_\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__26780\,
            I => \ALU.status_19_4_cascade_\
        );

    \I__2594\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__26771\,
            I => \ALU.status_17_I_15_c_RNOZ0\
        );

    \I__2591\ : InMux
    port map (
            O => \N__26768\,
            I => \CONTROL.addrstack_1_cry_0\
        );

    \I__2590\ : InMux
    port map (
            O => \N__26765\,
            I => \CONTROL.addrstack_1_cry_1\
        );

    \I__2589\ : InMux
    port map (
            O => \N__26762\,
            I => \CONTROL.addrstack_1_cry_2\
        );

    \I__2588\ : InMux
    port map (
            O => \N__26759\,
            I => \CONTROL.addrstack_1_cry_3\
        );

    \I__2587\ : InMux
    port map (
            O => \N__26756\,
            I => \CONTROL.addrstack_1_cry_4\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__26753\,
            I => \N__26747\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__26752\,
            I => \N__26744\
        );

    \I__2584\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26737\
        );

    \I__2583\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26737\
        );

    \I__2582\ : InMux
    port map (
            O => \N__26747\,
            I => \N__26737\
        );

    \I__2581\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26734\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__26737\,
            I => \N__26729\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__26734\,
            I => \N__26729\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__26729\,
            I => \CONTROL.addrstackptrZ0Z_6\
        );

    \I__2577\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26719\
        );

    \I__2576\ : InMux
    port map (
            O => \N__26725\,
            I => \N__26719\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__26724\,
            I => \N__26716\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26713\
        );

    \I__2573\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26710\
        );

    \I__2572\ : Odrv12
    port map (
            O => \N__26713\,
            I => \CONTROL.addrstack_1_6\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__26710\,
            I => \CONTROL.addrstack_1_6\
        );

    \I__2570\ : InMux
    port map (
            O => \N__26705\,
            I => \CONTROL.addrstack_1_cry_5\
        );

    \I__2569\ : InMux
    port map (
            O => \N__26702\,
            I => \CONTROL.addrstack_1_cry_6\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__26699\,
            I => \ALU.dout_3_ns_1_5_cascade_\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__26696\,
            I => \CONTROL.g0_3_cascade_\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__26693\,
            I => \CONTROL.addrstackptr_N_10_mux_0_0_0_cascade_\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__26690\,
            I => \N__26687\
        );

    \I__2564\ : InMux
    port map (
            O => \N__26687\,
            I => \N__26684\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__26684\,
            I => \N__26681\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__26681\,
            I => \N__26678\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__26678\,
            I => \CONTROL.addrstackptr_N_7_0_i\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__26675\,
            I => \CONTROL.N_6_1_cascade_\
        );

    \I__2559\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26669\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__26669\,
            I => \CONTROL.N_4_2\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__26666\,
            I => \CONTROL.N_4_2_cascade_\
        );

    \I__2556\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26660\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__26660\,
            I => \CONTROL.addrstackptr_N_10_mux_0_0_0\
        );

    \I__2554\ : InMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__26654\,
            I => \CONTROL.tempCounterZ0Z_13\
        );

    \I__2552\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__26648\,
            I => \N__26645\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__26645\,
            I => \CONTROL.tempCounterZ0Z_6\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__26642\,
            I => \PROM_ROMDATA_dintern_23ro_cascade_\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__26639\,
            I => \N__26636\
        );

    \I__2547\ : CascadeBuf
    port map (
            O => \N__26636\,
            I => \N__26633\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__26633\,
            I => \N__26630\
        );

    \I__2545\ : CascadeBuf
    port map (
            O => \N__26630\,
            I => \N__26627\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__2543\ : CascadeBuf
    port map (
            O => \N__26624\,
            I => \N__26621\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__26621\,
            I => \N__26618\
        );

    \I__2541\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26615\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__26615\,
            I => \N__26612\
        );

    \I__2539\ : Span4Mux_h
    port map (
            O => \N__26612\,
            I => \N__26609\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__26609\,
            I => \CONTROL_romAddReg_7_7\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__2536\ : CascadeBuf
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__26600\,
            I => \N__26597\
        );

    \I__2534\ : CascadeBuf
    port map (
            O => \N__26597\,
            I => \N__26594\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__26594\,
            I => \N__26591\
        );

    \I__2532\ : CascadeBuf
    port map (
            O => \N__26591\,
            I => \N__26588\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__26588\,
            I => \N__26585\
        );

    \I__2530\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__26582\,
            I => \N__26579\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__26579\,
            I => \CONTROL_romAddReg_7_6\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__26576\,
            I => \PROM.ROMDATA.m465_bm_cascade_\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__26573\,
            I => \PROM.ROMDATA.m471_ns_1_cascade_\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__26570\,
            I => \PROM.ROMDATA.m471_ns_cascade_\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__26567\,
            I => \controlWord_24_cascade_\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__26564\,
            I => \N__26561\
        );

    \I__2522\ : CascadeBuf
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__26558\,
            I => \N__26555\
        );

    \I__2520\ : CascadeBuf
    port map (
            O => \N__26555\,
            I => \N__26552\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__26552\,
            I => \N__26549\
        );

    \I__2518\ : CascadeBuf
    port map (
            O => \N__26549\,
            I => \N__26546\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__26546\,
            I => \N__26543\
        );

    \I__2516\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26540\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__26540\,
            I => \CONTROL_romAddReg_7_8\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__26537\,
            I => \N__26534\
        );

    \I__2513\ : CascadeBuf
    port map (
            O => \N__26534\,
            I => \N__26531\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__26531\,
            I => \N__26528\
        );

    \I__2511\ : CascadeBuf
    port map (
            O => \N__26528\,
            I => \N__26525\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__26525\,
            I => \N__26522\
        );

    \I__2509\ : CascadeBuf
    port map (
            O => \N__26522\,
            I => \N__26519\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__26519\,
            I => \N__26516\
        );

    \I__2507\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26513\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__26513\,
            I => \CONTROL_romAddReg_7_4\
        );

    \I__2505\ : IoInMux
    port map (
            O => \N__26510\,
            I => \N__26507\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__26507\,
            I => \N__26504\
        );

    \I__2503\ : Span4Mux_s1_h
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__26501\,
            I => \N__26498\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__26495\,
            I => \gpuAddress_10\
        );

    \I__2499\ : IoInMux
    port map (
            O => \N__26492\,
            I => \N__26489\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__26489\,
            I => \N__26486\
        );

    \I__2497\ : IoSpan4Mux
    port map (
            O => \N__26486\,
            I => \N__26483\
        );

    \I__2496\ : IoSpan4Mux
    port map (
            O => \N__26483\,
            I => \N__26480\
        );

    \I__2495\ : Sp12to4
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__2494\ : Odrv12
    port map (
            O => \N__26477\,
            I => \gpuAddress_12\
        );

    \I__2493\ : IoInMux
    port map (
            O => \N__26474\,
            I => \N__26471\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__26471\,
            I => \N__26468\
        );

    \I__2491\ : IoSpan4Mux
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__2490\ : IoSpan4Mux
    port map (
            O => \N__26465\,
            I => \N__26462\
        );

    \I__2489\ : Span4Mux_s1_h
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__2488\ : Span4Mux_h
    port map (
            O => \N__26459\,
            I => \N__26456\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__26456\,
            I => \gpuAddress_13\
        );

    \I__2486\ : IoInMux
    port map (
            O => \N__26453\,
            I => \N__26450\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__26450\,
            I => \N__26447\
        );

    \I__2484\ : IoSpan4Mux
    port map (
            O => \N__26447\,
            I => \N__26444\
        );

    \I__2483\ : IoSpan4Mux
    port map (
            O => \N__26444\,
            I => \N__26441\
        );

    \I__2482\ : Span4Mux_s2_h
    port map (
            O => \N__26441\,
            I => \N__26438\
        );

    \I__2481\ : Span4Mux_h
    port map (
            O => \N__26438\,
            I => \N__26435\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__26435\,
            I => \gpuAddress_15\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__26432\,
            I => \N__26429\
        );

    \I__2478\ : CascadeBuf
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__2476\ : CascadeBuf
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__2474\ : CascadeBuf
    port map (
            O => \N__26417\,
            I => \N__26414\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__26414\,
            I => \N__26411\
        );

    \I__2472\ : InMux
    port map (
            O => \N__26411\,
            I => \N__26408\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__26408\,
            I => \N__26405\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__26402\,
            I => \CONTROL_romAddReg_7_2\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__26399\,
            I => \N__26396\
        );

    \I__2467\ : CascadeBuf
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__2465\ : CascadeBuf
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__2463\ : CascadeBuf
    port map (
            O => \N__26384\,
            I => \N__26381\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__26381\,
            I => \N__26378\
        );

    \I__2461\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__26372\,
            I => \CONTROL_romAddReg_7_3\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__2457\ : CascadeBuf
    port map (
            O => \N__26366\,
            I => \N__26363\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__2455\ : CascadeBuf
    port map (
            O => \N__26360\,
            I => \N__26357\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__2453\ : CascadeBuf
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__2451\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26345\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__26345\,
            I => \N__26342\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__26339\,
            I => \CONTROL_romAddReg_7_5\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \DROM_ROMDATA_dintern_12ro_cascade_\
        );

    \I__2446\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26330\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__26330\,
            I => \DROM_ROMDATA_dintern_12ro\
        );

    \I__2444\ : IoInMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__2442\ : Span4Mux_s3_h
    port map (
            O => \N__26321\,
            I => \N__26317\
        );

    \I__2441\ : IoInMux
    port map (
            O => \N__26320\,
            I => \N__26314\
        );

    \I__2440\ : Span4Mux_v
    port map (
            O => \N__26317\,
            I => \N__26311\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__26314\,
            I => \N__26308\
        );

    \I__2438\ : Sp12to4
    port map (
            O => \N__26311\,
            I => \N__26305\
        );

    \I__2437\ : Span4Mux_s3_h
    port map (
            O => \N__26308\,
            I => \N__26302\
        );

    \I__2436\ : Span12Mux_s11_h
    port map (
            O => \N__26305\,
            I => \N__26299\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__26302\,
            I => \N__26296\
        );

    \I__2434\ : Span12Mux_h
    port map (
            O => \N__26299\,
            I => \N__26293\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__26296\,
            I => \N__26290\
        );

    \I__2432\ : Span12Mux_v
    port map (
            O => \N__26293\,
            I => \N__26287\
        );

    \I__2431\ : Span4Mux_v
    port map (
            O => \N__26290\,
            I => \N__26284\
        );

    \I__2430\ : Odrv12
    port map (
            O => \N__26287\,
            I => bus_12
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__26284\,
            I => bus_12
        );

    \I__2428\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__26276\,
            I => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_2\
        );

    \I__2426\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26266\
        );

    \I__2424\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26263\
        );

    \I__2423\ : Span4Mux_h
    port map (
            O => \N__26266\,
            I => \N__26258\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__26263\,
            I => \N__26258\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__26255\,
            I => \DROM.ROMDATA.dintern_0_3_NEW_2\
        );

    \I__2419\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26249\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__26249\,
            I => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_3\
        );

    \I__2417\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26242\
        );

    \I__2416\ : InMux
    port map (
            O => \N__26245\,
            I => \N__26239\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__26242\,
            I => \N__26234\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__26239\,
            I => \N__26234\
        );

    \I__2413\ : Span4Mux_v
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__26231\,
            I => \DROM.ROMDATA.dintern_0_3_NEW_3\
        );

    \I__2411\ : IoInMux
    port map (
            O => \N__26228\,
            I => \N__26225\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26221\
        );

    \I__2409\ : IoInMux
    port map (
            O => \N__26224\,
            I => \N__26218\
        );

    \I__2408\ : IoSpan4Mux
    port map (
            O => \N__26221\,
            I => \N__26215\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__26218\,
            I => \N__26212\
        );

    \I__2406\ : Span4Mux_s2_h
    port map (
            O => \N__26215\,
            I => \N__26209\
        );

    \I__2405\ : IoSpan4Mux
    port map (
            O => \N__26212\,
            I => \N__26206\
        );

    \I__2404\ : Sp12to4
    port map (
            O => \N__26209\,
            I => \N__26203\
        );

    \I__2403\ : Span4Mux_s0_h
    port map (
            O => \N__26206\,
            I => \N__26200\
        );

    \I__2402\ : Span12Mux_s10_h
    port map (
            O => \N__26203\,
            I => \N__26197\
        );

    \I__2401\ : Span4Mux_h
    port map (
            O => \N__26200\,
            I => \N__26194\
        );

    \I__2400\ : Span12Mux_h
    port map (
            O => \N__26197\,
            I => \N__26191\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__26194\,
            I => \N__26188\
        );

    \I__2398\ : Span12Mux_v
    port map (
            O => \N__26191\,
            I => \N__26185\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__26188\,
            I => \N__26182\
        );

    \I__2396\ : Odrv12
    port map (
            O => \N__26185\,
            I => bus_10
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__26182\,
            I => bus_10
        );

    \I__2394\ : IoInMux
    port map (
            O => \N__26177\,
            I => \N__26174\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__26174\,
            I => \N__26171\
        );

    \I__2392\ : Span4Mux_s0_h
    port map (
            O => \N__26171\,
            I => \N__26168\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__26168\,
            I => \N__26165\
        );

    \I__2390\ : Span4Mux_h
    port map (
            O => \N__26165\,
            I => \N__26162\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__26162\,
            I => \gpuAddress_0\
        );

    \I__2388\ : IoInMux
    port map (
            O => \N__26159\,
            I => \N__26156\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__26156\,
            I => \N__26153\
        );

    \I__2386\ : Span12Mux_s8_h
    port map (
            O => \N__26153\,
            I => \N__26150\
        );

    \I__2385\ : Odrv12
    port map (
            O => \N__26150\,
            I => \gpuAddress_1\
        );

    \I__2384\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__2383\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26141\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__26141\,
            I => \DROM_ROMDATA_dintern_8ro\
        );

    \I__2381\ : IoInMux
    port map (
            O => \N__26138\,
            I => \N__26135\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26132\
        );

    \I__2379\ : Span12Mux_s8_h
    port map (
            O => \N__26132\,
            I => \N__26128\
        );

    \I__2378\ : IoInMux
    port map (
            O => \N__26131\,
            I => \N__26125\
        );

    \I__2377\ : Span12Mux_v
    port map (
            O => \N__26128\,
            I => \N__26122\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__26125\,
            I => \N__26119\
        );

    \I__2375\ : Span12Mux_h
    port map (
            O => \N__26122\,
            I => \N__26116\
        );

    \I__2374\ : Span12Mux_s8_h
    port map (
            O => \N__26119\,
            I => \N__26113\
        );

    \I__2373\ : Odrv12
    port map (
            O => \N__26116\,
            I => bus_8
        );

    \I__2372\ : Odrv12
    port map (
            O => \N__26113\,
            I => bus_8
        );

    \I__2371\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26102\
        );

    \I__2370\ : InMux
    port map (
            O => \N__26107\,
            I => \N__26102\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__26102\,
            I => \DROM.ROMDATA.dintern_0_0_NEW_1\
        );

    \I__2368\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26096\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__26096\,
            I => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_1\
        );

    \I__2366\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26089\
        );

    \I__2365\ : InMux
    port map (
            O => \N__26092\,
            I => \N__26086\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__26089\,
            I => \N__26081\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__26086\,
            I => \N__26081\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__26081\,
            I => \N__26078\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__26078\,
            I => \DROM.ROMDATA.dintern_0_2_NEW_0\
        );

    \I__2360\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26072\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__26072\,
            I => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_0\
        );

    \I__2358\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26066\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__26066\,
            I => \ALU.log_1_3cf0_1_10\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__26063\,
            I => \ALU.log_1_3cf0_10_cascade_\
        );

    \I__2355\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26057\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__26057\,
            I => \ALU.log_1_3cf1_10\
        );

    \I__2353\ : InMux
    port map (
            O => \N__26054\,
            I => \N__26051\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__26051\,
            I => \ALU.log_1_3cf1_1_10\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__26048\,
            I => \CONTROL.bus_7_a0_2_8_cascade_\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__2349\ : InMux
    port map (
            O => \N__26042\,
            I => \N__26039\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__26039\,
            I => \N__26036\
        );

    \I__2347\ : Odrv12
    port map (
            O => \N__26036\,
            I => \ALU.status_18_cry_8_c_RNOZ0\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \DROM_ROMDATA_dintern_8ro_cascade_\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__26030\,
            I => \ALU.operand2_12_cascade_\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__26027\,
            I => \ALU.N_126_cascade_\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__26024\,
            I => \ALU.c_RNI670LZ0Z_12_cascade_\
        );

    \I__2342\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26018\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__26018\,
            I => \ALU.operand2_7_ns_1_12\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__26015\,
            I => \N__26012\
        );

    \I__2339\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__26009\,
            I => \ALU.d_RNI8FCTZ0Z_12\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__26006\,
            I => \N__26003\
        );

    \I__2336\ : InMux
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__26000\,
            I => \ALU.operand2_12\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__25997\,
            I => \N__25994\
        );

    \I__2333\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25991\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__25985\,
            I => \ALU.status_18_cry_12_c_RNOZ0\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__2328\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__25976\,
            I => \ALU.status_18_cry_10_c_RNOZ0\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__25973\,
            I => \N__25970\
        );

    \I__2325\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__25967\,
            I => \ALU.status_18_cry_13_c_RNOZ0\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__25964\,
            I => \CONTROL.busState_1_RNIG7366Z0Z_2_cascade_\
        );

    \I__2322\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__25958\,
            I => \CONTROL.busState_1_RNI1JVK1_0Z0Z_2\
        );

    \I__2320\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25952\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__2318\ : Span4Mux_v
    port map (
            O => \N__25949\,
            I => \N__25946\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__25946\,
            I => \N__25943\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__2315\ : Span4Mux_v
    port map (
            O => \N__25940\,
            I => \N__25937\
        );

    \I__2314\ : IoSpan4Mux
    port map (
            O => \N__25937\,
            I => \N__25934\
        );

    \I__2313\ : IoSpan4Mux
    port map (
            O => \N__25934\,
            I => \N__25931\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__25931\,
            I => \gpuOut_c_5\
        );

    \I__2311\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25925\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__25925\,
            I => \CONTROL.N_166\
        );

    \I__2309\ : CascadeMux
    port map (
            O => \N__25922\,
            I => \N__25918\
        );

    \I__2308\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25915\
        );

    \I__2307\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25912\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__25915\,
            I => \N__25909\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__25912\,
            I => \N__25906\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__25909\,
            I => \N__25901\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__25906\,
            I => \N__25901\
        );

    \I__2302\ : Sp12to4
    port map (
            O => \N__25901\,
            I => \N__25898\
        );

    \I__2301\ : Span12Mux_h
    port map (
            O => \N__25898\,
            I => \N__25895\
        );

    \I__2300\ : Span12Mux_v
    port map (
            O => \N__25895\,
            I => \N__25892\
        );

    \I__2299\ : Odrv12
    port map (
            O => \N__25892\,
            I => \D5_in_c\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__25889\,
            I => \CONTROL.N_166_cascade_\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__25886\,
            I => \N__25883\
        );

    \I__2296\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25880\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__25880\,
            I => \romOut_5\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__2293\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25871\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__25871\,
            I => \ALU.combOperand2_i_11\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__25868\,
            I => \N__25865\
        );

    \I__2290\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__25862\,
            I => \ALU.combOperand2_i_14\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__25859\,
            I => \N__25856\
        );

    \I__2287\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25853\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__25853\,
            I => \ALU.combOperand2_i_15\
        );

    \I__2285\ : InMux
    port map (
            O => \N__25850\,
            I => \bfn_9_13_0_\
        );

    \I__2284\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__25844\,
            I => \ALU.status_17_I_45_c_RNOZ0\
        );

    \I__2282\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__25838\,
            I => \ALU.combOperand2_i_1\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__2279\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__25826\,
            I => \ALU.status_17_I_27_c_RNOZ0\
        );

    \I__2276\ : InMux
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__25820\,
            I => \ALU.combOperand2_i_7\
        );

    \I__2274\ : InMux
    port map (
            O => \N__25817\,
            I => \bfn_9_10_0_\
        );

    \I__2273\ : InMux
    port map (
            O => \N__25814\,
            I => clkdiv_cry_22
        );

    \I__2272\ : IoInMux
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__2270\ : Span12Mux_s6_v
    port map (
            O => \N__25805\,
            I => \N__25801\
        );

    \I__2269\ : InMux
    port map (
            O => \N__25804\,
            I => \N__25798\
        );

    \I__2268\ : Odrv12
    port map (
            O => \N__25801\,
            I => \GPIO3_c\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__25798\,
            I => \GPIO3_c\
        );

    \I__2266\ : IoInMux
    port map (
            O => \N__25793\,
            I => \N__25788\
        );

    \I__2265\ : IoInMux
    port map (
            O => \N__25792\,
            I => \N__25785\
        );

    \I__2264\ : IoInMux
    port map (
            O => \N__25791\,
            I => \N__25782\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__25788\,
            I => \B_OE_c_i\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__25785\,
            I => \B_OE_c_i\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__25782\,
            I => \B_OE_c_i\
        );

    \I__2260\ : IoInMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__25772\,
            I => \N__25769\
        );

    \I__2258\ : Span4Mux_s2_h
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__2257\ : Sp12to4
    port map (
            O => \N__25766\,
            I => \N__25762\
        );

    \I__2256\ : InMux
    port map (
            O => \N__25765\,
            I => \N__25759\
        );

    \I__2255\ : Span12Mux_s11_v
    port map (
            O => \N__25762\,
            I => \N__25756\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__25759\,
            I => \N__25753\
        );

    \I__2253\ : Odrv12
    port map (
            O => \N__25756\,
            I => \B_OE_c\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__25753\,
            I => \B_OE_c\
        );

    \I__2251\ : IoInMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__25745\,
            I => \N__25742\
        );

    \I__2249\ : Span4Mux_s3_h
    port map (
            O => \N__25742\,
            I => \N__25739\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__25739\,
            I => \N__25736\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__25736\,
            I => \gpuAddress_11\
        );

    \I__2246\ : IoInMux
    port map (
            O => \N__25733\,
            I => \N__25730\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__25730\,
            I => \N__25727\
        );

    \I__2244\ : Span4Mux_s2_h
    port map (
            O => \N__25727\,
            I => \N__25724\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__25724\,
            I => \N__25721\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__25721\,
            I => \N__25718\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__25718\,
            I => \gpuAddress_14\
        );

    \I__2240\ : IoInMux
    port map (
            O => \N__25715\,
            I => \N__25712\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__25712\,
            I => \N__25709\
        );

    \I__2238\ : Span12Mux_s6_h
    port map (
            O => \N__25709\,
            I => \N__25706\
        );

    \I__2237\ : Odrv12
    port map (
            O => \N__25706\,
            I => \gpuAddress_9\
        );

    \I__2236\ : IoInMux
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__25700\,
            I => \N__25697\
        );

    \I__2234\ : IoSpan4Mux
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__2233\ : Span4Mux_s3_h
    port map (
            O => \N__25694\,
            I => \N__25691\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__25691\,
            I => \N_6_0\
        );

    \I__2231\ : IoInMux
    port map (
            O => \N__25688\,
            I => \N__25685\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__25685\,
            I => \N__25681\
        );

    \I__2229\ : IoInMux
    port map (
            O => \N__25684\,
            I => \N__25678\
        );

    \I__2228\ : IoSpan4Mux
    port map (
            O => \N__25681\,
            I => \N__25673\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__25678\,
            I => \N__25673\
        );

    \I__2226\ : Span4Mux_s2_h
    port map (
            O => \N__25673\,
            I => \N__25669\
        );

    \I__2225\ : IoInMux
    port map (
            O => \N__25672\,
            I => \N__25666\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__25669\,
            I => \N__25663\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__25666\,
            I => \N__25660\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__25663\,
            I => \RAM_un1_WR_i\
        );

    \I__2221\ : Odrv12
    port map (
            O => \N__25660\,
            I => \RAM_un1_WR_i\
        );

    \I__2220\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25652\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__25652\,
            I => \clkdivZ0Z_15\
        );

    \I__2218\ : InMux
    port map (
            O => \N__25649\,
            I => clkdiv_cry_14
        );

    \I__2217\ : InMux
    port map (
            O => \N__25646\,
            I => \N__25643\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__25643\,
            I => \clkdivZ0Z_16\
        );

    \I__2215\ : InMux
    port map (
            O => \N__25640\,
            I => \bfn_1_19_0_\
        );

    \I__2214\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25634\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__25634\,
            I => \clkdivZ0Z_17\
        );

    \I__2212\ : InMux
    port map (
            O => \N__25631\,
            I => clkdiv_cry_16
        );

    \I__2211\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25625\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__25625\,
            I => \clkdivZ0Z_18\
        );

    \I__2209\ : InMux
    port map (
            O => \N__25622\,
            I => clkdiv_cry_17
        );

    \I__2208\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25616\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__25616\,
            I => \clkdivZ0Z_19\
        );

    \I__2206\ : InMux
    port map (
            O => \N__25613\,
            I => clkdiv_cry_18
        );

    \I__2205\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25607\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__25607\,
            I => \clkdivZ0Z_20\
        );

    \I__2203\ : InMux
    port map (
            O => \N__25604\,
            I => clkdiv_cry_19
        );

    \I__2202\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25598\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__25598\,
            I => \clkdivZ0Z_21\
        );

    \I__2200\ : InMux
    port map (
            O => \N__25595\,
            I => clkdiv_cry_20
        );

    \I__2199\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__25589\,
            I => \clkdivZ0Z_22\
        );

    \I__2197\ : InMux
    port map (
            O => \N__25586\,
            I => clkdiv_cry_21
        );

    \I__2196\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25580\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__25580\,
            I => \clkdivZ0Z_7\
        );

    \I__2194\ : InMux
    port map (
            O => \N__25577\,
            I => clkdiv_cry_6
        );

    \I__2193\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25571\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__25571\,
            I => \clkdivZ0Z_8\
        );

    \I__2191\ : InMux
    port map (
            O => \N__25568\,
            I => \bfn_1_18_0_\
        );

    \I__2190\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__25562\,
            I => \clkdivZ0Z_9\
        );

    \I__2188\ : InMux
    port map (
            O => \N__25559\,
            I => clkdiv_cry_8
        );

    \I__2187\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__25553\,
            I => \clkdivZ0Z_10\
        );

    \I__2185\ : InMux
    port map (
            O => \N__25550\,
            I => clkdiv_cry_9
        );

    \I__2184\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25544\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__25544\,
            I => \clkdivZ0Z_11\
        );

    \I__2182\ : InMux
    port map (
            O => \N__25541\,
            I => clkdiv_cry_10
        );

    \I__2181\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__25535\,
            I => \clkdivZ0Z_12\
        );

    \I__2179\ : InMux
    port map (
            O => \N__25532\,
            I => clkdiv_cry_11
        );

    \I__2178\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__25526\,
            I => \clkdivZ0Z_13\
        );

    \I__2176\ : InMux
    port map (
            O => \N__25523\,
            I => clkdiv_cry_12
        );

    \I__2175\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__25517\,
            I => \clkdivZ0Z_14\
        );

    \I__2173\ : InMux
    port map (
            O => \N__25514\,
            I => clkdiv_cry_13
        );

    \I__2172\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25508\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__25508\,
            I => \clkdivZ0Z_0\
        );

    \I__2170\ : InMux
    port map (
            O => \N__25505\,
            I => \bfn_1_17_0_\
        );

    \I__2169\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25499\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__25499\,
            I => \clkdivZ0Z_1\
        );

    \I__2167\ : InMux
    port map (
            O => \N__25496\,
            I => clkdiv_cry_0
        );

    \I__2166\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25490\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__25490\,
            I => \clkdivZ0Z_2\
        );

    \I__2164\ : InMux
    port map (
            O => \N__25487\,
            I => clkdiv_cry_1
        );

    \I__2163\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25481\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__25481\,
            I => \clkdivZ0Z_3\
        );

    \I__2161\ : InMux
    port map (
            O => \N__25478\,
            I => clkdiv_cry_2
        );

    \I__2160\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25472\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__25472\,
            I => \clkdivZ0Z_4\
        );

    \I__2158\ : InMux
    port map (
            O => \N__25469\,
            I => clkdiv_cry_3
        );

    \I__2157\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__25463\,
            I => \clkdivZ0Z_5\
        );

    \I__2155\ : InMux
    port map (
            O => \N__25460\,
            I => clkdiv_cry_4
        );

    \I__2154\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25454\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__25454\,
            I => \clkdivZ0Z_6\
        );

    \I__2152\ : InMux
    port map (
            O => \N__25451\,
            I => clkdiv_cry_5
        );

    \INVCONTROL.ramAddReg_6C\ : INV
    port map (
            O => \INVCONTROL.ramAddReg_6C_net\,
            I => \N__73250\
        );

    \INVCONTROL.results_2C\ : INV
    port map (
            O => \INVCONTROL.results_2C_net\,
            I => \N__73249\
        );

    \INVCONTROL.results_1C\ : INV
    port map (
            O => \INVCONTROL.results_1C_net\,
            I => \N__73238\
        );

    \INVCONTROL.increment_1C\ : INV
    port map (
            O => \INVCONTROL.increment_1C_net\,
            I => \N__73207\
        );

    \INVCONTROL.aluOperation_6C\ : INV
    port map (
            O => \INVCONTROL.aluOperation_6C_net\,
            I => \N__73216\
        );

    \INVCONTROL.ramAddReg_3C\ : INV
    port map (
            O => \INVCONTROL.ramAddReg_3C_net\,
            I => \N__73206\
        );

    \INVCONTROL.dout_13C\ : INV
    port map (
            O => \INVCONTROL.dout_13C_net\,
            I => \N__73198\
        );

    \INVCONTROL.increment_0C\ : INV
    port map (
            O => \INVCONTROL.increment_0C_net\,
            I => \N__73245\
        );

    \INVCONTROL.dout_9C\ : INV
    port map (
            O => \INVCONTROL.dout_9C_net\,
            I => \N__73191\
        );

    \INVCONTROL.operand2_fast_ne_1C\ : INV
    port map (
            O => \INVCONTROL.operand2_fast_ne_1C_net\,
            I => \N__73182\
        );

    \INVCONTROL.operand2_2_rep1_neC\ : INV
    port map (
            O => \INVCONTROL.operand2_2_rep1_neC_net\,
            I => \N__73171\
        );

    \INVCONTROL.addrstackptr_2C\ : INV
    port map (
            O => \INVCONTROL.addrstackptr_2C_net\,
            I => \N__73215\
        );

    \INVCONTROL.aluOperation_ne_5C\ : INV
    port map (
            O => \INVCONTROL.aluOperation_ne_5C_net\,
            I => \N__73197\
        );

    \INVCONTROL.dout_2C\ : INV
    port map (
            O => \INVCONTROL.dout_2C_net\,
            I => \N__73201\
        );

    \INVCONTROL.aluOperation_4C\ : INV
    port map (
            O => \INVCONTROL.aluOperation_4C_net\,
            I => \N__73195\
        );

    \INVCONTROL.aluParams_1_ne_1C\ : INV
    port map (
            O => \INVCONTROL.aluParams_1_ne_1C_net\,
            I => \N__73189\
        );

    \INVCONTROL.aluParams_1_0C\ : INV
    port map (
            O => \INVCONTROL.aluParams_1_0C_net\,
            I => \N__73178\
        );

    \INVCONTROL.operand1_ne_0C\ : INV
    port map (
            O => \INVCONTROL.operand1_ne_0C_net\,
            I => \N__73167\
        );

    \INVCONTROL.operand2_fast_ne_2C\ : INV
    port map (
            O => \INVCONTROL.operand2_fast_ne_2C_net\,
            I => \N__73152\
        );

    \INVCONTROL.ramWriteC\ : INV
    port map (
            O => \INVCONTROL.ramWriteC_net\,
            I => \N__73223\
        );

    \INVCONTROL.aluOperation_ne_1C\ : INV
    port map (
            O => \INVCONTROL.aluOperation_ne_1C_net\,
            I => \N__73214\
        );

    \INVCONTROL.addrstackptr_3C\ : INV
    port map (
            O => \INVCONTROL.addrstackptr_3C_net\,
            I => \N__73205\
        );

    \INVCONTROL.operand1_fast_ne_1C\ : INV
    port map (
            O => \INVCONTROL.operand1_fast_ne_1C_net\,
            I => \N__73170\
        );

    \INVCONTROL.tempCounter_4C\ : INV
    port map (
            O => \INVCONTROL.tempCounter_4C_net\,
            I => \N__73255\
        );

    \INVCONTROL.tempCounter_0C\ : INV
    port map (
            O => \INVCONTROL.tempCounter_0C_net\,
            I => \N__73244\
        );

    \INVCONTROL.dout_1C\ : INV
    port map (
            O => \INVCONTROL.dout_1C_net\,
            I => \N__73222\
        );

    \INVCONTROL.busState_1_1C\ : INV
    port map (
            O => \INVCONTROL.busState_1_1C_net\,
            I => \N__73213\
        );

    \INVCONTROL.busState_1_2C\ : INV
    port map (
            O => \INVCONTROL.busState_1_2C_net\,
            I => \N__73204\
        );

    \INVCONTROL.operand1_ne_1C\ : INV
    port map (
            O => \INVCONTROL.operand1_ne_1C_net\,
            I => \N__73180\
        );

    \INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C_net\,
            I => \N__73149\
        );

    \INVCONTROL.ramAddReg_14C\ : INV
    port map (
            O => \INVCONTROL.ramAddReg_14C_net\,
            I => \N__73272\
        );

    \INVCONTROL.addrstackptr_1C\ : INV
    port map (
            O => \INVCONTROL.addrstackptr_1C_net\,
            I => \N__73254\
        );

    \INVCONTROL.ramAddReg_0C\ : INV
    port map (
            O => \INVCONTROL.ramAddReg_0C_net\,
            I => \N__73243\
        );

    \INVCONTROL.dout_15C\ : INV
    port map (
            O => \INVCONTROL.dout_15C_net\,
            I => \N__73231\
        );

    \INVCONTROL.dout_10C\ : INV
    port map (
            O => \INVCONTROL.dout_10C_net\,
            I => \N__73221\
        );

    \INVCONTROL.aluReadBusC\ : INV
    port map (
            O => \INVCONTROL.aluReadBusC_net\,
            I => \N__73203\
        );

    \INVCONTROL.dout_11C\ : INV
    port map (
            O => \INVCONTROL.dout_11C_net\,
            I => \N__73196\
        );

    \INVCONTROL.dout_14C\ : INV
    port map (
            O => \INVCONTROL.dout_14C_net\,
            I => \N__73179\
        );

    \INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C_net\,
            I => \N__73169\
        );

    \INVCONTROL.addrstackptr_4C\ : INV
    port map (
            O => \INVCONTROL.addrstackptr_4C_net\,
            I => \N__73242\
        );

    \INVCONTROL.ramAddReg_5C\ : INV
    port map (
            O => \INVCONTROL.ramAddReg_5C_net\,
            I => \N__73230\
        );

    \INVCONTROL.gpuWriteC\ : INV
    port map (
            O => \INVCONTROL.gpuWriteC_net\,
            I => \N__73220\
        );

    \INVCONTROL.gpuAddReg_2C\ : INV
    port map (
            O => \INVCONTROL.gpuAddReg_2C_net\,
            I => \N__73212\
        );

    \INVCONTROL.dout_7C\ : INV
    port map (
            O => \INVCONTROL.dout_7C_net\,
            I => \N__73202\
        );

    \INVCONTROL.addrstackptr_0C\ : INV
    port map (
            O => \INVCONTROL.addrstackptr_0C_net\,
            I => \N__73139\
        );

    \INVCONTROL.tempCounter_10C\ : INV
    port map (
            O => \INVCONTROL.tempCounter_10C_net\,
            I => \N__73276\
        );

    \INVCONTROL.ramAddReg_13C\ : INV
    port map (
            O => \INVCONTROL.ramAddReg_13C_net\,
            I => \N__73229\
        );

    \INVCONTROL.busState_1_0C\ : INV
    port map (
            O => \INVCONTROL.busState_1_0C_net\,
            I => \N__73219\
        );

    \INVCONTROL.romAddReg_10C\ : INV
    port map (
            O => \INVCONTROL.romAddReg_10C_net\,
            I => \N__73211\
        );

    \INVCONTROL.tempCounter_11C\ : INV
    port map (
            O => \INVCONTROL.tempCounter_11C_net\,
            I => \N__73275\
        );

    \INVCONTROL.addrstackptr_5C\ : INV
    port map (
            O => \INVCONTROL.addrstackptr_5C_net\,
            I => \N__73262\
        );

    \INVCONTROL.dout_6C\ : INV
    port map (
            O => \INVCONTROL.dout_6C_net\,
            I => \N__73252\
        );

    \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            I => \N__73241\
        );

    \INVCONTROL.aluOperation_ne_0C\ : INV
    port map (
            O => \INVCONTROL.aluOperation_ne_0C_net\,
            I => \N__73228\
        );

    \INVCONTROL.romAddReg_13C\ : INV
    port map (
            O => \INVCONTROL.romAddReg_13C_net\,
            I => \N__73218\
        );

    \INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C_net\,
            I => \N__73210\
        );

    \INVCONTROL.tempCounter_13C\ : INV
    port map (
            O => \INVCONTROL.tempCounter_13C_net\,
            I => \N__73282\
        );

    \INVCONTROL.addrstackptr_6C\ : INV
    port map (
            O => \INVCONTROL.addrstackptr_6C_net\,
            I => \N__73277\
        );

    \INVCONTROL.dout_3C\ : INV
    port map (
            O => \INVCONTROL.dout_3C_net\,
            I => \N__73268\
        );

    \INVCONTROL.gpuAddReg_0C\ : INV
    port map (
            O => \INVCONTROL.gpuAddReg_0C_net\,
            I => \N__73261\
        );

    \INVCONTROL.aluOperation_3C\ : INV
    port map (
            O => \INVCONTROL.aluOperation_3C_net\,
            I => \N__73251\
        );

    \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net\,
            I => \N__73240\
        );

    \INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C_net\,
            I => \N__73227\
        );

    \INVCONTROL.dout_5C\ : INV
    port map (
            O => \INVCONTROL.dout_5C_net\,
            I => \N__73200\
        );

    \INVCONTROL.gpuAddReg_9C\ : INV
    port map (
            O => \INVCONTROL.gpuAddReg_9C_net\,
            I => \N__73273\
        );

    \INVCONTROL.gpuAddReg_14C\ : INV
    port map (
            O => \INVCONTROL.gpuAddReg_14C_net\,
            I => \N__73259\
        );

    \INVCONTROL.gpuAddReg_11C\ : INV
    port map (
            O => \INVCONTROL.gpuAddReg_11C_net\,
            I => \N__73280\
        );

    \INVDROM.ROMDATA.dintern_0_0RCLKN\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_0RCLKN_net\,
            I => \N__73239\
        );

    \INVDROM.ROMDATA.dintern_0_1RCLKN\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_1RCLKN_net\,
            I => \N__73260\
        );

    \INVDROM.ROMDATA.dintern_0_2RCLKN\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_2RCLKN_net\,
            I => \N__73274\
        );

    \INVDROM.ROMDATA.dintern_0_3RCLKN\ : INV
    port map (
            O => \INVDROM.ROMDATA.dintern_0_3RCLKN_net\,
            I => \N__73281\
        );

    \INVCONTROL.addrstack_addrstack_0_0RCLKN\ : INV
    port map (
            O => \INVCONTROL.addrstack_addrstack_0_0RCLKN_net\,
            I => \N__73291\
        );

    \IN_MUX_bfv_23_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_14_0_\
        );

    \IN_MUX_bfv_23_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.addsub_cry_6\,
            carryinitout => \bfn_23_15_0_\
        );

    \IN_MUX_bfv_23_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.addsub_cry_14\,
            carryinitout => \bfn_23_16_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \CONTROL.programCounter_1_cry_7\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.status_18_cry_7\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.status_18_4\,
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.status_17_data_tmp_7\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.mult_3_c10\,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.mult_1_c8\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_20_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_10_0_\
        );

    \IN_MUX_bfv_19_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_10_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.mult_7_c14\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.mult_5_c12\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_7,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clkdiv_cry_15,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_23_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_7_0_\
        );

    \IN_MUX_bfv_23_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.status_19_cry_7\,
            carryinitout => \bfn_23_8_0_\
        );

    \IN_MUX_bfv_23_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.status_19Z0Z_5\,
            carryinitout => \bfn_23_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.mult_17_c9\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.mult_25_c11\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_19_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_9_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU.mult_19_c13\,
            carryinitout => \bfn_15_10_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \clkdiv_0_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25511\,
            in2 => \_gnd_net_\,
            in3 => \N__25505\,
            lcout => \clkdivZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => clkdiv_cry_0,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_1_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25502\,
            in2 => \_gnd_net_\,
            in3 => \N__25496\,
            lcout => \clkdivZ0Z_1\,
            ltout => OPEN,
            carryin => clkdiv_cry_0,
            carryout => clkdiv_cry_1,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_2_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25493\,
            in2 => \_gnd_net_\,
            in3 => \N__25487\,
            lcout => \clkdivZ0Z_2\,
            ltout => OPEN,
            carryin => clkdiv_cry_1,
            carryout => clkdiv_cry_2,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_3_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25484\,
            in2 => \_gnd_net_\,
            in3 => \N__25478\,
            lcout => \clkdivZ0Z_3\,
            ltout => OPEN,
            carryin => clkdiv_cry_2,
            carryout => clkdiv_cry_3,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_4_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25475\,
            in2 => \_gnd_net_\,
            in3 => \N__25469\,
            lcout => \clkdivZ0Z_4\,
            ltout => OPEN,
            carryin => clkdiv_cry_3,
            carryout => clkdiv_cry_4,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_5_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25466\,
            in2 => \_gnd_net_\,
            in3 => \N__25460\,
            lcout => \clkdivZ0Z_5\,
            ltout => OPEN,
            carryin => clkdiv_cry_4,
            carryout => clkdiv_cry_5,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_6_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25457\,
            in2 => \_gnd_net_\,
            in3 => \N__25451\,
            lcout => \clkdivZ0Z_6\,
            ltout => OPEN,
            carryin => clkdiv_cry_5,
            carryout => clkdiv_cry_6,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_7_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25583\,
            in2 => \_gnd_net_\,
            in3 => \N__25577\,
            lcout => \clkdivZ0Z_7\,
            ltout => OPEN,
            carryin => clkdiv_cry_6,
            carryout => clkdiv_cry_7,
            clk => \N__73286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_8_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25574\,
            in2 => \_gnd_net_\,
            in3 => \N__25568\,
            lcout => \clkdivZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => clkdiv_cry_8,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_9_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25565\,
            in2 => \_gnd_net_\,
            in3 => \N__25559\,
            lcout => \clkdivZ0Z_9\,
            ltout => OPEN,
            carryin => clkdiv_cry_8,
            carryout => clkdiv_cry_9,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_10_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25556\,
            in2 => \_gnd_net_\,
            in3 => \N__25550\,
            lcout => \clkdivZ0Z_10\,
            ltout => OPEN,
            carryin => clkdiv_cry_9,
            carryout => clkdiv_cry_10,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_11_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25547\,
            in2 => \_gnd_net_\,
            in3 => \N__25541\,
            lcout => \clkdivZ0Z_11\,
            ltout => OPEN,
            carryin => clkdiv_cry_10,
            carryout => clkdiv_cry_11,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_12_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25538\,
            in2 => \_gnd_net_\,
            in3 => \N__25532\,
            lcout => \clkdivZ0Z_12\,
            ltout => OPEN,
            carryin => clkdiv_cry_11,
            carryout => clkdiv_cry_12,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_13_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25529\,
            in2 => \_gnd_net_\,
            in3 => \N__25523\,
            lcout => \clkdivZ0Z_13\,
            ltout => OPEN,
            carryin => clkdiv_cry_12,
            carryout => clkdiv_cry_13,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_14_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25520\,
            in2 => \_gnd_net_\,
            in3 => \N__25514\,
            lcout => \clkdivZ0Z_14\,
            ltout => OPEN,
            carryin => clkdiv_cry_13,
            carryout => clkdiv_cry_14,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_15_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25655\,
            in2 => \_gnd_net_\,
            in3 => \N__25649\,
            lcout => \clkdivZ0Z_15\,
            ltout => OPEN,
            carryin => clkdiv_cry_14,
            carryout => clkdiv_cry_15,
            clk => \N__73290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_16_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25646\,
            in2 => \_gnd_net_\,
            in3 => \N__25640\,
            lcout => \clkdivZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => clkdiv_cry_16,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_17_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25637\,
            in2 => \_gnd_net_\,
            in3 => \N__25631\,
            lcout => \clkdivZ0Z_17\,
            ltout => OPEN,
            carryin => clkdiv_cry_16,
            carryout => clkdiv_cry_17,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_18_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25628\,
            in2 => \_gnd_net_\,
            in3 => \N__25622\,
            lcout => \clkdivZ0Z_18\,
            ltout => OPEN,
            carryin => clkdiv_cry_17,
            carryout => clkdiv_cry_18,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_19_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25619\,
            in2 => \_gnd_net_\,
            in3 => \N__25613\,
            lcout => \clkdivZ0Z_19\,
            ltout => OPEN,
            carryin => clkdiv_cry_18,
            carryout => clkdiv_cry_19,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_20_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25610\,
            in2 => \_gnd_net_\,
            in3 => \N__25604\,
            lcout => \clkdivZ0Z_20\,
            ltout => OPEN,
            carryin => clkdiv_cry_19,
            carryout => clkdiv_cry_20,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_21_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25601\,
            in2 => \_gnd_net_\,
            in3 => \N__25595\,
            lcout => \clkdivZ0Z_21\,
            ltout => OPEN,
            carryin => clkdiv_cry_20,
            carryout => clkdiv_cry_21,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_22_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25592\,
            in2 => \_gnd_net_\,
            in3 => \N__25586\,
            lcout => \clkdivZ0Z_22\,
            ltout => OPEN,
            carryin => clkdiv_cry_21,
            carryout => clkdiv_cry_22,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clkdiv_23_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25804\,
            in2 => \_gnd_net_\,
            in3 => \N__25814\,
            lcout => \GPIO3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GPU.BUFFER.B_OE_c_i_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25765\,
            lcout => \B_OE_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GPU.BUFFER.OE_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__29474\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__73304\,
            lcout => \B_OE_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_11_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31234\,
            in1 => \N__70795\,
            in2 => \N__58004\,
            in3 => \N__70552\,
            lcout => \gpuAddress_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_11C_net\,
            ce => \N__30760\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_14_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31411\,
            in1 => \N__70794\,
            in2 => \N__57869\,
            in3 => \N__70548\,
            lcout => \gpuAddress_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_14C_net\,
            ce => \N__30761\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_25dflt_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72376\,
            in2 => \_gnd_net_\,
            in3 => \N__72248\,
            lcout => \controlWord_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_9_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31123\,
            in1 => \N__70761\,
            in2 => \N__37970\,
            in3 => \N__70535\,
            lcout => \gpuAddress_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_9C_net\,
            ce => \N__30752\,
            sr => \_gnd_net_\
        );

    \RAM.OE_i_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__73302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34989\,
            lcout => \N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM.un1_WR_i_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__73303\,
            in1 => \N__34990\,
            in2 => \N__29387\,
            in3 => \N__28148\,
            lcout => \RAM_un1_WR_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_1_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28598\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \ALU.status_17_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_9_c_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32464\,
            in2 => \N__27683\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_17_data_tmp_0\,
            carryout => \ALU.status_17_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_15_c_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26777\,
            in2 => \N__32479\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_17_data_tmp_1\,
            carryout => \ALU.status_17_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_27_c_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32456\,
            in2 => \N__25835\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_17_data_tmp_2\,
            carryout => \ALU.status_17_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_45_c_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25847\,
            in2 => \N__32481\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_17_data_tmp_3\,
            carryout => \ALU.status_17_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_33_c_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32457\,
            in2 => \N__26828\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_17_data_tmp_4\,
            carryout => \ALU.status_17_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_39_c_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37403\,
            in2 => \N__32480\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_17_data_tmp_5\,
            carryout => \ALU.status_17_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_21_c_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53030\,
            in2 => \N__32482\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_17_data_tmp_6\,
            carryout => \ALU.status_17_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_0_3_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69529\,
            in1 => \N__45448\,
            in2 => \N__56627\,
            in3 => \N__25817\,
            lcout => \aluStatus_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_45_c_RNO_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__61935\,
            in1 => \N__62890\,
            in2 => \N__62956\,
            in3 => \N__55817\,
            lcout => \ALU.status_17_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_0_c_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60617\,
            in2 => \N__35324\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \ALU.status_18_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_1_c_inv_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25841\,
            in2 => \N__65574\,
            in3 => \N__66048\,
            lcout => \ALU.combOperand2_i_1\,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_0\,
            carryout => \ALU.status_18_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_2_c_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66313\,
            in2 => \N__32378\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_1\,
            carryout => \ALU.status_18_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_3_c_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60261\,
            in2 => \N__27044\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_2\,
            carryout => \ALU.status_18_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_4_c_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59873\,
            in2 => \N__26861\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_3\,
            carryout => \ALU.status_18_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_5_c_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59503\,
            in2 => \N__34016\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_4\,
            carryout => \ALU.status_18_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_27_c_RNO_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111101011"
        )
    port map (
            in0 => \N__55993\,
            in1 => \N__26813\,
            in2 => \N__62579\,
            in3 => \N__62186\,
            lcout => \ALU.status_17_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_5\,
            carryout => \ALU.status_18_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_7_c_inv_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25823\,
            in2 => \N__62234\,
            in3 => \N__55992\,
            lcout => \ALU.combOperand2_i_7\,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_6\,
            carryout => \ALU.status_18_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_8_c_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61947\,
            in2 => \N__26045\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \ALU.status_18_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_9_c_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62891\,
            in2 => \N__62957\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_8\,
            carryout => \ALU.status_18_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_10_c_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61681\,
            in2 => \N__25982\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_9\,
            carryout => \ALU.status_18_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_11_c_inv_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61433\,
            in2 => \N__25877\,
            in3 => \N__57031\,
            lcout => \ALU.combOperand2_i_11\,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_10\,
            carryout => \ALU.status_18_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_12_c_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61193\,
            in2 => \N__25997\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_11\,
            carryout => \ALU.status_18_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_13_c_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60995\,
            in2 => \N__25973\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_12\,
            carryout => \ALU.status_18_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_14_c_inv_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63847\,
            in2 => \N__25868\,
            in3 => \N__56753\,
            lcout => \ALU.combOperand2_i_14\,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_13\,
            carryout => \ALU.status_18_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_15_c_inv_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63674\,
            in2 => \N__25859\,
            in3 => \N__74608\,
            lcout => \ALU.combOperand2_i_15\,
            ltout => OPEN,
            carryin => \ALU.status_18_cry_14\,
            carryout => \ALU.status_18_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_4_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69530\,
            in1 => \N__40729\,
            in2 => \N__56623\,
            in3 => \N__25850\,
            lcout => \aluStatus_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_10_c_RNO_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__61682\,
            in1 => \N__71452\,
            in2 => \N__26906\,
            in3 => \N__37120\,
            lcout => \ALU.status_18_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3D2O61_2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__56900\,
            in1 => \N__60246\,
            in2 => \N__56824\,
            in3 => \N__66292\,
            lcout => \ALU.d_RNI3D2O61Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_13_c_RNO_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__39674\,
            in1 => \N__39651\,
            in2 => \N__61013\,
            in3 => \N__71453\,
            lcout => \ALU.status_18_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIG7366_2_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__50225\,
            in1 => \N__59587\,
            in2 => \N__25886\,
            in3 => \N__49596\,
            lcout => OPEN,
            ltout => \CONTROL.busState_1_RNIG7366Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI3G078_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__25961\,
            in1 => \_gnd_net_\,
            in2 => \N__25964\,
            in3 => \N__49829\,
            lcout => bus_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI1JVK1_0_2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__50224\,
            in1 => \N__25928\,
            in2 => \N__25922\,
            in3 => \N__49595\,
            lcout => \CONTROL.busState_1_RNI1JVK1_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI6MOJ_5_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25955\,
            in1 => \N__45673\,
            in2 => \_gnd_net_\,
            in3 => \N__50222\,
            lcout => \CONTROL.N_166\,
            ltout => \CONTROL.N_166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI1JVK1_2_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__50223\,
            in1 => \N__25921\,
            in2 => \N__25889\,
            in3 => \N__49594\,
            lcout => \N_182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI6OIF1_1_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__28920\,
            in1 => \N__27905\,
            in2 => \N__26996\,
            in3 => \N__27962\,
            lcout => \romOut_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_5_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__40912\,
            in1 => \N__50620\,
            in2 => \N__79532\,
            in3 => \N__38801\,
            lcout => \CONTROL.ctrlOut_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_5C_net\,
            ce => \N__44461\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_21dflt_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__79523\,
            in2 => \N__50621\,
            in3 => \N__40911\,
            lcout => \controlWord_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1C0D5_12_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__53967\,
            in1 => \N__26921\,
            in2 => \N__26015\,
            in3 => \N__26021\,
            lcout => \ALU.operand2_12\,
            ltout => \ALU.operand2_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0UD4G_12_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31755\,
            in2 => \N__26030\,
            in3 => \N__71449\,
            lcout => \ALU.N_126\,
            ltout => \ALU.N_126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9UI0K_1_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26027\,
            in3 => \N__65563\,
            lcout => \ALU.d_RNI9UI0KZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8I8I5_0_10_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26895\,
            in2 => \_gnd_net_\,
            in3 => \N__71450\,
            lcout => \ALU.log_1_3cf0_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI670L_12_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52411\,
            in1 => \N__67556\,
            in2 => \_gnd_net_\,
            in3 => \N__43307\,
            lcout => OPEN,
            ltout => \ALU.c_RNI670LZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIHJ2L2_12_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__46841\,
            in1 => \N__53966\,
            in2 => \N__26024\,
            in3 => \N__28952\,
            lcout => \ALU.operand2_7_ns_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8FCT_12_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__57946\,
            in1 => \N__65096\,
            in2 => \_gnd_net_\,
            in3 => \N__43308\,
            lcout => \ALU.d_RNI8FCTZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_12_c_RNO_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__61199\,
            in1 => \N__31756\,
            in2 => \N__26006\,
            in3 => \N__71451\,
            lcout => \ALU.status_18_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIIBVU9_10_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101110010010"
        )
    port map (
            in0 => \N__63247\,
            in1 => \N__26069\,
            in2 => \N__74889\,
            in3 => \N__61662\,
            lcout => OPEN,
            ltout => \ALU.log_1_3cf0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJPU5U_10_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26060\,
            in2 => \N__26063\,
            in3 => \N__37113\,
            lcout => \ALU.log_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIIBVU9_0_10_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111001101000"
        )
    port map (
            in0 => \N__63246\,
            in1 => \N__26054\,
            in2 => \N__74888\,
            in3 => \N__61661\,
            lcout => \ALU.log_1_3cf1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8I8I5_10_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__71424\,
            in1 => \_gnd_net_\,
            in2 => \N__26905\,
            in3 => \_gnd_net_\,
            lcout => \ALU.log_1_3cf1_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIMSAK1_0_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__49587\,
            in1 => \N__50298\,
            in2 => \N__49824\,
            in3 => \N__50190\,
            lcout => \CONTROL.bus_7_a0_2_8\,
            ltout => \CONTROL.bus_7_a0_2_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIF208A_0_0_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27194\,
            in2 => \N__26048\,
            in3 => \N__29056\,
            lcout => bus_0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_8_c_RNO_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__57094\,
            in1 => \N__26957\,
            in2 => \N__61948\,
            in3 => \N__71425\,
            lcout => \ALU.status_18_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIA8EO_0_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32308\,
            in1 => \N__26075\,
            in2 => \_gnd_net_\,
            in3 => \N__26092\,
            lcout => \DROM_ROMDATA_dintern_8ro\,
            ltout => \DROM_ROMDATA_dintern_8ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI05PC2_0_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26033\,
            in3 => \N__27268\,
            lcout => \busState_1_RNI05PC2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIA6749_0_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__27269\,
            in1 => \N__26146\,
            in2 => \_gnd_net_\,
            in3 => \N__29120\,
            lcout => bus_0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIA6749_0_0_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001111"
        )
    port map (
            in0 => \N__27270\,
            in1 => \N__26147\,
            in2 => \N__27842\,
            in3 => \_gnd_net_\,
            lcout => bus_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI7LJL_1_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26099\,
            in1 => \N__26107\,
            in2 => \_gnd_net_\,
            in3 => \N__32307\,
            lcout => \DROM_ROMDATA_dintern_1ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_1_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26108\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_1C_net\,
            ce => \N__32324\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_1_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27068\,
            lcout => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net\,
            ce => \N__32321\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_2_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26273\,
            lcout => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net\,
            ce => \N__32321\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_3_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26246\,
            lcout => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net\,
            ce => \N__32321\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_0_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26093\,
            lcout => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_3_OLD_ne_1C_net\,
            ce => \N__32321\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_RNICIR11_0_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27353\,
            in1 => \N__27376\,
            in2 => \_gnd_net_\,
            in3 => \N__32302\,
            lcout => \DROM_ROMDATA_dintern_12ro\,
            ltout => \DROM_ROMDATA_dintern_12ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI8R4IA_0_0_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30541\,
            in2 => \N__26336\,
            in3 => \N__27283\,
            lcout => bus_0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_3_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__36689\,
            in1 => \N__69766\,
            in2 => \N__38140\,
            in3 => \N__41504\,
            lcout => \aluOperation_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluOperation_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI8R4IA_0_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__26333\,
            in1 => \N__30542\,
            in2 => \_gnd_net_\,
            in3 => \N__27284\,
            lcout => bus_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIDBEO_3_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27383\,
            in1 => \N__27400\,
            in2 => \_gnd_net_\,
            in3 => \N__32300\,
            lcout => \DROM_ROMDATA_dintern_11ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIEKR11_2_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32301\,
            in1 => \N__26279\,
            in2 => \_gnd_net_\,
            in3 => \N__26269\,
            lcout => \DROM_ROMDATA_dintern_14ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIFLR11_3_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26252\,
            in1 => \N__26245\,
            in2 => \_gnd_net_\,
            in3 => \N__32303\,
            lcout => \DROM_ROMDATA_dintern_15ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIF208A_0_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__29057\,
            in1 => \N__27193\,
            in2 => \_gnd_net_\,
            in3 => \N__27285\,
            lcout => bus_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__33317\,
            in1 => \N__70785\,
            in2 => \N__70544\,
            in3 => \N__37565\,
            lcout => \gpuAddress_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_0C_net\,
            ce => \N__30739\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_1_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__70541\,
            in1 => \N__37520\,
            in2 => \N__70798\,
            in3 => \N__33257\,
            lcout => \gpuAddress_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_0C_net\,
            ce => \N__30739\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_10_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31276\,
            in1 => \N__70542\,
            in2 => \N__58241\,
            in3 => \N__70786\,
            lcout => \gpuAddress_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_0C_net\,
            ce => \N__30739\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_12_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__57950\,
            in1 => \N__70543\,
            in2 => \N__28229\,
            in3 => \N__70787\,
            lcout => \gpuAddress_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_0C_net\,
            ce => \N__30739\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_13_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__70539\,
            in1 => \N__27988\,
            in2 => \N__70796\,
            in3 => \N__57908\,
            lcout => \gpuAddress_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_0C_net\,
            ce => \N__30739\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_15_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__70540\,
            in1 => \N__54194\,
            in2 => \N__70797\,
            in3 => \N__45010\,
            lcout => \gpuAddress_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_0C_net\,
            ce => \N__30739\,
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_2_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__29596\,
            in1 => \N__72212\,
            in2 => \N__35570\,
            in3 => \N__71822\,
            lcout => \CONTROL_romAddReg_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_3_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__71825\,
            in1 => \N__37745\,
            in2 => \N__72289\,
            in3 => \N__44278\,
            lcout => \CONTROL_romAddReg_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_3_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__44279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__72220\,
            lcout => \CONTROL.ctrlOut_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_3C_net\,
            ce => \N__44462\,
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_5_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__40148\,
            in1 => \N__72213\,
            in2 => \N__29451\,
            in3 => \N__71823\,
            lcout => \CONTROL_romAddReg_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m461_ns_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100010001"
        )
    port map (
            in0 => \N__47762\,
            in1 => \N__72773\,
            in2 => \N__55505\,
            in3 => \N__74072\,
            lcout => \PROM_ROMDATA_dintern_23ro\,
            ltout => \PROM_ROMDATA_dintern_23ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_7_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__72247\,
            in1 => \N__48872\,
            in2 => \N__26642\,
            in3 => \N__71824\,
            lcout => \CONTROL_romAddReg_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_6_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__71826\,
            in1 => \N__35760\,
            in2 => \N__72288\,
            in3 => \N__70815\,
            lcout => \CONTROL_romAddReg_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m465_bm_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__64022\,
            in1 => \N__76625\,
            in2 => \N__65033\,
            in3 => \N__76015\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m465_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m471_ns_1_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__33416\,
            in1 => \N__79500\,
            in2 => \N__26576\,
            in3 => \N__79896\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m471_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m471_ns_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__79501\,
            in1 => \N__40985\,
            in2 => \N__26573\,
            in3 => \N__29615\,
            lcout => \PROM.ROMDATA.m471_ns\,
            ltout => \PROM.ROMDATA.m471_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_24dflt_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__47494\,
            in1 => \N__72774\,
            in2 => \N__26570\,
            in3 => \N__72221\,
            lcout => \controlWord_24\,
            ltout => \controlWord_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_8_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__71873\,
            in1 => \N__72223\,
            in2 => \N__26567\,
            in3 => \N__50438\,
            lcout => \CONTROL_romAddReg_7_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_4_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__44178\,
            in1 => \N__72222\,
            in2 => \N__35807\,
            in3 => \N__71874\,
            lcout => \CONTROL_romAddReg_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI2UPI1_5_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34769\,
            in1 => \N__57819\,
            in2 => \N__60735\,
            in3 => \N__27499\,
            lcout => OPEN,
            ltout => \CONTROL.g0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI6P3NN91_4_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38443\,
            in1 => \N__60813\,
            in2 => \N__26696\,
            in3 => \N__41986\,
            lcout => \CONTROL.addrstackptr_N_10_mux_0_0_0\,
            ltout => \CONTROL.addrstackptr_N_10_mux_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNIEKK1Q82_6_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__26750\,
            in1 => \N__26725\,
            in2 => \N__26693\,
            in3 => \N__26672\,
            lcout => \CONTROL.addrstackptr_N_7_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_19_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36470\,
            in1 => \N__42261\,
            in2 => \N__45368\,
            in3 => \N__38184\,
            lcout => OPEN,
            ltout => \CONTROL.N_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIDB191V_7_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38516\,
            in1 => \N__42044\,
            in2 => \N__26675\,
            in3 => \N__41503\,
            lcout => \CONTROL.N_4_2\,
            ltout => \CONTROL.N_4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_6_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__26726\,
            in1 => \N__26751\,
            in2 => \N__26666\,
            in3 => \N__26663\,
            lcout => \CONTROL.addrstackptrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.addrstackptr_6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI73QI1_6_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34770\,
            in1 => \N__27498\,
            in2 => \N__26753\,
            in3 => \N__38442\,
            lcout => \CONTROL.g1_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_13_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28343\,
            lcout => \CONTROL.tempCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_13C_net\,
            ce => \N__34970\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_6_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47839\,
            lcout => \CONTROL.tempCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_13C_net\,
            ce => \N__34970\,
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_0_c_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57791\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \CONTROL.addrstack_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_0_c_RNIDDJK_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38431\,
            in2 => \N__32567\,
            in3 => \N__26768\,
            lcout => \CONTROL.addrstack_1_1\,
            ltout => OPEN,
            carryin => \CONTROL.addrstack_1_cry_0\,
            carryout => \CONTROL.addrstack_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_1_c_RNIFGKK_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32554\,
            in2 => \N__60734\,
            in3 => \N__26765\,
            lcout => \CONTROL.addrstack_1_2\,
            ltout => OPEN,
            carryin => \CONTROL.addrstack_1_cry_1\,
            carryout => \CONTROL.addrstack_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_2_c_RNIHJLK_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34768\,
            in2 => \N__32568\,
            in3 => \N__26762\,
            lcout => \CONTROL.addrstack_1_3\,
            ltout => OPEN,
            carryin => \CONTROL.addrstack_1_cry_2\,
            carryout => \CONTROL.addrstack_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_3_c_RNIJMMK_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32558\,
            in2 => \N__60812\,
            in3 => \N__26759\,
            lcout => \CONTROL.addrstack_1_4\,
            ltout => OPEN,
            carryin => \CONTROL.addrstack_1_cry_3\,
            carryout => \CONTROL.addrstack_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_4_c_RNILPNK_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27500\,
            in2 => \N__32569\,
            in3 => \N__26756\,
            lcout => \CONTROL.addrstack_1_5\,
            ltout => OPEN,
            carryin => \CONTROL.addrstack_1_cry_4\,
            carryout => \CONTROL.addrstack_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_5_c_RNINSOK_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32562\,
            in2 => \N__26752\,
            in3 => \N__26705\,
            lcout => \CONTROL.addrstack_1_6\,
            ltout => OPEN,
            carryin => \CONTROL.addrstack_1_cry_5\,
            carryout => \CONTROL.addrstack_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_1_cry_6_c_RNIPVPK_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42287\,
            in2 => \_gnd_net_\,
            in3 => \N__26702\,
            lcout => \CONTROL.addrstack_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI69B31_5_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__40036\,
            in1 => \N__34568\,
            in2 => \N__40070\,
            in3 => \N__43931\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIE8D02_5_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__40144\,
            in1 => \N__40097\,
            in2 => \N__26699\,
            in3 => \N__47212\,
            lcout => \ALU.N_1090\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI8FH51_5_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__39932\,
            in1 => \N__34567\,
            in2 => \N__39972\,
            in3 => \N__43930\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIKPK1_5_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__40239\,
            in1 => \N__40220\,
            in2 => \N__26795\,
            in3 => \N__47213\,
            lcout => OPEN,
            ltout => \ALU.N_1138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI31LU3_5_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54143\,
            in2 => \N__26792\,
            in3 => \N__26789\,
            lcout => \aluOut_5\,
            ltout => \aluOut_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJRM75_5_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__53289\,
            in1 => \N__49607\,
            in2 => \N__26783\,
            in3 => \N__50220\,
            lcout => \ALU.d_RNIJRM75Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILKJ1I_5_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__59486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56077\,
            lcout => \ALU.d_RNILKJ1IZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIK31N31_10_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__61427\,
            in1 => \N__56377\,
            in2 => \N__68517\,
            in3 => \N__61667\,
            lcout => \ALU.c_RNIK31N31Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7BDMH_7_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62185\,
            in2 => \_gnd_net_\,
            in3 => \N__56078\,
            lcout => \ALU.d_RNI7BDMHZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILEAFE_5_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__40585\,
            in1 => \N__28933\,
            in2 => \N__28921\,
            in3 => \N__28876\,
            lcout => \ALU.status_19_4\,
            ltout => \ALU.status_19_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI07V431_2_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__56378\,
            in1 => \N__60245\,
            in2 => \N__26780\,
            in3 => \N__66296\,
            lcout => \ALU.d_RNI07V431Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_15_c_RNO_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101111010111"
        )
    port map (
            in0 => \N__34012\,
            in1 => \N__59881\,
            in2 => \N__26857\,
            in3 => \N__59487\,
            lcout => \ALU.status_17_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIUEFBI_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65558\,
            in2 => \_gnd_net_\,
            in3 => \N__56196\,
            lcout => \ALU.d_RNIUEFBIZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIALE3I_6_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__26812\,
            in1 => \_gnd_net_\,
            in2 => \N__63292\,
            in3 => \N__62506\,
            lcout => \ALU.d_RNIALE3IZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIJU2E_0_6_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__26933\,
            in1 => \N__27345\,
            in2 => \N__32693\,
            in3 => \N__40581\,
            lcout => \ALU.combOperand2_0_6\,
            ltout => \ALU.combOperand2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA9P4I_6_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001110000110"
        )
    port map (
            in0 => \N__63265\,
            in1 => \N__74890\,
            in2 => \N__26801\,
            in3 => \N__62505\,
            lcout => \ALU.N_22_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI67HQ21_0_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__65545\,
            in1 => \N__60593\,
            in2 => \N__68506\,
            in3 => \N__56328\,
            lcout => \ALU.d_RNI67HQ21Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIJU2E_6_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111111"
        )
    port map (
            in0 => \N__40580\,
            in1 => \N__32689\,
            in2 => \N__27347\,
            in3 => \N__26932\,
            lcout => \ALU.status_19_5\,
            ltout => \ALU.status_19_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5NE641_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__65544\,
            in1 => \N__60594\,
            in2 => \N__26798\,
            in3 => \N__56223\,
            lcout => \ALU.d_RNI5NE641Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBLU321_6_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__55989\,
            in1 => \N__62504\,
            in2 => \N__62324\,
            in3 => \N__55801\,
            lcout => \ALU.d_RNIBLU321Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI73D441_6_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__62503\,
            in1 => \N__56076\,
            in2 => \N__62316\,
            in3 => \N__56224\,
            lcout => \ALU.d_RNI73D441Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVPV6E_0_4_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__27755\,
            in1 => \N__26870\,
            in2 => \N__40592\,
            in3 => \N__28013\,
            lcout => \ALU.combOperand2_0_4\,
            ltout => \ALU.combOperand2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7BF7I_4_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \N__59802\,
            in1 => \_gnd_net_\,
            in2 => \N__26876\,
            in3 => \N__63260\,
            lcout => \ALU.d_RNI7BF7IZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un14_log_a0_2_15_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__50216\,
            in1 => \N__53232\,
            in2 => \N__49606\,
            in3 => \N__50327\,
            lcout => \ALU.un14_log_a0_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIU83C1_2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__37994\,
            in1 => \N__49600\,
            in2 => \N__33143\,
            in3 => \N__50217\,
            lcout => OPEN,
            ltout => \N_181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVKK66_4_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__53233\,
            in1 => \N__71440\,
            in2 => \N__26873\,
            in3 => \N__27797\,
            lcout => \ALU.d_RNIVKK66Z0Z_4\,
            ltout => \ALU.d_RNIVKK66Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVPV6E_4_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__28012\,
            in1 => \N__40576\,
            in2 => \N__26864\,
            in3 => \N__27754\,
            lcout => \ALU.status_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7VP8I_4_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101110010010"
        )
    port map (
            in0 => \N__63261\,
            in1 => \N__26844\,
            in2 => \N__74903\,
            in3 => \N__59801\,
            lcout => \ALU.log_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8JFO21_6_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__68438\,
            in1 => \N__62502\,
            in2 => \N__62302\,
            in3 => \N__56345\,
            lcout => \ALU.d_RNI8JFO21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_33_c_RNO_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__57033\,
            in1 => \N__61463\,
            in2 => \N__61718\,
            in3 => \N__55549\,
            lcout => \ALU.status_17_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI1QK5K_10_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__55548\,
            in1 => \_gnd_net_\,
            in2 => \N__63293\,
            in3 => \N__61714\,
            lcout => \ALU.c_RNI1QK5KZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIRRB4I_11_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__57032\,
            in1 => \N__63269\,
            in2 => \_gnd_net_\,
            in3 => \N__61464\,
            lcout => \ALU.c_RNIRRB4IZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC0VE6_5_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__71441\,
            in1 => \N__26939\,
            in2 => \N__53291\,
            in3 => \N__40001\,
            lcout => \ALU.d_RNIC0VE6Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI18J1J_3_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60219\,
            in2 => \_gnd_net_\,
            in3 => \N__55547\,
            lcout => \ALU.d_RNI18J1JZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKHEQH_7_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62274\,
            in2 => \_gnd_net_\,
            in3 => \N__56346\,
            lcout => \ALU.d_RNIKHEQHZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMCVI41_2_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__60220\,
            in1 => \N__55546\,
            in2 => \N__55670\,
            in3 => \N__66299\,
            lcout => \ALU.d_RNIMCVI41Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4BCT_10_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__43304\,
            in1 => \_gnd_net_\,
            in2 => \N__36034\,
            in3 => \N__58234\,
            lcout => \ALU.d_RNI4BCTZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0SI26_6_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111111"
        )
    port map (
            in0 => \N__49798\,
            in1 => \N__27572\,
            in2 => \N__71448\,
            in3 => \N__27818\,
            lcout => \ALU.combOperand2_0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI4VJC1_12_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43306\,
            in1 => \N__57685\,
            in2 => \_gnd_net_\,
            in3 => \N__39818\,
            lcout => \ALU.b_RNI4VJC1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI0RJC1_10_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36003\,
            in1 => \N__39137\,
            in2 => \_gnd_net_\,
            in3 => \N__43305\,
            lcout => OPEN,
            ltout => \ALU.b_RNI0RJC1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHRVC5_10_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__26915\,
            in1 => \N__27857\,
            in2 => \N__26909\,
            in3 => \N__53965\,
            lcout => \ALU.operand2_10\,
            ltout => \ALU.operand2_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINK8QF_10_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__71410\,
            in1 => \_gnd_net_\,
            in2 => \N__26981\,
            in3 => \N__37112\,
            lcout => \ALU.status_19_9\,
            ltout => \ALU.status_19_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0LDMJ_1_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26978\,
            in3 => \N__65562\,
            lcout => \ALU.d_RNI0LDMJZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIBHMN_8_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46280\,
            in1 => \N__48745\,
            in2 => \_gnd_net_\,
            in3 => \N__46944\,
            lcout => OPEN,
            ltout => \ALU.e_RNIBHMNZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI34KF2_8_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__27968\,
            in1 => \N__53909\,
            in2 => \N__26975\,
            in3 => \N__46840\,
            lcout => \ALU.operand2_7_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIINJ_8_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48141\,
            in1 => \N__51580\,
            in2 => \_gnd_net_\,
            in3 => \N__43277\,
            lcout => \ALU.d_RNIIINJZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIE6BV_8_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49045\,
            in1 => \N__48326\,
            in2 => \_gnd_net_\,
            in3 => \N__43279\,
            lcout => OPEN,
            ltout => \ALU.b_RNIE6BVZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI77KG4_8_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__26972\,
            in1 => \N__26966\,
            in2 => \N__26960\,
            in3 => \N__53910\,
            lcout => \ALU.operand2_8\,
            ltout => \ALU.operand2_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI844QD_8_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011111100"
        )
    port map (
            in0 => \N__26948\,
            in1 => \N__71423\,
            in2 => \N__26942\,
            in3 => \N__27835\,
            lcout => \ALU.status_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI230L_10_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43278\,
            in1 => \N__35722\,
            in2 => \_gnd_net_\,
            in3 => \N__36136\,
            lcout => \ALU.c_RNI230LZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_3_c_RNO_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__38058\,
            in1 => \N__60218\,
            in2 => \N__33057\,
            in3 => \N__53238\,
            lcout => \ALU.status_18_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIUV6T5_2_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000101"
        )
    port map (
            in0 => \N__28576\,
            in1 => \N__49524\,
            in2 => \N__60247\,
            in3 => \N__50203\,
            lcout => \N_228_0\,
            ltout => \N_228_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHMDUU_3_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010001"
        )
    port map (
            in0 => \N__38057\,
            in1 => \N__53237\,
            in2 => \N__27029\,
            in3 => \N__68939\,
            lcout => \ALU.lshift62_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_3_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_3C_net\,
            ce => \N__32299\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI9NJL_3_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27026\,
            in1 => \N__32295\,
            in2 => \_gnd_net_\,
            in3 => \N__27019\,
            lcout => OPEN,
            ltout => \DROM_ROMDATA_dintern_3ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIDU0U1_2_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__49561\,
            in1 => \N__50280\,
            in2 => \N__27008\,
            in3 => \N__50202\,
            lcout => \busState_1_RNIDU0U1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_adflt_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__27936\,
            in1 => \N__27898\,
            in2 => \_gnd_net_\,
            in3 => \N__27119\,
            lcout => \DROM_ROMDATA_dintern_adflt\,
            ltout => \DROM_ROMDATA_dintern_adflt_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIBS0U1_2_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__27005\,
            in1 => \N__49523\,
            in2 => \N__26999\,
            in3 => \N__50201\,
            lcout => \busState_1_RNIBS0U1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_adflt_3_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27113\,
            in1 => \N__27088\,
            in2 => \N__27938\,
            in3 => \N__27101\,
            lcout => \DROM.ROMDATA.dintern_adfltZ0Z_3\,
            ltout => \DROM.ROMDATA.dintern_adfltZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI5NIF1_0_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__27897\,
            in1 => \N__28003\,
            in2 => \N__27122\,
            in3 => \N__27955\,
            lcout => \romOut_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_RNIDE6K_12_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27954\,
            in1 => \N__27896\,
            in2 => \N__27937\,
            in3 => \N__50127\,
            lcout => \CONTROL.bus_6_a0_sx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_adflt_sx_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27099\,
            in1 => \N__27111\,
            in2 => \N__27089\,
            in3 => \N__27953\,
            lcout => \DROM.ROMDATA.dintern_adflt_sxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_adflt_3_x_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__27112\,
            in1 => \N__27087\,
            in2 => \_gnd_net_\,
            in3 => \N__27100\,
            lcout => dintern_adflt_3_x,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_13_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__27989\,
            in1 => \N__72102\,
            in2 => \N__52357\,
            in3 => \N__71870\,
            lcout => \dataRomAddress_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.romAddReg_13C_net\,
            ce => \N__28111\,
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_14_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__71869\,
            in1 => \N__52304\,
            in2 => \N__31412\,
            in3 => \N__72104\,
            lcout => \dataRomAddress_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.romAddReg_13C_net\,
            ce => \N__28111\,
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_15_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__45009\,
            in1 => \N__72103\,
            in2 => \N__50405\,
            in3 => \N__71871\,
            lcout => \dataRomAddress_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.romAddReg_13C_net\,
            ce => \N__28111\,
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_ne_0_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__41432\,
            in1 => \N__71872\,
            in2 => \_gnd_net_\,
            in3 => \N__54689\,
            lcout => \aluOperation_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluOperation_ne_0C_net\,
            ce => \N__38144\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_RNIDJR11_1_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27074\,
            in1 => \N__27067\,
            in2 => \_gnd_net_\,
            in3 => \N__32264\,
            lcout => \DROM_ROMDATA_dintern_13ro\,
            ltout => \DROM_ROMDATA_dintern_13ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIN5MIA_0_0_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34456\,
            in2 => \N__27293\,
            in3 => \N__27286\,
            lcout => bus_0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIN5MIA_0_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101010101"
        )
    port map (
            in0 => \N__34457\,
            in1 => \_gnd_net_\,
            in2 => \N__27290\,
            in3 => \N__27248\,
            lcout => bus_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_RNICAEO_2_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32263\,
            in1 => \N__27410\,
            in2 => \_gnd_net_\,
            in3 => \N__27433\,
            lcout => \DROM_ROMDATA_dintern_10ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI9V0V_1_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27155\,
            in1 => \N__27178\,
            in2 => \_gnd_net_\,
            in3 => \N__32260\,
            lcout => \DROM_ROMDATA_dintern_5ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIA01V_2_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32261\,
            in1 => \N__27128\,
            in2 => \_gnd_net_\,
            in3 => \N__27145\,
            lcout => \DROM_ROMDATA_dintern_6ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_RNIB9EO_1_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27443\,
            in1 => \N__27466\,
            in2 => \_gnd_net_\,
            in3 => \N__32262\,
            lcout => \DROM_ROMDATA_dintern_9ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_0_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28033\,
            lcout => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_1_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27179\,
            lcout => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_2_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27149\,
            lcout => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_3_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28061\,
            lcout => \DROM.ROMDATA.dintern_0_1_OLDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_1_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27467\,
            lcout => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_2_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27434\,
            lcout => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_2_OLD_ne_3_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27404\,
            lcout => \DROM.ROMDATA.dintern_0_2_OLDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_3_OLD_ne_0_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27377\,
            lcout => \DROM.ROMDATA.dintern_0_3_OLDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_1_OLD_ne_0C_net\,
            ce => \N__32320\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_6_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__40892\,
            in1 => \N__43744\,
            in2 => \N__79531\,
            in3 => \N__71579\,
            lcout => \CONTROL.ctrlOut_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_6C_net\,
            ce => \N__44457\,
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI5P5Q5_1_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__62556\,
            in1 => \N__50324\,
            in2 => \N__27346\,
            in3 => \N__50113\,
            lcout => OPEN,
            ltout => \CONTROL.N_199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIF3TV7_0_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__49786\,
            in1 => \N__27571\,
            in2 => \N__27314\,
            in3 => \N__49553\,
            lcout => bus_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI8OOJ_6_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27311\,
            in1 => \N__45583\,
            in2 => \_gnd_net_\,
            in3 => \N__50111\,
            lcout => OPEN,
            ltout => \CONTROL.N_167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI4TRD1_2_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__50112\,
            in1 => \N__27596\,
            in2 => \N__27575\,
            in3 => \N__49552\,
            lcout => \N_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_22dflt_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__71578\,
            in1 => \N__79514\,
            in2 => \N__43745\,
            in3 => \N__40889\,
            lcout => \controlWord_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_4_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__40891\,
            in1 => \N__65236\,
            in2 => \N__79530\,
            in3 => \N__74213\,
            lcout => \CONTROL.ctrlOut_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_6C_net\,
            ce => \N__44457\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_20dflt_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__74212\,
            in1 => \N__79515\,
            in2 => \N__65237\,
            in3 => \N__40890\,
            lcout => \controlWord_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI37DAN91_3_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34771\,
            in1 => \N__57821\,
            in2 => \N__27659\,
            in3 => \N__41982\,
            lcout => \CONTROL.addrstackptr_N_8_mux_1_0\,
            ltout => \CONTROL.addrstackptr_N_8_mux_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNIAEEIH92_5_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__27493\,
            in1 => \N__27529\,
            in2 => \N__27557\,
            in3 => \N__27536\,
            lcout => \CONTROL.addrstackptr_N_6_0_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIO2O5VB_0_7_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__54681\,
            in1 => \N__41488\,
            in2 => \N__71876\,
            in3 => \N__44696\,
            lcout => OPEN,
            ltout => \CONTROL.g0_3_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIFRI6PV_0_7_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__27665\,
            in1 => \N__38185\,
            in2 => \N__27539\,
            in3 => \N__27671\,
            lcout => \CONTROL.N_4_0\,
            ltout => \CONTROL.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_5_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__27530\,
            in1 => \N__27494\,
            in2 => \N__27509\,
            in3 => \N__27506\,
            lcout => \CONTROL.addrstackptrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.addrstackptr_5C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_1_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101111111"
        )
    port map (
            in0 => \N__42265\,
            in1 => \N__55470\,
            in2 => \N__72284\,
            in3 => \N__54680\,
            lcout => \CONTROL.g0_3_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_a7_2_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__54679\,
            in1 => \N__40676\,
            in2 => \N__63485\,
            in3 => \N__38272\,
            lcout => \CONTROL.g0_3_i_a7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI1E361_4_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__38441\,
            in1 => \_gnd_net_\,
            in2 => \N__60814\,
            in3 => \N__60723\,
            lcout => \CONTROL.g0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_12_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27647\,
            lcout => \CONTROL.addrstack_reto_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_11_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27632\,
            lcout => \CONTROL_addrstack_reto_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_13_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43676\,
            lcout => \CONTROL.dout_reto_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_7_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27620\,
            lcout => \CONTROL.addrstack_reto_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_14_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27608\,
            lcout => \CONTROL.addrstack_reto_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIJDJ31_3_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__73668\,
            in1 => \N__64532\,
            in2 => \_gnd_net_\,
            in3 => \N__64487\,
            lcout => \CONTROL.programCounter_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_11_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29726\,
            lcout => \CONTROL.tempCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_11C_net\,
            ce => \N__34966\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_15_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.tempCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_11C_net\,
            ce => \N__34966\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_14_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29648\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.tempCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_11C_net\,
            ce => \N__34966\,
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_8_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27701\,
            lcout => \CONTROL_addrstack_reto_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_9_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27692\,
            lcout => \CONTROL.addrstack_reto_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHJSI82_4_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__59842\,
            in1 => \N__59585\,
            in2 => \N__28472\,
            in3 => \N__65953\,
            lcout => \ALU.N_860\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFGGBO_0_6_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__62570\,
            in1 => \N__62307\,
            in2 => \_gnd_net_\,
            in3 => \N__66735\,
            lcout => \ALU.N_609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_9_c_RNO_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__68270\,
            in1 => \N__66298\,
            in2 => \N__60262\,
            in3 => \N__68825\,
            lcout => \ALU.status_17_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI0QV651_10_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__56240\,
            in1 => \N__61426\,
            in2 => \N__61668\,
            in3 => \N__56394\,
            lcout => \ALU.c_RNI0QV651Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIOFVDI_5_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59483\,
            in2 => \_gnd_net_\,
            in3 => \N__56239\,
            lcout => \ALU.d_RNIOFVDIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPNF141_4_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__59840\,
            in1 => \N__55681\,
            in2 => \N__55816\,
            in3 => \N__59485\,
            lcout => \ALU.d_RNIPNF141Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI88K161_4_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__59484\,
            in1 => \N__59841\,
            in2 => \N__55688\,
            in3 => \N__55585\,
            lcout => \ALU.d_RNI88K161Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_2_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39479\,
            in1 => \N__39611\,
            in2 => \_gnd_net_\,
            in3 => \N__39539\,
            lcout => h_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73148\,
            ce => \N__69458\,
            sr => \_gnd_net_\
        );

    \ALU.h_4_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57421\,
            in1 => \N__42549\,
            in2 => \_gnd_net_\,
            in3 => \N__39377\,
            lcout => h_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73148\,
            ce => \N__69458\,
            sr => \_gnd_net_\
        );

    \ALU.h_5_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57422\,
            in1 => \N__39319\,
            in2 => \_gnd_net_\,
            in3 => \N__52635\,
            lcout => h_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73148\,
            ce => \N__69458\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNITPMMO_0_6_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__62551\,
            in1 => \N__59479\,
            in2 => \_gnd_net_\,
            in3 => \N__66733\,
            lcout => \ALU.N_608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITPMMO_6_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__66734\,
            in1 => \_gnd_net_\,
            in2 => \N__59540\,
            in3 => \N__62552\,
            lcout => \ALU.N_833\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2RK5I_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59476\,
            in2 => \_gnd_net_\,
            in3 => \N__56360\,
            lcout => \ALU.d_RNI2RK5IZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6HBMG_5_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__59477\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55985\,
            lcout => \ALU.d_RNI6HBMGZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIB5POH_5_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59478\,
            in2 => \_gnd_net_\,
            in3 => \N__55768\,
            lcout => \ALU.d_RNIB5POHZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMQM8I_5_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59549\,
            lcout => \ALU.d_RNIMQM8IZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISSV4I_9_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__56202\,
            in1 => \N__62829\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ALU.d_RNISSV4IZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIK9E841_6_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__56359\,
            in1 => \N__62518\,
            in2 => \N__62315\,
            in3 => \N__56201\,
            lcout => \ALU.d_RNIK9E841Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJ0U031_2_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56068\,
            in1 => \N__60190\,
            in2 => \N__56229\,
            in3 => \N__66297\,
            lcout => \ALU.d_RNIJ0U031Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIV1LMH_3_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56200\,
            lcout => \ALU.d_RNIV1LMHZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9DAEH_3_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60188\,
            in2 => \_gnd_net_\,
            in3 => \N__56357\,
            lcout => \ALU.d_RNI9DAEHZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIITFA41_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__65539\,
            in1 => \N__60589\,
            in2 => \N__56228\,
            in3 => \N__56358\,
            lcout => \ALU.d_RNIITFA41Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISP66I_1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55660\,
            in2 => \_gnd_net_\,
            in3 => \N__65541\,
            lcout => \ALU.d_RNISP66IZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKRBVN_4_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__60192\,
            in1 => \_gnd_net_\,
            in2 => \N__59866\,
            in3 => \N__66662\,
            lcout => \ALU.N_831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKG0L11_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56327\,
            in1 => \N__60196\,
            in2 => \N__68505\,
            in3 => \N__66269\,
            lcout => \ALU.d_RNIKG0L11Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI12A911_2_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__66270\,
            in1 => \N__55959\,
            in2 => \N__60241\,
            in3 => \N__56082\,
            lcout => \ALU.d_RNI12A911Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINIF011_2_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__60227\,
            in1 => \N__55767\,
            in2 => \N__55984\,
            in3 => \N__66271\,
            lcout => \ALU.d_RNINIF011Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJTUN21_4_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__59817\,
            in1 => \N__55960\,
            in2 => \N__56096\,
            in3 => \N__59550\,
            lcout => \ALU.d_RNIJTUN21Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIS69AH_3_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60191\,
            in2 => \_gnd_net_\,
            in3 => \N__56069\,
            lcout => \ALU.d_RNIS69AHZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8Q43I_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__65540\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56326\,
            lcout => \ALU.d_RNI8Q43IZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_3_c_RNIGCKVJ5_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__59672\,
            in1 => \N__66976\,
            in2 => \_gnd_net_\,
            in3 => \N__35282\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_3_c_RNIGCKVJZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_3_c_RNIM4CUT9_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__34178\,
            in1 => \N__48554\,
            in2 => \N__27746\,
            in3 => \N__68431\,
            lcout => \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9\,
            ltout => \ALU.addsub_cry_3_c_RNIM4CUTZ0Z9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_4_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__42550\,
            in1 => \N__57406\,
            in2 => \N__27743\,
            in3 => \_gnd_net_\,
            lcout => \ALU.aZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73168\,
            ce => \N__71212\,
            sr => \_gnd_net_\
        );

    \ALU.e_RNI26JM_4_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__44000\,
            in1 => \_gnd_net_\,
            in2 => \N__32663\,
            in3 => \N__27782\,
            lcout => OPEN,
            ltout => \ALU.e_RNI26JMZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIFKVD2_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__53956\,
            in1 => \N__53435\,
            in2 => \N__27740\,
            in3 => \N__27791\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI19244_4_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__43325\,
            in1 => \N__53957\,
            in2 => \N__27800\,
            in3 => \N__43430\,
            lcout => \ALU.operand2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI6IVQ_4_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35796\,
            in1 => \N__35852\,
            in2 => \_gnd_net_\,
            in3 => \N__43999\,
            lcout => \ALU.c_RNI6IVQZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI6DH51_4_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__43448\,
            in1 => \N__34560\,
            in2 => \N__44155\,
            in3 => \N__43920\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEGPK1_4_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__43348\,
            in1 => \N__43386\,
            in2 => \N__27785\,
            in3 => \N__47203\,
            lcout => \ALU.N_1137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI47B31_4_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__27781\,
            in1 => \N__34561\,
            in2 => \N__32662\,
            in3 => \N__43921\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIA4D02_4_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__35797\,
            in1 => \N__35851\,
            in2 => \N__27770\,
            in3 => \N__47204\,
            lcout => OPEN,
            ltout => \ALU.N_1089_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIROKU3_4_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54138\,
            in2 => \N__27767\,
            in3 => \N__27764\,
            lcout => \aluOut_4\,
            ltout => \aluOut_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBJM75_4_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__53245\,
            in1 => \N__49583\,
            in2 => \N__27758\,
            in3 => \N__50199\,
            lcout => \ALU.d_RNIBJM75Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI990621_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__55994\,
            in1 => \N__65538\,
            in2 => \N__60609\,
            in3 => \N__55724\,
            lcout => \ALU.d_RNI990621Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRU9M31_6_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__62265\,
            in1 => \N__55647\,
            in2 => \N__62572\,
            in3 => \N__55726\,
            lcout => \ALU.d_RNIRU9M31Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIINE1H_3_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60157\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55725\,
            lcout => \ALU.d_RNIINE1HZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKDVI51_4_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__59800\,
            in1 => \N__59595\,
            in2 => \N__57024\,
            in3 => \N__55558\,
            lcout => \ALU.d_RNIKDVI51Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJP1AE_9_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111111"
        )
    port map (
            in0 => \N__40593\,
            in1 => \N__40540\,
            in2 => \N__40494\,
            in3 => \N__40520\,
            lcout => \ALU.status_19_8\,
            ltout => \ALU.status_19_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITCCHH_3_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27824\,
            in3 => \N__60158\,
            lcout => \ALU.d_RNITCCHHZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIPLDD2_6_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__27806\,
            in1 => \N__27878\,
            in2 => \N__53969\,
            in3 => \N__46831\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJIG34_6_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__27872\,
            in1 => \N__27812\,
            in2 => \N__27821\,
            in3 => \N__53961\,
            lcout => \ALU.operand2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI9JSP_6_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39899\,
            in1 => \N__70585\,
            in2 => \_gnd_net_\,
            in3 => \N__46943\,
            lcout => \ALU.b_RNI9JSPZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI6AJM_6_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43998\,
            in1 => \N__32732\,
            in2 => \_gnd_net_\,
            in3 => \N__42937\,
            lcout => \ALU.e_RNI6AJMZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIAMVQ_6_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35768\,
            in1 => \N__35834\,
            in2 => \_gnd_net_\,
            in3 => \N__43997\,
            lcout => \ALU.c_RNIAMVQZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDV8E_6_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46942\,
            in1 => \N__37438\,
            in2 => \_gnd_net_\,
            in3 => \N__36062\,
            lcout => \ALU.d_RNIDV8EZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIUI741_10_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32635\,
            in1 => \N__37076\,
            in2 => \_gnd_net_\,
            in3 => \N__43287\,
            lcout => OPEN,
            ltout => \ALU.a_RNIUI741Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI9B2L2_10_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__46832\,
            in1 => \N__27866\,
            in2 => \N__27860\,
            in3 => \N__53962\,
            lcout => \ALU.operand2_7_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNISTG51_8_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__48325\,
            in1 => \N__32825\,
            in2 => \N__49044\,
            in3 => \N__36341\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBFGH1_8_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__48142\,
            in1 => \N__51587\,
            in2 => \N__27851\,
            in3 => \N__54297\,
            lcout => \ALU_N_1141\,
            ltout => \ALU_N_1141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_RNIEQRR4_0_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__34481\,
            in1 => \N__54141\,
            in2 => \N__27848\,
            in3 => \N__29026\,
            lcout => OPEN,
            ltout => \CONTROL.bus_0_sx_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIA1EN6_0_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49758\,
            in2 => \N__27845\,
            in3 => \N__33166\,
            lcout => \CONTROL_bus_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIQNA31_8_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__48752\,
            in1 => \N__32824\,
            in2 => \N__46279\,
            in3 => \N__36340\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI734T1_8_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__50431\,
            in1 => \N__46378\,
            in2 => \N__27971\,
            in3 => \N__54296\,
            lcout => \ALU_N_1093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFT2S_8_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46379\,
            in1 => \N__50430\,
            in2 => \_gnd_net_\,
            in3 => \N__46946\,
            lcout => \ALU.c_RNIFT2SZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_10_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__31277\,
            in1 => \N__72008\,
            in2 => \N__35723\,
            in3 => \N__71867\,
            lcout => \dataRomAddress_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.romAddReg_10C_net\,
            ce => \N__28110\,
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_12_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__71866\,
            in1 => \N__28228\,
            in2 => \N__72140\,
            in3 => \N__52412\,
            lcout => \dataRomAddress_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.romAddReg_10C_net\,
            ce => \N__28110\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_adflt_4_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28310\,
            in1 => \N__28286\,
            in2 => \N__29747\,
            in3 => \N__28418\,
            lcout => \PROM.ROMDATA.dintern_adfltZ0Z_4\,
            ltout => \PROM.ROMDATA.dintern_adfltZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_adflt_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__28442\,
            in1 => \N__30346\,
            in2 => \N__27917\,
            in3 => \N__28519\,
            lcout => \PROM_ROMDATA_dintern_adflt\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_12dflt_0_1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__30373\,
            in1 => \N__64663\,
            in2 => \N__30407\,
            in3 => \N__28441\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.dintern_12dflt_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_12dflt_0_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__72712\,
            in1 => \N__28520\,
            in2 => \N__27914\,
            in3 => \N__27911\,
            lcout => \PROM.ROMDATA.dintern_12dfltZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_11_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__35678\,
            in1 => \N__72009\,
            in2 => \N__31233\,
            in3 => \N__71868\,
            lcout => \dataRomAddress_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.romAddReg_10C_net\,
            ce => \N__28110\,
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNO_0_0_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010001"
        )
    port map (
            in0 => \N__35141\,
            in1 => \N__35189\,
            in2 => \N__41702\,
            in3 => \N__30794\,
            lcout => OPEN,
            ltout => \CONTROL.busState_1_e_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_0_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100011"
        )
    port map (
            in0 => \N__28079\,
            in1 => \N__40636\,
            in2 => \N__28130\,
            in3 => \N__49742\,
            lcout => \busState_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.busState_1_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState_1_sqmuxa_i_0_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__38713\,
            in1 => \N__31466\,
            in2 => \N__29539\,
            in3 => \N__30793\,
            lcout => \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0\,
            ltout => \CONTROL.un1_busState_1_sqmuxa_iZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState_1_sqmuxa_i_i_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__36621\,
            in1 => \N__38715\,
            in2 => \N__28127\,
            in3 => \N__54750\,
            lcout => \N_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m11_0_a2_1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__38714\,
            in1 => \N__41260\,
            in2 => \N__29540\,
            in3 => \N__41431\,
            lcout => \CONTROL.N_352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_sr_en_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__38716\,
            in1 => \N__54751\,
            in2 => \N__36626\,
            in3 => \N__28073\,
            lcout => \DROM.ROMDATA.dintern_0_0_sr_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.busState_1_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_RNIB11V_3_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28067\,
            in1 => \N__28057\,
            in2 => \_gnd_net_\,
            in3 => \N__32246\,
            lcout => \DROM_ROMDATA_dintern_7ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_1_OLD_ne_RNI8U0V_0_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32247\,
            in1 => \N__28040\,
            in2 => \_gnd_net_\,
            in3 => \N__28034\,
            lcout => \DROM_ROMDATA_dintern_4ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_29dflt_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__76637\,
            in1 => \N__43690\,
            in2 => \N__44324\,
            in3 => \N__43721\,
            lcout => \controlWord_29\,
            ltout => \controlWord_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_13_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__70462\,
            in1 => \N__57621\,
            in2 => \N__28232\,
            in3 => \N__70763\,
            lcout => \A13_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_13C_net\,
            ce => \N__70340\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_28dflt_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__72741\,
            in1 => \N__47477\,
            in2 => \N__65149\,
            in3 => \N__72133\,
            lcout => \controlWord_28\,
            ltout => \controlWord_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_12_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__70461\,
            in1 => \N__57675\,
            in2 => \N__28208\,
            in3 => \N__70762\,
            lcout => \A12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_13C_net\,
            ce => \N__70340\,
            sr => \_gnd_net_\
        );

    \RAM.un1_WR_105_0_10_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__28186\,
            in1 => \N__44021\,
            in2 => \_gnd_net_\,
            in3 => \N__28159\,
            lcout => \RAM.un1_WR_105_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m520_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__79871\,
            in1 => \N__44320\,
            in2 => \N__79529\,
            in3 => \N__76636\,
            lcout => \PROM.ROMDATA.m520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_29dflt_1_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__79522\,
            in1 => \N__79872\,
            in2 => \N__72772\,
            in3 => \N__72132\,
            lcout => \PROM.ROMDATA.dintern_29dfltZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m514_ns_1_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__79870\,
            in1 => \N__76635\,
            in2 => \N__79528\,
            in3 => \N__75985\,
            lcout => \PROM.ROMDATA.m514_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_0_c_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36728\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \CONTROL.programCounter_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_0_c_RNI26EE1_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29789\,
            in2 => \_gnd_net_\,
            in3 => \N__28136\,
            lcout => \CONTROL.programCounter_1_1\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_0\,
            carryout => \CONTROL.programCounter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_1_c_RNIRV7S1_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__78065\,
            in2 => \_gnd_net_\,
            in3 => \N__28133\,
            lcout => \CONTROL.programCounter_1_2\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_1\,
            carryout => \CONTROL.programCounter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_2_c_RNIAGGE1_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28271\,
            in2 => \_gnd_net_\,
            in3 => \N__28259\,
            lcout => \CONTROL.programCounter_1_3\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_2\,
            carryout => \CONTROL.programCounter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_3_c_RNIELHE1_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47330\,
            in2 => \_gnd_net_\,
            in3 => \N__28256\,
            lcout => \CONTROL.programCounter_1_4\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_3\,
            carryout => \CONTROL.programCounter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_4_c_RNI5AT91_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36743\,
            in2 => \_gnd_net_\,
            in3 => \N__28253\,
            lcout => \CONTROL.programCounter_1_5\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_4\,
            carryout => \CONTROL.programCounter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_5_c_RNIOM9I1_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__79486\,
            in2 => \_gnd_net_\,
            in3 => \N__28250\,
            lcout => \CONTROL.programCounter_1_6\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_5\,
            carryout => \CONTROL.programCounter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_6_c_RNIDKV91_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72737\,
            in2 => \_gnd_net_\,
            in3 => \N__28247\,
            lcout => \CONTROL.programCounter_1_7\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_6\,
            carryout => \CONTROL.programCounter_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_7_c_RNIHP0A1_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28376\,
            in2 => \_gnd_net_\,
            in3 => \N__28244\,
            lcout => \CONTROL.programCounter_1_8\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \CONTROL.programCounter_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_8_c_RNI39V71_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28547\,
            in2 => \_gnd_net_\,
            in3 => \N__28241\,
            lcout => \CONTROL.programCounter_1_9\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_8\,
            carryout => \CONTROL.programCounter_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_9_c_RNI67I81_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28440\,
            in2 => \_gnd_net_\,
            in3 => \N__28238\,
            lcout => \CONTROL.programCounter_1_10\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_9\,
            carryout => \CONTROL.programCounter_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_10_c_RNIHFO21_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30350\,
            in2 => \_gnd_net_\,
            in3 => \N__28235\,
            lcout => \CONTROL.programCounter_1_11\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_10\,
            carryout => \CONTROL.programCounter_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_11_c_RNIBCO41_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28417\,
            in2 => \_gnd_net_\,
            in3 => \N__28355\,
            lcout => \CONTROL.programCounter_1_12\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_11\,
            carryout => \CONTROL.programCounter_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_12_c_RNIFHP41_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28309\,
            in2 => \_gnd_net_\,
            in3 => \N__28352\,
            lcout => \CONTROL.programCounter_1_13\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_12\,
            carryout => \CONTROL.programCounter_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_13_c_RNIJMQ41_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28285\,
            in2 => \_gnd_net_\,
            in3 => \N__28349\,
            lcout => \CONTROL.programCounter_1_14\,
            ltout => OPEN,
            carryin => \CONTROL.programCounter_1_cry_13\,
            carryout => \CONTROL.programCounter_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_14_c_RNINRR41_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29740\,
            in2 => \_gnd_net_\,
            in3 => \N__28346\,
            lcout => \CONTROL.programCounter_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_13_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28342\,
            lcout => \CONTROL.programCounter_1_reto_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI3EMQ_13_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28325\,
            in1 => \N__28319\,
            in2 => \_gnd_net_\,
            in3 => \N__42080\,
            lcout => OPEN,
            ltout => \CONTROL.N_428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI7NCV_13_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29822\,
            in2 => \N__28313\,
            in3 => \N__28448\,
            lcout => \progRomAddress_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIAQCV_14_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29823\,
            in1 => \_gnd_net_\,
            in2 => \N__28295\,
            in3 => \N__29510\,
            lcout => \progRomAddress_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_13_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28463\,
            lcout => \CONTROL.addrstack_reto_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI8MDT_10_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28391\,
            in1 => \N__64619\,
            in2 => \_gnd_net_\,
            in3 => \N__29795\,
            lcout => \progRomAddress_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI4KCV_12_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28424\,
            in1 => \N__36701\,
            in2 => \_gnd_net_\,
            in3 => \N__29821\,
            lcout => \progRomAddress_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_10_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28403\,
            lcout => \CONTROL.addrstack_reto_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_8_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33586\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIK8GE_8_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28385\,
            in1 => \N__29504\,
            in2 => \_gnd_net_\,
            in3 => \N__45121\,
            lcout => \N_423\,
            ltout => \N_423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNILCUU_8_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__73687\,
            in2 => \N__28379\,
            in3 => \N__28538\,
            lcout => \CONTROL.programCounter_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_9_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28496\,
            lcout => \CONTROL.programCounter_1_reto_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_addrstack_0_0_RNO_0_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50836\,
            in2 => \_gnd_net_\,
            in3 => \N__50903\,
            lcout => \CONTROL.programCounter10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNID2FG_9_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29753\,
            in1 => \N__28562\,
            in2 => \_gnd_net_\,
            in3 => \N__42086\,
            lcout => OPEN,
            ltout => \CONTROL.N_424_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI6QRS_9_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28556\,
            in2 => \N__28550\,
            in3 => \N__29824\,
            lcout => \progRomAddress_9\,
            ltout => \progRomAddress_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_adflt_3_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__28537\,
            in1 => \N__28529\,
            in2 => \N__28523\,
            in3 => \N__64655\,
            lcout => \PROM.ROMDATA.dintern_adfltZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_10_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29842\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.tempCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_10C_net\,
            ce => \N__34964\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_9_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28495\,
            lcout => \CONTROL.tempCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_10C_net\,
            ce => \N__34964\,
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57728\,
            in2 => \_gnd_net_\,
            in3 => \N__41990\,
            lcout => \CONTROL.addrstack_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.addrstackptr_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNINS3U7_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33101\,
            in1 => \N__28640\,
            in2 => \_gnd_net_\,
            in3 => \N__49817\,
            lcout => bus_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN3QUB1_0_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__66602\,
            in1 => \N__66312\,
            in2 => \N__60263\,
            in3 => \N__65951\,
            lcout => \ALU.rshift_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5SIF41_4_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__59586\,
            in1 => \N__59874\,
            in2 => \N__56268\,
            in3 => \N__56115\,
            lcout => \ALU.d_RNI5SIF41Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_1_c_RNO_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__65952\,
            in1 => \N__65570\,
            in2 => \N__60629\,
            in3 => \N__66603\,
            lcout => \ALU.status_17_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0PI3E1_8_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__65965\,
            in1 => \N__62874\,
            in2 => \N__61976\,
            in3 => \N__68823\,
            lcout => \ALU.d_RNI0PI3E1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFGGBO_6_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__62273\,
            in1 => \_gnd_net_\,
            in2 => \N__62585\,
            in3 => \N__66601\,
            lcout => OPEN,
            ltout => \ALU.N_834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMQD952_6_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__65963\,
            in1 => \_gnd_net_\,
            in2 => \N__28586\,
            in3 => \N__42772\,
            lcout => \ALU.N_864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIUFQIG_7_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__62271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68256\,
            lcout => \ALU.d_RNIUFQIGZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIC6EBM2_2_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__68824\,
            in1 => \N__47985\,
            in2 => \N__45723\,
            in3 => \N__65964\,
            lcout => \ALU.d_RNIC6EBM2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITLGIL_7_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62270\,
            in2 => \_gnd_net_\,
            in3 => \N__68822\,
            lcout => \ALU.d_RNITLGILZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIB692D1_6_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__62272\,
            in1 => \N__65962\,
            in2 => \N__62584\,
            in3 => \N__66600\,
            lcout => \ALU.mult_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISRIE42_2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__66653\,
            in1 => \N__68940\,
            in2 => \N__68280\,
            in3 => \N__66010\,
            lcout => \ALU.lshift62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9OBVC_3_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__38065\,
            in1 => \N__28583\,
            in2 => \N__53288\,
            in3 => \N__34586\,
            lcout => \ALU.status_19_2\,
            ltout => \ALU.status_19_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJBM6G_3_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28661\,
            in3 => \N__60197\,
            lcout => \ALU.d_RNIJBM6GZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFBJI61_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__68941\,
            in1 => \N__65550\,
            in2 => \N__60628\,
            in3 => \N__68231\,
            lcout => \ALU.d_RNIFBJI61Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITK2D51_2_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__68232\,
            in1 => \N__66288\,
            in2 => \N__60264\,
            in3 => \N__68942\,
            lcout => \ALU.d_RNITK2D51Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI04H8G_3_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__60198\,
            in1 => \N__63289\,
            in2 => \_gnd_net_\,
            in3 => \N__68233\,
            lcout => \ALU.d_RNI04H8GZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI7U266_2_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__59865\,
            in1 => \N__49605\,
            in2 => \N__28658\,
            in3 => \N__50221\,
            lcout => \CONTROL.busState_1_RNI7U266Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_95_c_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34046\,
            in2 => \N__28847\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \ALU.mult_3_c3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_95_c_RNINLQ452_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30206\,
            in2 => \N__28859\,
            in3 => \N__28631\,
            lcout => \ALU.mult_3_4\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c3\,
            carryout => \ALU.mult_3_c4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_101_c_RNIKJVKQ1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30245\,
            in2 => \N__28628\,
            in3 => \N__28619\,
            lcout => \ALU.mult_3_5\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c4\,
            carryout => \ALU.mult_3_c5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_107_c_RNIILDTH1_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28616\,
            in2 => \N__28610\,
            in3 => \N__28601\,
            lcout => \ALU.mult_3_6\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c5\,
            carryout => \ALU.mult_3_c6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_113_c_RNIH8VLK1_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28790\,
            in2 => \N__28784\,
            in3 => \N__28772\,
            lcout => \ALU.mult_3_7\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c6\,
            carryout => \ALU.mult_3_c7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_119_c_RNI03FQK1_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28769\,
            in2 => \N__28763\,
            in3 => \N__28754\,
            lcout => \ALU.mult_3_8\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c7\,
            carryout => \ALU.mult_3_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_125_c_RNI84ENI1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28751\,
            in2 => \N__28745\,
            in3 => \N__28736\,
            lcout => \ALU.mult_3_9\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c8\,
            carryout => \ALU.mult_3_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_131_c_RNICCA4H1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28733\,
            in2 => \N__28808\,
            in3 => \N__28727\,
            lcout => \ALU.mult_3_10\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c9\,
            carryout => \ALU.mult_3_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_137_c_RNI7M9PJ1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28724\,
            in2 => \N__28820\,
            in3 => \N__28715\,
            lcout => \ALU.mult_3_11\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \ALU.mult_3_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_143_c_RNIUMAAM1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28712\,
            in2 => \N__28700\,
            in3 => \N__28685\,
            lcout => \ALU.mult_3_12\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c11\,
            carryout => \ALU.mult_3_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_149_c_RNIK33CN1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28682\,
            in2 => \N__28829\,
            in3 => \N__28667\,
            lcout => \ALU.mult_3_13\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c12\,
            carryout => \ALU.mult_3_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_155_c_RNI2IBOL1_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28796\,
            in2 => \N__28964\,
            in3 => \N__28664\,
            lcout => \ALU.mult_3_14\,
            ltout => OPEN,
            carryin => \ALU.mult_3_c13\,
            carryout => \ALU.mult_3_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_3_c14_THRU_LUT4_0_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28832\,
            lcout => \ALU.mult_3_c14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9E4F21_4_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55800\,
            in1 => \N__59588\,
            in2 => \N__55990\,
            in3 => \N__59833\,
            lcout => \ALU.d_RNI9E4F21Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIH49MH_1_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__65543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55799\,
            lcout => \ALU.d_RNIH49MHZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRJ3VH_1_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65542\,
            in2 => \_gnd_net_\,
            in3 => \N__56086\,
            lcout => \ALU.d_RNIRJ3VHZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI371041_8_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__62845\,
            in1 => \N__56116\,
            in2 => \N__56272\,
            in3 => \N__61901\,
            lcout => \ALU.d_RNI371041Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2IA441_2_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__66249\,
            in1 => \N__60213\,
            in2 => \N__57029\,
            in3 => \N__55577\,
            lcout => \ALU.d_RNI2IA441Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7SQI21_2_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55674\,
            in1 => \N__60209\,
            in2 => \N__55823\,
            in3 => \N__66248\,
            lcout => \ALU.d_RNI7SQI21Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIK8R951_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__60598\,
            in1 => \N__65493\,
            in2 => \N__57028\,
            in3 => \N__55578\,
            lcout => \ALU.d_RNIK8R951Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID31VF_3_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60208\,
            in2 => \_gnd_net_\,
            in3 => \N__55957\,
            lcout => \ALU.d_RNID31VFZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBRFE41_2_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__66250\,
            in1 => \N__60214\,
            in2 => \N__57030\,
            in3 => \N__56905\,
            lcout => \ALU.d_RNIBRFE41Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN3H0D_3_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010110000"
        )
    port map (
            in0 => \N__33058\,
            in1 => \N__53165\,
            in2 => \N__70012\,
            in3 => \N__38066\,
            lcout => \ALU.d_RNIN3H0DZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9IN2H_3_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60101\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57015\,
            lcout => \ALU.d_RNI9IN2HZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRD18N_2_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__60118\,
            in1 => \N__66251\,
            in2 => \_gnd_net_\,
            in3 => \N__66377\,
            lcout => \ALU.N_767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI2N741_12_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48269\,
            in2 => \N__51421\,
            in3 => \N__43309\,
            lcout => \ALU.a_RNI2N741Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILEAFE_0_5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__40594\,
            in1 => \N__28940\,
            in2 => \N__28922\,
            in3 => \N__28877\,
            lcout => \ALU.combOperand2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI693UN_3_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65929\,
            lcout => \ALU.d_RNI693UNZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_95_c_RNO_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60099\,
            in2 => \_gnd_net_\,
            in3 => \N__66376\,
            lcout => \ALU.mult_95_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI42AE1_11_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__39841\,
            in1 => \N__47284\,
            in2 => \N__35968\,
            in3 => \N__54304\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI88772_11_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__57981\,
            in1 => \N__36188\,
            in2 => \N__28835\,
            in3 => \N__47210\,
            lcout => \ALU.N_1144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI2TJC1_11_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__39842\,
            in1 => \_gnd_net_\,
            in2 => \N__35969\,
            in3 => \N__43310\,
            lcout => \ALU.b_RNI2TJC1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI4OEM1_11_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__36104\,
            in1 => \N__29081\,
            in2 => \N__35671\,
            in3 => \N__47211\,
            lcout => OPEN,
            ltout => \ALU.N_1096_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIF4474_11_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29015\,
            in2 => \N__29009\,
            in3 => \N__54142\,
            lcout => \aluOut_11\,
            ltout => \aluOut_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNICV1S5_1_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__29006\,
            in1 => \N__50341\,
            in2 => \N__28994\,
            in3 => \N__50219\,
            lcout => \N_204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBH5A2_11_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__29087\,
            in1 => \N__53936\,
            in2 => \N__28973\,
            in3 => \N__46836\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN5325_11_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__53937\,
            in1 => \N__36170\,
            in2 => \N__28991\,
            in3 => \N__28988\,
            lcout => OPEN,
            ltout => \ALU.operand2_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMR627_11_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30677\,
            in2 => \N__28979\,
            in3 => \N__71399\,
            lcout => OPEN,
            ltout => \ALU.d_RNIMR627Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVUCRD_11_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__30664\,
            in1 => \N__53161\,
            in2 => \N__28976\,
            in3 => \N__49588\,
            lcout => \ALU.status_19_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNIV5PU_11_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46935\,
            in2 => \N__37265\,
            in3 => \N__32599\,
            lcout => \ALU.a_RNIV5PUZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3MHF_11_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__35664\,
            in1 => \N__36103\,
            in2 => \N__46945\,
            in3 => \_gnd_net_\,
            lcout => \ALU.c_RNI3MHFZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI2QT51_11_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__37261\,
            in1 => \N__47285\,
            in2 => \N__32606\,
            in3 => \N__54303\,
            lcout => \ALU.dout_3_ns_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNICADA1_10_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__37075\,
            in1 => \N__36338\,
            in2 => \N__32636\,
            in3 => \N__32822\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBCLN1_10_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__35712\,
            in1 => \N__36137\,
            in2 => \N__29075\,
            in3 => \N__54292\,
            lcout => \ALU.N_1095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIEIPI1_10_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__39133\,
            in1 => \N__36339\,
            in2 => \N__36004\,
            in3 => \N__32823\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFSD82_10_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__58227\,
            in1 => \N__36035\,
            in2 => \N__29072\,
            in3 => \N__54293\,
            lcout => OPEN,
            ltout => \ALU.N_1143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNITCH94_10_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54128\,
            in1 => \_gnd_net_\,
            in2 => \N__29069\,
            in3 => \N__29066\,
            lcout => \aluOut_10\,
            ltout => \aluOut_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIDR6R7_0_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__30833\,
            in1 => \N__34482\,
            in2 => \N__29060\,
            in3 => \N__49785\,
            lcout => \CONTROL.bus_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILM2O3_8_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29033\,
            in1 => \N__54129\,
            in2 => \_gnd_net_\,
            in3 => \N__29027\,
            lcout => \aluOut_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.combOperand2_d_bm_7_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__29183\,
            in1 => \N__49532\,
            in2 => \N__29174\,
            in3 => \N__50124\,
            lcout => \ALU.combOperand2_d_bmZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_7_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29141\,
            in2 => \_gnd_net_\,
            in3 => \N__72101\,
            lcout => \CONTROL.ctrlOut_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_7C_net\,
            ce => \N__44452\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNIAQOJ_7_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29204\,
            in1 => \N__33391\,
            in2 => \_gnd_net_\,
            in3 => \N__50123\,
            lcout => \N_168\,
            ltout => \N_168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI77OM1_2_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__50126\,
            in1 => \N__49544\,
            in2 => \N__29177\,
            in3 => \N__29173\,
            lcout => OPEN,
            ltout => \CONTROL.bus_7_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNITSIT7_0_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000101"
        )
    port map (
            in0 => \N__49711\,
            in1 => \N__49534\,
            in2 => \N__29144\,
            in3 => \N__43769\,
            lcout => bus_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_23dflt_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29140\,
            in2 => \_gnd_net_\,
            in3 => \N__72100\,
            lcout => \controlWord_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIP3P31_0_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__49709\,
            in1 => \N__49533\,
            in2 => \_gnd_net_\,
            in3 => \N__50125\,
            lcout => \CONTROL.bus_7_a1_1_8\,
            ltout => \CONTROL.bus_7_a1_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIA1EN6_0_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__33167\,
            in1 => \N__61836\,
            in2 => \N__29123\,
            in3 => \N__49710\,
            lcout => \CONTROL.bus_sx_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_2_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__29597\,
            in1 => \N__70708\,
            in2 => \N__34399\,
            in3 => \N__70458\,
            lcout => \gpuAddress_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_2C_net\,
            ce => \N__30759\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_3_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__70455\,
            in1 => \N__58610\,
            in2 => \N__70764\,
            in3 => \N__44255\,
            lcout => \gpuAddress_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_2C_net\,
            ce => \N__30759\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_4_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__70514\,
            in1 => \N__70709\,
            in2 => \N__43403\,
            in3 => \N__44188\,
            lcout => \gpuAddress_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_2C_net\,
            ce => \N__30759\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_5_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__70456\,
            in1 => \N__29455\,
            in2 => \N__70765\,
            in3 => \N__40268\,
            lcout => \gpuAddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_2C_net\,
            ce => \N__30759\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_6_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__70828\,
            in1 => \N__70710\,
            in2 => \N__37445\,
            in3 => \N__70459\,
            lcout => \gpuAddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_2C_net\,
            ce => \N__30759\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_7_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__70457\,
            in1 => \N__43835\,
            in2 => \N__70766\,
            in3 => \N__29368\,
            lcout => \gpuAddress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_2C_net\,
            ce => \N__30759\,
            sr => \_gnd_net_\
        );

    \CONTROL.gpuAddReg_8_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31084\,
            in1 => \N__70711\,
            in2 => \N__48146\,
            in3 => \N__70460\,
            lcout => \gpuAddress_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuAddReg_2C_net\,
            ce => \N__30759\,
            sr => \_gnd_net_\
        );

    \CONTROL.ramWrite_5_m9_0_a2_0_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38597\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30790\,
            lcout => \CONTROL.N_346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuWrite_RNO_3_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000100"
        )
    port map (
            in0 => \N__41430\,
            in1 => \N__41241\,
            in2 => \N__36404\,
            in3 => \N__54688\,
            lcout => OPEN,
            ltout => \CONTROL.un1_busState119_1_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuWrite_RNO_1_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__41596\,
            in1 => \_gnd_net_\,
            in2 => \N__29207\,
            in3 => \N__54746\,
            lcout => \CONTROL.N_66_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuWrite_RNO_2_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__31462\,
            in1 => \N__38595\,
            in2 => \N__41698\,
            in3 => \N__41595\,
            lcout => OPEN,
            ltout => \CONTROL.gpuWrite_RNOZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuWrite_RNO_0_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__38596\,
            in1 => \N__38324\,
            in2 => \N__29498\,
            in3 => \N__30789\,
            lcout => \CONTROL.gpuWrite_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState101_3_0_a2_1_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__54687\,
            in1 => \N__44899\,
            in2 => \N__44773\,
            in3 => \N__44714\,
            lcout => \CONTROL.busState96\,
            ltout => \CONTROL.busState96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState101_3_0_1_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001111"
        )
    port map (
            in0 => \N__36605\,
            in1 => \_gnd_net_\,
            in2 => \N__29495\,
            in3 => \N__36494\,
            lcout => \CONTROL.un1_busState101_3_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.gpuWrite_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010001"
        )
    port map (
            in0 => \N__29492\,
            in1 => \N__29486\,
            in2 => \N__29473\,
            in3 => \N__29480\,
            lcout => \gpuWrite\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.gpuWriteC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_5_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__39986\,
            in1 => \N__70722\,
            in2 => \N__29456\,
            in3 => \N__70467\,
            lcout => \A5_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_5C_net\,
            ce => \N__70317\,
            sr => \_gnd_net_\
        );

    \RAM.un1_WR_105_0_3_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__29557\,
            in1 => \N__29344\,
            in2 => \_gnd_net_\,
            in3 => \N__31294\,
            lcout => OPEN,
            ltout => \RAM.un1_WR_105_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM.un1_WR_105_0_11_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__70369\,
            in1 => \N__31151\,
            in2 => \N__29417\,
            in3 => \N__29398\,
            lcout => \RAM.un1_WR_105_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_7_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__29369\,
            in1 => \N__70723\,
            in2 => \N__49091\,
            in3 => \N__70468\,
            lcout => \A7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_5C_net\,
            ce => \N__70317\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_18dflt_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__45767\,
            in1 => \N__72775\,
            in2 => \N__41012\,
            in3 => \N__72131\,
            lcout => \controlWord_18\,
            ltout => \controlWord_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_2_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35636\,
            in1 => \N__70721\,
            in2 => \N__29579\,
            in3 => \N__70466\,
            lcout => \A2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_5C_net\,
            ce => \N__70317\,
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_4_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111111111111"
        )
    port map (
            in0 => \N__42266\,
            in1 => \N__54659\,
            in2 => \N__72315\,
            in3 => \N__55471\,
            lcout => OPEN,
            ltout => \CONTROL.g0_3_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIFRI6PV_7_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__29516\,
            in1 => \N__38501\,
            in2 => \N__29546\,
            in3 => \N__38186\,
            lcout => \CONTROL.N_4_1\,
            ltout => \CONTROL.N_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_4_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__29708\,
            in1 => \N__60780\,
            in2 => \N__29543\,
            in3 => \N__29675\,
            lcout => \CONTROL.addrstackptrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.addrstackptr_4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI1MMTM91_3_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41977\,
            in1 => \N__34772\,
            in2 => \N__31481\,
            in3 => \N__60730\,
            lcout => \CONTROL.un1_addrstackptr_c4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_7_174_i_i_o2_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__44701\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54657\,
            lcout => \CONTROL.N_81_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_a7_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__45221\,
            in1 => \N__54658\,
            in2 => \N__63481\,
            in3 => \N__38273\,
            lcout => \CONTROL.g0_3_i_a7_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI5GMQ_14_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29603\,
            in1 => \N__29633\,
            in2 => \_gnd_net_\,
            in3 => \N__42081\,
            lcout => \CONTROL.N_429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_8_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31346\,
            lcout => \CONTROL.dout_reto_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIDTCV_15_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__33482\,
            in1 => \_gnd_net_\,
            in2 => \N__31424\,
            in3 => \N__29825\,
            lcout => \progRomAddress_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_11_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI5PM5H92_4_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__29707\,
            in1 => \N__29681\,
            in2 => \N__60805\,
            in3 => \N__29674\,
            lcout => \CONTROL.addrstackptr_8_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_14_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29647\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI8INO_11_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29627\,
            in1 => \N__29621\,
            in2 => \_gnd_net_\,
            in3 => \N__45120\,
            lcout => \N_426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_11_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30650\,
            lcout => \CONTROL.dout_reto_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m470_am_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__76624\,
            in1 => \N__75908\,
            in2 => \N__64265\,
            in3 => \N__64973\,
            lcout => \PROM.ROMDATA.m470_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_14_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30452\,
            lcout => \CONTROL.dout_reto_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50837\,
            in2 => \_gnd_net_\,
            in3 => \N__50904\,
            lcout => \CONTROL.un1_programCounter9_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_10_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29846\,
            lcout => \CONTROL.programCounter_1_reto_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_35_rep1_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__50905\,
            in1 => \_gnd_net_\,
            in2 => \N__50843\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter11_reto_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI6GNO_10_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45119\,
            in1 => \N__34895\,
            in2 => \_gnd_net_\,
            in3 => \N__29801\,
            lcout => \CONTROL.N_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNID7J31_1_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__73686\,
            in1 => \N__73574\,
            in2 => \_gnd_net_\,
            in3 => \N__73820\,
            lcout => \CONTROL.programCounter_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI45TU352_1_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__31492\,
            in1 => \N__31444\,
            in2 => \N__31531\,
            in3 => \N__31541\,
            lcout => \CONTROL.addrstackptr_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI19JNL91_0_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57761\,
            in2 => \_gnd_net_\,
            in3 => \N__41981\,
            lcout => \CONTROL.addrstackptr_RNI19JNL91Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_9_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40322\,
            lcout => \CONTROL.dout_reto_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_5_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57321\,
            in1 => \N__52637\,
            in2 => \_gnd_net_\,
            in3 => \N__39323\,
            lcout => \ALU.aZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73138\,
            ce => \N__71215\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIET09P_0_12_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__61195\,
            in1 => \N__61462\,
            in2 => \_gnd_net_\,
            in3 => \N__66598\,
            lcout => \ALU.N_614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICP0UG_5_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__59583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68281\,
            lcout => \ALU.d_RNICP0UGZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBK47O_8_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__61977\,
            in1 => \N__62872\,
            in2 => \_gnd_net_\,
            in3 => \N__66597\,
            lcout => \ALU.N_836\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6CL331_4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__59584\,
            in1 => \N__59894\,
            in2 => \N__68394\,
            in3 => \N__56401\,
            lcout => \ALU.d_RNI6CL331Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_173_c_RNO_0_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59582\,
            in2 => \_gnd_net_\,
            in3 => \N__66596\,
            lcout => \ALU.mult_173_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILJMRC1_8_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__66599\,
            in1 => \N__61978\,
            in2 => \N__62320\,
            in3 => \N__65954\,
            lcout => OPEN,
            ltout => \ALU.d_RNILJMRC1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITH0GI3_8_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30326\,
            in2 => \N__29861\,
            in3 => \N__48232\,
            lcout => \ALU.N_642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_239_c_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31721\,
            in2 => \N__31730\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \ALU.mult_7_c7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_239_c_RNI6DER62_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32864\,
            in2 => \N__29870\,
            in3 => \N__29858\,
            lcout => \ALU.mult_7_8\,
            ltout => OPEN,
            carryin => \ALU.mult_7_c7\,
            carryout => \ALU.mult_7_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_245_c_RNISI9DS1_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29855\,
            in2 => \N__29879\,
            in3 => \N__29849\,
            lcout => \ALU.mult_7_9\,
            ltout => OPEN,
            carryin => \ALU.mult_7_c8\,
            carryout => \ALU.mult_7_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_251_c_RNIH3GMJ1_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29993\,
            in2 => \N__29987\,
            in3 => \N__29969\,
            lcout => \ALU.mult_7_10\,
            ltout => OPEN,
            carryin => \ALU.mult_7_c9\,
            carryout => \ALU.mult_7_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_257_c_RNIP79EM1_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29966\,
            in2 => \N__29951\,
            in3 => \N__29933\,
            lcout => \ALU.mult_7_11\,
            ltout => OPEN,
            carryin => \ALU.mult_7_c10\,
            carryout => \ALU.mult_7_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_263_c_RNIVGHJM1_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29930\,
            in2 => \N__30098\,
            in3 => \N__29915\,
            lcout => \ALU.mult_7_12\,
            ltout => OPEN,
            carryin => \ALU.mult_7_c11\,
            carryout => \ALU.mult_7_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_269_c_RNIG3OFK1_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29912\,
            in2 => \N__37001\,
            in3 => \N__29900\,
            lcout => \ALU.mult_7_13\,
            ltout => OPEN,
            carryin => \ALU.mult_7_c12\,
            carryout => \ALU.mult_7_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_275_c_RNIKBKSI1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29897\,
            in2 => \N__46586\,
            in3 => \N__29885\,
            lcout => \ALU.mult_7_14\,
            ltout => OPEN,
            carryin => \ALU.mult_7_c13\,
            carryout => \ALU.mult_7_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_7_c14_THRU_LUT4_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29882\,
            lcout => \ALU.mult_7_c14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFGNR61_4_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__68745\,
            in1 => \N__59864\,
            in2 => \N__59599\,
            in3 => \N__68229\,
            lcout => \ALU.d_RNIFGNR61Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHNHG61_6_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__68230\,
            in1 => \N__62285\,
            in2 => \N__62557\,
            in3 => \N__68746\,
            lcout => \ALU.d_RNIHNHG61Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4LU7E1_6_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__68744\,
            in1 => \N__62519\,
            in2 => \N__62306\,
            in3 => \N__66011\,
            lcout => \ALU.d_RNI4LU7E1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJAJOO_0_10_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__62873\,
            in1 => \N__61666\,
            in2 => \_gnd_net_\,
            in3 => \N__66652\,
            lcout => \ALU.N_612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA6P2I_7_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62281\,
            in2 => \_gnd_net_\,
            in3 => \N__56267\,
            lcout => \ALU.d_RNIA6P2IZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIOGRG_1_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65520\,
            in2 => \_gnd_net_\,
            in3 => \N__68228\,
            lcout => \ALU.d_RNIIOGRGZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_5_c_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32063\,
            in2 => \N__30503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \ALU.mult_1_c1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_5_c_RNIFR9072_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32402\,
            in2 => \N__32411\,
            in3 => \N__30086\,
            lcout => \ALU.mult_1_2\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c1\,
            carryout => \ALU.mult_1_c2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_11_c_RNIL35NS1_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32099\,
            in2 => \N__30083\,
            in3 => \N__30074\,
            lcout => \ALU.mult_1_3\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c2\,
            carryout => \ALU.mult_1_c3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_17_c_RNIJ5JVJ1_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30071\,
            in2 => \N__30065\,
            in3 => \N__30050\,
            lcout => \ALU.mult_1_4\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c3\,
            carryout => \ALU.mult_1_c4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_23_c_RNIIO4OM1_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30047\,
            in2 => \N__30035\,
            in3 => \N__30023\,
            lcout => \ALU.mult_1_5\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c4\,
            carryout => \ALU.mult_1_c5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_29_c_RNI1JKSM1_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30020\,
            in2 => \N__30008\,
            in3 => \N__29996\,
            lcout => \ALU.mult_1_6\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c5\,
            carryout => \ALU.mult_1_c6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_35_c_RNI9KJPK1_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40163\,
            in2 => \N__30197\,
            in3 => \N__30185\,
            lcout => \ALU.mult_1_7\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c6\,
            carryout => \ALU.mult_1_c7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_41_c_RNIDSF6J1_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30182\,
            in2 => \N__33977\,
            in3 => \N__30170\,
            lcout => \ALU.mult_1_8\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c7\,
            carryout => \ALU.mult_1_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_47_c_RNI86FRL1_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30167\,
            in2 => \N__30254\,
            in3 => \N__30161\,
            lcout => \ALU.mult_1_9\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \ALU.mult_1_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_53_c_RNIV6GCO1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30260\,
            in2 => \N__30158\,
            in3 => \N__30146\,
            lcout => \ALU.mult_1_10\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c9\,
            carryout => \ALU.mult_1_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_59_c_RNILJ8EP1_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30143\,
            in2 => \N__30131\,
            in3 => \N__30122\,
            lcout => \ALU.mult_1_11\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c10\,
            carryout => \ALU.mult_1_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_65_c_RNI32HQN1_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30236\,
            in2 => \N__30575\,
            in3 => \N__30119\,
            lcout => \ALU.mult_1_12\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c11\,
            carryout => \ALU.mult_1_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_71_c_RNIPD3ES1_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30116\,
            in2 => \N__37205\,
            in3 => \N__30104\,
            lcout => \ALU.mult_1_13\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c12\,
            carryout => \ALU.mult_1_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_77_c_RNIF6U9Q1_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30230\,
            in2 => \N__30221\,
            in3 => \N__30101\,
            lcout => \ALU.mult_1_14\,
            ltout => OPEN,
            carryin => \ALU.mult_1_c13\,
            carryout => \ALU.mult_1_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_83_c_RNIKEU6B2_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30212\,
            in1 => \N__30284\,
            in2 => \N__30278\,
            in3 => \N__30263\,
            lcout => \ALU.mult_83_c_RNIKEU6BZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI83GO51_0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60542\,
            in1 => \N__65481\,
            in2 => \N__55686\,
            in3 => \N__55576\,
            lcout => \ALU.d_RNI83GO51Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPIBO31_0_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__65483\,
            in1 => \N__60541\,
            in2 => \N__55685\,
            in3 => \N__55821\,
            lcout => \ALU.d_RNIPIBO31Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIHC6L_3_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68658\,
            in2 => \_gnd_net_\,
            in3 => \N__60206\,
            lcout => \ALU.d_RNIIHC6LZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITH0K51_0_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__57039\,
            in1 => \N__56904\,
            in2 => \N__65546\,
            in3 => \N__60543\,
            lcout => \ALU.d_RNITH0K51Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0H41K_1_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56805\,
            in2 => \_gnd_net_\,
            in3 => \N__65479\,
            lcout => \ALU.d_RNI0H41KZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIETL861_0_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__65482\,
            in1 => \N__56737\,
            in2 => \N__56823\,
            in3 => \N__60544\,
            lcout => \ALU.d_RNIETL861Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8FM541_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__60545\,
            in1 => \N__74609\,
            in2 => \N__56748\,
            in3 => \N__65480\,
            lcout => \ALU.d_RNI8FM541Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGIF4D1_2_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__60207\,
            in1 => \N__66241\,
            in2 => \N__68733\,
            in3 => \N__66012\,
            lcout => \ALU.d_RNIGIF4D1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINLH9L_2_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001101000"
        )
    port map (
            in0 => \N__68720\,
            in1 => \N__74834\,
            in2 => \N__63290\,
            in3 => \N__66252\,
            lcout => \ALU.log_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN178L_2_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__66253\,
            in1 => \N__63248\,
            in2 => \_gnd_net_\,
            in3 => \N__68719\,
            lcout => \ALU.d_RNIN178LZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIBPDT_11_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30406\,
            in1 => \N__30377\,
            in2 => \_gnd_net_\,
            in3 => \N__64664\,
            lcout => \progRomAddress_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILJMRC1_0_8_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__62261\,
            in1 => \N__66441\,
            in2 => \N__61975\,
            in3 => \N__65930\,
            lcout => \ALU.d_RNILJMRC1_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI58QFI_5_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__59625\,
            in1 => \N__63249\,
            in2 => \_gnd_net_\,
            in3 => \N__33993\,
            lcout => \ALU.d_RNI58QFIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.combOperand2_1_0_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011011"
        )
    port map (
            in0 => \N__53145\,
            in1 => \N__36918\,
            in2 => \N__32846\,
            in3 => \N__38847\,
            lcout => OPEN,
            ltout => \ALU.combOperand2_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFFCPG_0_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001110"
        )
    port map (
            in0 => \N__71395\,
            in1 => \N__53146\,
            in2 => \N__30314\,
            in3 => \N__37870\,
            lcout => \ALU.status_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI6KJL_0_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32318\,
            in1 => \N__30473\,
            in2 => \_gnd_net_\,
            in3 => \N__30490\,
            lcout => OPEN,
            ltout => \DROM_ROMDATA_dintern_0ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIAR0U1_2_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__49562\,
            in1 => \N__30311\,
            in2 => \N__30299\,
            in3 => \N__30296\,
            lcout => \busState_1_RNIAR0U1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.combOperand2_a0_0_6_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71394\,
            in2 => \_gnd_net_\,
            in3 => \N__49793\,
            lcout => \ALU.combOperand2_a0_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIR8PGB_0_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__38848\,
            in1 => \N__49797\,
            in2 => \N__36925\,
            in3 => \N__32845\,
            lcout => bus_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_5_c_RNO_0_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__65351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66375\,
            lcout => \ALU.mult_5_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_0_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30491\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_0C_net\,
            ce => \N__32319\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_14_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30994\,
            in2 => \_gnd_net_\,
            in3 => \N__40915\,
            lcout => \CONTROL.ctrlOut_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_14C_net\,
            ce => \N__44453\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI6ADU_14_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30467\,
            in1 => \N__30445\,
            in2 => \_gnd_net_\,
            in3 => \N__50147\,
            lcout => OPEN,
            ltout => \CONTROL.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIHTF52_2_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__50148\,
            in1 => \N__30434\,
            in2 => \N__30413\,
            in3 => \N__49572\,
            lcout => \N_191\,
            ltout => \N_191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNISBR29_0_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__49573\,
            in1 => \N__47072\,
            in2 => \N__30410\,
            in3 => \N__49815\,
            lcout => bus_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_30dflt_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30993\,
            in2 => \_gnd_net_\,
            in3 => \N__40914\,
            lcout => \controlWord_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIRA1I6_2_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__49574\,
            in1 => \N__34099\,
            in2 => \N__50200\,
            in3 => \N__65408\,
            lcout => OPEN,
            ltout => \CONTROL.busState_1_RNIRA1I6Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI2BDF8_0_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49816\,
            in1 => \_gnd_net_\,
            in2 => \N__30578\,
            in3 => \N__33032\,
            lcout => bus_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8VHNH_1_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56987\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65407\,
            lcout => \ALU.d_RNI8VHNHZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI13B91_12_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__48265\,
            in1 => \N__43917\,
            in2 => \N__51422\,
            in3 => \N__32821\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI49JM1_12_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__52410\,
            in1 => \N__67549\,
            in2 => \N__30560\,
            in3 => \N__54294\,
            lcout => \ALU.N_1097\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI4EQI1_12_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__39817\,
            in1 => \N__34542\,
            in2 => \N__57686\,
            in3 => \N__43916\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9SE82_12_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__57934\,
            in1 => \N__65089\,
            in2 => \N__30557\,
            in3 => \N__54295\,
            lcout => OPEN,
            ltout => \ALU.N_1145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIG9G84_12_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30554\,
            in2 => \N__30548\,
            in3 => \N__54130\,
            lcout => \aluOut_12\,
            ltout => \aluOut_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI6CUR7_0_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__30587\,
            in1 => \N__34483\,
            in2 => \N__30545\,
            in3 => \N__49810\,
            lcout => \CONTROL.bus_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI04DU_11_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50106\,
            in1 => \N__30527\,
            in2 => \_gnd_net_\,
            in3 => \N__30643\,
            lcout => OPEN,
            ltout => \CONTROL.N_172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI8VQQ1_2_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__49494\,
            in1 => \N__30701\,
            in2 => \N__30680\,
            in3 => \N__50107\,
            lcout => \N_188\,
            ltout => \N_188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIQBOE8_0_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__30668\,
            in1 => \N__49811\,
            in2 => \N__30653\,
            in3 => \N__49495\,
            lcout => bus_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_11_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__72129\,
            in1 => \N__47475\,
            in2 => \N__72768\,
            in3 => \N__36950\,
            lcout => \CONTROL.ctrlOut_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_11C_net\,
            ce => \N__44415\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_27dflt_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__36949\,
            in1 => \N__72713\,
            in2 => \N__47488\,
            in3 => \N__72128\,
            lcout => \controlWord_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_12_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__72130\,
            in1 => \N__65150\,
            in2 => \N__72769\,
            in3 => \N__47476\,
            lcout => \CONTROL.ctrlOut_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_11C_net\,
            ce => \N__44415\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI26DU_12_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50104\,
            in1 => \N__30632\,
            in2 => \_gnd_net_\,
            in3 => \N__38764\,
            lcout => OPEN,
            ltout => \CONTROL.N_173_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIB9N32_2_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__49493\,
            in1 => \N__30611\,
            in2 => \N__30590\,
            in3 => \N__50105\,
            lcout => \CONTROL.N_189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState14_1_i_o2_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41245\,
            in1 => \N__41408\,
            in2 => \N__36883\,
            in3 => \N__54677\,
            lcout => \CONTROL.un1_busState14_1_i_o2_0\,
            ltout => \CONTROL.un1_busState14_1_i_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState12_2_i_a2_d_0_tz_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__30880\,
            in1 => \N__36433\,
            in2 => \N__30581\,
            in3 => \N__41246\,
            lcout => OPEN,
            ltout => \CONTROL.un1_busState12_2_i_a2_0_1_tz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState12_2_i_a2_0_i_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__36821\,
            in1 => \N__35171\,
            in2 => \N__30821\,
            in3 => \N__30791\,
            lcout => \CONTROL.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_1_sqmuxa_0_a2_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__30881\,
            in1 => \N__38717\,
            in2 => \N__36448\,
            in3 => \N__41248\,
            lcout => \CONTROL.aluReadBus_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState119_i_i_a2_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__36684\,
            in1 => \N__54678\,
            in2 => \N__41259\,
            in3 => \N__44708\,
            lcout => \CONTROL.N_244\,
            ltout => \CONTROL.N_244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36578\,
            in1 => \N__30809\,
            in2 => \N__30818\,
            in3 => \N__71314\,
            lcout => \aluReadBus\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluReadBusC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState98_1_1_0_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__41249\,
            in1 => \N__36443\,
            in2 => \_gnd_net_\,
            in3 => \N__33473\,
            lcout => \CONTROL.un1_busState98_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState14_1_i_a2_1_i_1_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__30879\,
            in1 => \N__30815\,
            in2 => \N__36447\,
            in3 => \N__41247\,
            lcout => \CONTROL.un1_busState14_1_i_a2_1_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_RNO_0_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__41429\,
            in1 => \N__30707\,
            in2 => \N__36609\,
            in3 => \N__44898\,
            lcout => \CONTROL.aluReadBus_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState14_1_i_a2_1_i_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__38323\,
            in1 => \N__30800\,
            in2 => \N__38657\,
            in3 => \N__30792\,
            lcout => \CONTROL.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState101_3_0_m2_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__41428\,
            in1 => \N__55474\,
            in2 => \N__36884\,
            in3 => \N__54670\,
            lcout => \CONTROL.N_89\,
            ltout => \CONTROL.N_89_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState101_3_0_0_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41594\,
            in2 => \N__30887\,
            in3 => \N__36688\,
            lcout => \CONTROL.un1_busState101_3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState103_0_o2_0_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44705\,
            in1 => \N__54668\,
            in2 => \N__41435\,
            in3 => \N__44897\,
            lcout => \CONTROL.N_101_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState97_1_0_o2_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__54669\,
            in1 => \N__55473\,
            in2 => \_gnd_net_\,
            in3 => \N__44707\,
            lcout => \CONTROL.N_87_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_1_sqmuxa_0_a2_0_0_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__55472\,
            in1 => \N__42244\,
            in2 => \_gnd_net_\,
            in3 => \N__72181\,
            lcout => OPEN,
            ltout => \CONTROL.aluReadBus_1_sqmuxa_0_a2_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100100111"
        )
    port map (
            in0 => \N__44896\,
            in1 => \N__36506\,
            in2 => \N__30884\,
            in3 => \N__44706\,
            lcout => \CONTROL.aluReadBus_1_sqmuxa_0_o2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_10_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010001010"
        )
    port map (
            in0 => \N__72191\,
            in1 => \N__73945\,
            in2 => \N__72790\,
            in3 => \N__62609\,
            lcout => \CONTROL.ctrlOut_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_10C_net\,
            ce => \N__44445\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNIU1DU_10_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30869\,
            in1 => \N__34906\,
            in2 => \_gnd_net_\,
            in3 => \N__50019\,
            lcout => OPEN,
            ltout => \CONTROL.N_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI5LU12_2_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__50021\,
            in1 => \N__30854\,
            in2 => \N__30836\,
            in3 => \N__49391\,
            lcout => \CONTROL.N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_26dflt_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100000000"
        )
    port map (
            in0 => \N__62608\,
            in1 => \N__72777\,
            in2 => \N__73946\,
            in3 => \N__72189\,
            lcout => \controlWord_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_0_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010001010"
        )
    port map (
            in0 => \N__72190\,
            in1 => \N__64057\,
            in2 => \N__72789\,
            in3 => \N__74330\,
            lcout => \CONTROL.ctrlOut_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_10C_net\,
            ce => \N__44445\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNISBOJ_0_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31028\,
            in1 => \N__45076\,
            in2 => \_gnd_net_\,
            in3 => \N__50020\,
            lcout => OPEN,
            ltout => \CONTROL.N_161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNII0IO1_2_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__50022\,
            in1 => \N__31010\,
            in2 => \N__30998\,
            in3 => \N__49392\,
            lcout => \N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_16dflt_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100000000"
        )
    port map (
            in0 => \N__74329\,
            in1 => \N__72776\,
            in2 => \N__64058\,
            in3 => \N__72188\,
            lcout => \controlWord_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.combOperand2_d_bm_15_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__50005\,
            in1 => \N__30941\,
            in2 => \N__30935\,
            in3 => \N__49545\,
            lcout => \ALU.combOperand2_d_bmZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_15_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__72193\,
            in1 => \N__30992\,
            in2 => \N__72791\,
            in3 => \N__47490\,
            lcout => \CONTROL.ctrlOut_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_15C_net\,
            ce => \N__44435\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31dflt_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__47489\,
            in1 => \N__72784\,
            in2 => \N__30995\,
            in3 => \N__72192\,
            lcout => \controlWord_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI8CDU_15_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30962\,
            in1 => \N__33433\,
            in2 => \_gnd_net_\,
            in3 => \N__50004\,
            lcout => \N_176\,
            ltout => \N_176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIK7CU1_2_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101110111"
        )
    port map (
            in0 => \N__50006\,
            in1 => \N__30934\,
            in2 => \N__30890\,
            in3 => \N__49546\,
            lcout => \CONTROL.bus_7_ns_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_8_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__31376\,
            in1 => \N__72785\,
            in2 => \N__47495\,
            in3 => \N__72194\,
            lcout => \CONTROL.ctrlOut_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_15C_net\,
            ce => \N__44435\,
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNICSOJ_8_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31367\,
            in1 => \N__31345\,
            in2 => \_gnd_net_\,
            in3 => \N__50003\,
            lcout => \CONTROL.N_169\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_0_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__33313\,
            in1 => \N__70754\,
            in2 => \N__49136\,
            in3 => \N__70525\,
            lcout => \A0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_0C_net\,
            ce => \N__70318\,
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_1_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__70523\,
            in1 => \N__33247\,
            in2 => \N__49181\,
            in3 => \N__70759\,
            lcout => \A1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_0C_net\,
            ce => \N__70318\,
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_10_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31275\,
            in1 => \N__70755\,
            in2 => \N__36008\,
            in3 => \N__70526\,
            lcout => \A10_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_0C_net\,
            ce => \N__70318\,
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_11_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__70522\,
            in1 => \N__35967\,
            in2 => \N__31238\,
            in3 => \N__70758\,
            lcout => \A11_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_0C_net\,
            ce => \N__70318\,
            sr => \_gnd_net_\
        );

    \RAM.un1_WR_105_0_9_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31039\,
            in1 => \N__31192\,
            in2 => \N__31168\,
            in3 => \N__31096\,
            lcout => \RAM.un1_WR_105_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_9_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__48998\,
            in1 => \N__70756\,
            in2 => \N__31136\,
            in3 => \N__70527\,
            lcout => \A9_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_0C_net\,
            ce => \N__70318\,
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_8_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__70524\,
            in1 => \N__49052\,
            in2 => \N__31085\,
            in3 => \N__70760\,
            lcout => \A8_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_0C_net\,
            ce => \N__70318\,
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI0N94M91_1_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__38415\,
            in1 => \N__57809\,
            in2 => \_gnd_net_\,
            in3 => \N__41960\,
            lcout => \CONTROL.g1_0\,
            ltout => \CONTROL.g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_1_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__31445\,
            in1 => \N__31535\,
            in2 => \N__31499\,
            in3 => \N__31493\,
            lcout => \CONTROL.addrstackptrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.addrstackptr_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_1_i_a6_4_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__42264\,
            in1 => \N__36281\,
            in2 => \N__48488\,
            in3 => \N__38216\,
            lcout => OPEN,
            ltout => \CONTROL.g0_1_i_a6Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_1_i_a6_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40709\,
            in2 => \N__31496\,
            in3 => \N__40691\,
            lcout => \CONTROL.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNITQCP_1_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38411\,
            in2 => \_gnd_net_\,
            in3 => \N__57808\,
            lcout => \CONTROL.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState_1_sqmuxa_i_a2_2_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__42263\,
            in1 => \N__55399\,
            in2 => \N__72306\,
            in3 => \N__71854\,
            lcout => \CONTROL.N_366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI94D27G_7_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__72271\,
            in1 => \N__55475\,
            in2 => \N__36650\,
            in3 => \N__41496\,
            lcout => \CONTROL.g0_1_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_15_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31433\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.addrstack_reto_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_14_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31404\,
            in1 => \N__70757\,
            in2 => \N__57593\,
            in3 => \N__70521\,
            lcout => \A14_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_14C_net\,
            ce => \N__70328\,
            sr => \_gnd_net_\
        );

    \ALU.mult_173_c_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33713\,
            in2 => \N__31688\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \ALU.mult_5_c5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_173_c_RNIFBQH72_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33947\,
            in2 => \N__32093\,
            in3 => \N__31679\,
            lcout => \ALU.mult_5_6\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c5\,
            carryout => \ALU.mult_5_c6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_179_c_RNIE2T2T1_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31676\,
            in2 => \N__33959\,
            in3 => \N__31667\,
            lcout => \ALU.mult_5_7\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c6\,
            carryout => \ALU.mult_5_c7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_185_c_RNI3J3CK1_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31664\,
            in2 => \N__31658\,
            in3 => \N__31649\,
            lcout => \ALU.mult_5_8\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c7\,
            carryout => \ALU.mult_5_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_191_c_RNI26L4N1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31646\,
            in2 => \N__33773\,
            in3 => \N__31634\,
            lcout => \ALU.mult_5_9\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c8\,
            carryout => \ALU.mult_5_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_197_c_RNIH059N1_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31631\,
            in2 => \N__31619\,
            in3 => \N__31607\,
            lcout => \ALU.mult_5_10\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c9\,
            carryout => \ALU.mult_5_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_203_c_RNIG7BVK1_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31604\,
            in2 => \N__31589\,
            in3 => \N__31574\,
            lcout => \ALU.mult_5_11\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c10\,
            carryout => \ALU.mult_5_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_209_c_RNIT0FBJ1_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31571\,
            in2 => \N__31559\,
            in3 => \N__31544\,
            lcout => \ALU.mult_5_12\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c11\,
            carryout => \ALU.mult_5_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_215_c_RNIFP61M1_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31862\,
            in2 => \N__31850\,
            in3 => \N__31838\,
            lcout => \ALU.mult_5_13\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \ALU.mult_5_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_221_c_RNI6Q7IO1_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31835\,
            in2 => \N__31826\,
            in3 => \N__31811\,
            lcout => \ALU.mult_5_14\,
            ltout => OPEN,
            carryin => \ALU.mult_5_c13\,
            carryout => \ALU.mult_5_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_227_c_RNIBPRV92_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31808\,
            in1 => \N__31802\,
            in2 => \N__31787\,
            in3 => \N__31769\,
            lcout => \ALU.mult_227_c_RNIBPRVZ0Z92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILTVJG3_3_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001111"
        )
    port map (
            in0 => \N__57238\,
            in1 => \N__56465\,
            in2 => \N__70016\,
            in3 => \N__31766\,
            lcout => \ALU.d_RNILTVJG3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_239_c_RNO_0_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__62269\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66570\,
            lcout => \ALU.mult_239_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_239_c_RNO_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__65828\,
            in1 => \N__62314\,
            in2 => \N__66696\,
            in3 => \N__62523\,
            lcout => \ALU.mult_239_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_5_c_RNI6LDHN2_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__31714\,
            in1 => \N__33806\,
            in2 => \N__31715\,
            in3 => \_gnd_net_\,
            lcout => \ALU.mult_2\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \ALU.mult_17_c2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_388_c_RNI23SO83_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34112\,
            in2 => \N__31700\,
            in3 => \N__31691\,
            lcout => \ALU.mult_3\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c2\,
            carryout => \ALU.mult_17_c3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_391_c_RNIQB68P3_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32057\,
            in2 => \N__32045\,
            in3 => \N__32036\,
            lcout => \ALU.mult_17_4\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c3\,
            carryout => \ALU.mult_17_c4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_394_c_RNIP20HH3_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32033\,
            in2 => \N__32027\,
            in3 => \N__32012\,
            lcout => \ALU.mult_17_5\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c4\,
            carryout => \ALU.mult_17_c5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_397_c_RNI951U83_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32009\,
            in2 => \N__32000\,
            in3 => \N__31985\,
            lcout => \ALU.mult_17_6\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c5\,
            carryout => \ALU.mult_17_c6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_400_c_RNI1KKT93_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31982\,
            in2 => \N__31976\,
            in3 => \N__31961\,
            lcout => \ALU.mult_17_7\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c6\,
            carryout => \ALU.mult_17_c7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_403_c_RNINS3F83_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31958\,
            in2 => \N__31952\,
            in3 => \N__31937\,
            lcout => \ALU.mult_17_8\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c7\,
            carryout => \ALU.mult_17_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_406_c_RNITD5193_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31934\,
            in2 => \N__31925\,
            in3 => \N__31910\,
            lcout => \ALU.mult_17_9\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c8\,
            carryout => \ALU.mult_17_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_409_c_RNIRS5V93_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31907\,
            in2 => \N__31898\,
            in3 => \N__31889\,
            lcout => \ALU.mult_17_10\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \ALU.mult_17_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_412_c_RNI68PMD3_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31886\,
            in2 => \N__31880\,
            in3 => \N__31865\,
            lcout => \ALU.mult_17_11\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c10\,
            carryout => \ALU.mult_17_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_415_c_RNIET5KE3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32189\,
            in2 => \N__32183\,
            in3 => \N__32168\,
            lcout => \ALU.mult_17_12\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c11\,
            carryout => \ALU.mult_17_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_418_c_RNITRJ9K3_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32165\,
            in2 => \N__32159\,
            in3 => \N__32144\,
            lcout => \ALU.mult_17_13\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c12\,
            carryout => \ALU.mult_17_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_421_c_RNIRNI2G3_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32141\,
            in2 => \N__32135\,
            in3 => \N__32120\,
            lcout => \ALU.mult_17_14\,
            ltout => OPEN,
            carryin => \ALU.mult_17_c13\,
            carryout => \ALU.mult_17_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_424_c_RNIUVTAL4_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32117\,
            in1 => \N__32108\,
            in2 => \N__33815\,
            in3 => \N__32102\,
            lcout => \ALU.mult_424_c_RNIUVTALZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHU6RL_1_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65521\,
            in2 => \_gnd_net_\,
            in3 => \N__68728\,
            lcout => \ALU.d_RNIHU6RLZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2E4JE1_4_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__65715\,
            in1 => \N__68660\,
            in2 => \N__59624\,
            in3 => \N__59903\,
            lcout => \ALU.d_RNI2E4JE1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISLOMK_0_1_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101010011"
        )
    port map (
            in0 => \N__34100\,
            in1 => \N__34685\,
            in2 => \N__53249\,
            in3 => \N__34067\,
            lcout => \ALU.addsub_axb_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFCCRV4_4_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39229\,
            in1 => \N__68661\,
            in2 => \_gnd_net_\,
            in3 => \N__32078\,
            lcout => \ALU.N_920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_5_c_RNO_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__60539\,
            in1 => \N__65446\,
            in2 => \N__66755\,
            in3 => \N__65711\,
            lcout => \ALU.mult_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI290AE1_0_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__65445\,
            in1 => \N__68659\,
            in2 => \N__65826\,
            in3 => \N__60540\,
            lcout => \ALU.d_RNI290AE1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5MTIO_1_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65444\,
            in2 => \_gnd_net_\,
            in3 => \N__65710\,
            lcout => \ALU.d_RNI5MTIOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNICT0U1_2_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__49519\,
            in1 => \N__50337\,
            in2 => \N__32357\,
            in3 => \N__50197\,
            lcout => \busState_1_RNICT0U1_2\,
            ltout => \busState_1_RNICT0U1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8U1VH_2_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111000100"
        )
    port map (
            in0 => \N__32758\,
            in1 => \N__53204\,
            in2 => \N__32396\,
            in3 => \N__32937\,
            lcout => \ALU.status_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8U1VH_0_2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111000100"
        )
    port map (
            in0 => \N__32759\,
            in1 => \N__53205\,
            in2 => \N__32393\,
            in3 => \N__32938\,
            lcout => \ALU.lshift_15_0_sx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNILM6T5_2_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__66228\,
            in1 => \N__32392\,
            in2 => \N__49582\,
            in3 => \N__50198\,
            lcout => \N_227_0\,
            ltout => \N_227_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_2_c_RNO_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__53216\,
            in1 => \N__66229\,
            in2 => \N__32381\,
            in3 => \N__32939\,
            lcout => \ALU.status_18_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_RNI8MJL_2_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32330\,
            in1 => \N__32347\,
            in2 => \_gnd_net_\,
            in3 => \N__32322\,
            lcout => \DROM_ROMDATA_dintern_2ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DROM.ROMDATA.dintern_0_0_OLD_ne_2_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DROM.ROMDATA.dintern_0_0_OLDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDROM.ROMDATA.dintern_0_0_OLD_ne_2C_net\,
            ce => \N__32323\,
            sr => \_gnd_net_\
        );

    \ALU.e_2_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39456\,
            in1 => \N__39604\,
            in2 => \_gnd_net_\,
            in3 => \N__39516\,
            lcout => \ALU.eZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73153\,
            ce => \N__69244\,
            sr => \_gnd_net_\
        );

    \ALU.e_4_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39391\,
            in1 => \N__57420\,
            in2 => \_gnd_net_\,
            in3 => \N__42551\,
            lcout => \ALU.eZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73153\,
            ce => \N__69244\,
            sr => \_gnd_net_\
        );

    \ALU.e_5_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57419\,
            in1 => \N__52627\,
            in2 => \_gnd_net_\,
            in3 => \N__39322\,
            lcout => \ALU.eZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73153\,
            ce => \N__69244\,
            sr => \_gnd_net_\
        );

    \ALU.e_6_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43067\,
            in1 => \N__43121\,
            in2 => \_gnd_net_\,
            in3 => \N__42991\,
            lcout => \ALU.eZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73153\,
            ce => \N__69244\,
            sr => \_gnd_net_\
        );

    \ALU.e_3_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__58799\,
            in1 => \N__58757\,
            in2 => \_gnd_net_\,
            in3 => \N__58666\,
            lcout => \ALU.eZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73153\,
            ce => \N__69244\,
            sr => \_gnd_net_\
        );

    \ALU.e_10_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58510\,
            in1 => \N__58371\,
            in2 => \_gnd_net_\,
            in3 => \N__58300\,
            lcout => \ALU.eZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73153\,
            ce => \N__69244\,
            sr => \_gnd_net_\
        );

    \ALU.e_11_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58194\,
            in2 => \N__58126\,
            in3 => \N__58058\,
            lcout => \ALU.eZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73153\,
            ce => \N__69244\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIAHH51_6_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__43912\,
            in1 => \N__70603\,
            in2 => \N__39895\,
            in3 => \N__34556\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMOPK1_6_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__37434\,
            in1 => \N__36055\,
            in2 => \N__32735\,
            in3 => \N__47188\,
            lcout => \ALU.N_1139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI8BB31_6_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__43913\,
            in1 => \N__42941\,
            in2 => \N__32728\,
            in3 => \N__34557\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIICD02_6_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__35764\,
            in1 => \N__35833\,
            in2 => \N__32708\,
            in3 => \N__47189\,
            lcout => OPEN,
            ltout => \ALU.N_1091_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIB9LU3_6_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54110\,
            in2 => \N__32705\,
            in3 => \N__32702\,
            lcout => \aluOut_6\,
            ltout => \aluOut_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIR3N75_6_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__53144\,
            in1 => \N__49563\,
            in2 => \N__32696\,
            in3 => \N__50143\,
            lcout => \ALU.d_RNIR3N75Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI3N941_1_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__47144\,
            in1 => \N__49164\,
            in2 => \N__47271\,
            in3 => \N__48410\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5KHJ1_1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__37512\,
            in1 => \N__47145\,
            in2 => \N__32675\,
            in3 => \N__52165\,
            lcout => \ALU_N_1134\,
            ltout => \ALU_N_1134_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_RNIR8FK7_0_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32669\,
            in2 => \N__32672\,
            in3 => \N__34286\,
            lcout => \operand1_ne_RNIR8FK7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_RNIBQE03_0_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__54113\,
            in1 => \N__50131\,
            in2 => \N__49579\,
            in3 => \N__34298\,
            lcout => \CONTROL.operand1_ne_RNIBQE03Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI9P5V3_2_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__50132\,
            in1 => \N__49512\,
            in2 => \_gnd_net_\,
            in3 => \N__66127\,
            lcout => \busState_1_RNI9P5V3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI1H321_1_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__37234\,
            in1 => \N__47142\,
            in2 => \N__46351\,
            in3 => \N__47246\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI185V1_1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__47143\,
            in1 => \N__48942\,
            in2 => \N__32747\,
            in3 => \N__46462\,
            lcout => \ALU_N_1086\,
            ltout => \ALU_N_1086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI905S3_1_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54114\,
            in1 => \_gnd_net_\,
            in2 => \N__32744\,
            in3 => \N__32741\,
            lcout => \aluOut_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_1_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100001110"
        )
    port map (
            in0 => \N__79431\,
            in1 => \N__72722\,
            in2 => \N__34433\,
            in3 => \N__54362\,
            lcout => \aluOperand1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_ne_1C_net\,
            ce => \N__36240\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_fast_ne_2_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101001010"
        )
    port map (
            in0 => \N__72721\,
            in1 => \N__50487\,
            in2 => \N__45059\,
            in3 => \N__41052\,
            lcout => \aluOperand1_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_ne_1C_net\,
            ce => \N__36240\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_2_rep1_ne_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__45050\,
            in1 => \N__41053\,
            in2 => \N__50494\,
            in3 => \N__72723\,
            lcout => \aluOperand1_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_ne_1C_net\,
            ce => \N__36240\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_2_rep2_ne_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101001010"
        )
    port map (
            in0 => \N__72720\,
            in1 => \N__50486\,
            in2 => \N__45058\,
            in3 => \N__41051\,
            lcout => \aluOperand1_2_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_ne_1C_net\,
            ce => \N__36240\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_2_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__45051\,
            in1 => \N__41054\,
            in2 => \N__50495\,
            in3 => \N__72724\,
            lcout => \aluOperand1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_ne_1C_net\,
            ce => \N__36240\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPTT4O_0_8_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__61881\,
            in1 => \N__62191\,
            in2 => \_gnd_net_\,
            in3 => \N__66569\,
            lcout => \ALU.N_610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHD7AO_7_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62190\,
            in2 => \_gnd_net_\,
            in3 => \N__65931\,
            lcout => \ALU.d_RNIHD7AOZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNICDG51_0_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__48376\,
            in1 => \N__36315\,
            in2 => \N__49132\,
            in3 => \N__32809\,
            lcout => \ALU.dout_6_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_RNIHKCU2_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__50103\,
            in1 => \N__54061\,
            in2 => \N__49528\,
            in3 => \N__32767\,
            lcout => OPEN,
            ltout => \CONTROL.operand1_ne_RNIHKCU2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_RNIDN8E7_0_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32776\,
            in2 => \N__32849\,
            in3 => \N__32783\,
            lcout => \operand1_ne_RNIDN8E7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBEFH1_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__51971\,
            in1 => \N__54236\,
            in2 => \N__37561\,
            in3 => \N__32831\,
            lcout => \ALU_N_1133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIA7A31_0_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__46324\,
            in1 => \N__32810\,
            in2 => \N__37589\,
            in3 => \N__36316\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI723T1_0_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__48900\,
            in1 => \N__46433\,
            in2 => \N__32789\,
            in3 => \N__54235\,
            lcout => \ALU_N_1085\,
            ltout => \ALU_N_1085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_RNIHKCU2_0_0_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__54060\,
            in1 => \N__49431\,
            in2 => \N__32786\,
            in3 => \N__50102\,
            lcout => \CONTROL.operand1_ne_RNIHKCU2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILK0O3_0_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32777\,
            in1 => \N__54062\,
            in2 => \_gnd_net_\,
            in3 => \N__32768\,
            lcout => \aluOut_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI1C5B1_2_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__53584\,
            in1 => \N__35632\,
            in2 => \N__39422\,
            in3 => \N__53480\,
            lcout => \ALU.operand2_6_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIV5V81_2_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__34352\,
            in1 => \N__53583\,
            in2 => \N__34334\,
            in3 => \N__53479\,
            lcout => OPEN,
            ltout => \ALU.operand2_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI0C2B2_2_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__35566\,
            in1 => \N__35876\,
            in2 => \N__32960\,
            in3 => \N__53429\,
            lcout => \ALU.N_1199\,
            ltout => \ALU.N_1199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJ1JO4_2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__43494\,
            in1 => \N__71320\,
            in2 => \N__32957\,
            in3 => \N__53941\,
            lcout => \ALU.c_RNIJ1JO4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJ1JO4_0_2_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__53942\,
            in1 => \N__32954\,
            in2 => \N__71384\,
            in3 => \N__43495\,
            lcout => OPEN,
            ltout => \ALU.c_RNIJ1JO4_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIARKGB_2_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32918\,
            in2 => \N__32948\,
            in3 => \N__32945\,
            lcout => \ALU.d_RNIARKGBZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4OEV1_2_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__36083\,
            in1 => \N__32924\,
            in2 => \N__34403\,
            in3 => \N__53430\,
            lcout => \ALU.N_1247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI48DU_13_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32912\,
            in1 => \N__43669\,
            in2 => \_gnd_net_\,
            in3 => \N__50009\,
            lcout => OPEN,
            ltout => \CONTROL.N_174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIEJJS1_2_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__50010\,
            in1 => \N__32891\,
            in2 => \N__32867\,
            in3 => \N__49341\,
            lcout => \CONTROL.N_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIAHKF1_2_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__49340\,
            in1 => \N__33200\,
            in2 => \N__33191\,
            in3 => \N__50008\,
            lcout => \CONTROL.N_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_2_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__41615\,
            in1 => \N__40625\,
            in2 => \N__49505\,
            in3 => \N__34697\,
            lcout => \busState_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.busState_1_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIU83C1_0_2_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__49342\,
            in1 => \N__37993\,
            in2 => \N__33139\,
            in3 => \N__50011\,
            lcout => \CONTROL.busState_1_RNIU83C1_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIOKAQ1_2_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__49339\,
            in1 => \N__34829\,
            in2 => \N__33086\,
            in3 => \N__50007\,
            lcout => \N_179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIBKBS7_0_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__33065\,
            in1 => \N__33380\,
            in2 => \_gnd_net_\,
            in3 => \N__49802\,
            lcout => bus_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNILAEH1_2_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__49946\,
            in1 => \N__49322\,
            in2 => \N__32993\,
            in3 => \N__32984\,
            lcout => \CONTROL.busState_1_RNILAEH1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNIUDOJ_1_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33017\,
            in1 => \N__50662\,
            in2 => \_gnd_net_\,
            in3 => \N__49942\,
            lcout => \N_162\,
            ltout => \N_162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.combOperand2_d_bm_1_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__49943\,
            in1 => \N__32983\,
            in2 => \N__32963\,
            in3 => \N__49320\,
            lcout => \ALU.combOperand2_d_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_1_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__34868\,
            in1 => \N__40637\,
            in2 => \N__50186\,
            in3 => \N__34712\,
            lcout => \busState_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.busState_1_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_a7_3_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__39779\,
            in1 => \N__45410\,
            in2 => \N__45515\,
            in3 => \N__54660\,
            lcout => \CONTROL.g0_3_i_a7_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIRU6J1_2_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__49323\,
            in1 => \N__33344\,
            in2 => \N__33353\,
            in3 => \N__49947\,
            lcout => \CONTROL.N_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI2IOJ_3_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49944\,
            in1 => \N__33374\,
            in2 => \_gnd_net_\,
            in3 => \N__45280\,
            lcout => \N_164\,
            ltout => \N_164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.combOperand2_d_bm_3_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__49321\,
            in1 => \N__33343\,
            in2 => \N__33320\,
            in3 => \N__49945\,
            lcout => \ALU.combOperand2_d_bmZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_0_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__71828\,
            in1 => \N__33306\,
            in2 => \N__48914\,
            in3 => \N__72178\,
            lcout => \CONTROL_romAddReg_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_17dflt_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__72177\,
            in1 => \N__38869\,
            in2 => \N__63968\,
            in3 => \N__72681\,
            lcout => \controlWord_17\,
            ltout => \controlWord_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_1_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__71829\,
            in1 => \N__48950\,
            in2 => \N__33236\,
            in3 => \N__72179\,
            lcout => \CONTROL_romAddReg_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m375_am_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110001011"
        )
    port map (
            in0 => \N__74480\,
            in1 => \N__76593\,
            in2 => \N__73394\,
            in3 => \N__75969\,
            lcout => \PROM.ROMDATA.m375_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_1_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__72682\,
            in1 => \N__63967\,
            in2 => \N__38873\,
            in3 => \N__72180\,
            lcout => \CONTROL.ctrlOut_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_1C_net\,
            ce => \N__44434\,
            sr => \_gnd_net_\
        );

    \CONTROL.busState104_2_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__72176\,
            in1 => \N__71827\,
            in2 => \_gnd_net_\,
            in3 => \N__44679\,
            lcout => \CONTROL.N_384_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_35_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50841\,
            in2 => \_gnd_net_\,
            in3 => \N__50906\,
            lcout => \CONTROL_programCounter11_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI7IMQ_15_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33440\,
            in1 => \N__33422\,
            in2 => \_gnd_net_\,
            in3 => \N__42082\,
            lcout => \CONTROL.N_430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState98_1_1_0_0_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111001"
        )
    port map (
            in0 => \N__44702\,
            in1 => \N__36680\,
            in2 => \N__41261\,
            in3 => \N__54655\,
            lcout => \CONTROL.un1_busState98_1_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_15_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_15_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33434\,
            lcout => \CONTROL.dout_reto_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m465_am_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__74491\,
            in1 => \N__76633\,
            in2 => \_gnd_net_\,
            in3 => \N__75973\,
            lcout => \PROM.ROMDATA.m465_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m299_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000100000"
        )
    port map (
            in0 => \N__78853\,
            in1 => \N__78060\,
            in2 => \N__76004\,
            in3 => \N__77308\,
            lcout => \PROM.ROMDATA.m299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_7_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33401\,
            lcout => \CONTROL.dout_reto_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_0_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__47408\,
            in1 => \N__73636\,
            in2 => \_gnd_net_\,
            in3 => \N__50969\,
            lcout => \CONTROL.tempCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_0C_net\,
            ce => \N__34954\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_5_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41740\,
            lcout => \CONTROL.tempCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_0C_net\,
            ce => \N__34954\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_3_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51148\,
            lcout => \CONTROL.tempCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_0C_net\,
            ce => \N__34954\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_8_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33587\,
            lcout => \CONTROL.tempCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_0C_net\,
            ce => \N__34954\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_4_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.tempCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_4C_net\,
            ce => \N__34965\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_1_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45188\,
            lcout => \CONTROL.tempCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_4C_net\,
            ce => \N__34965\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_7_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__73348\,
            lcout => \CONTROL.tempCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_4C_net\,
            ce => \N__34965\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_12_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36778\,
            lcout => \CONTROL.tempCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_4C_net\,
            ce => \N__34965\,
            sr => \_gnd_net_\
        );

    \CONTROL.tempCounter_2_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45316\,
            lcout => \CONTROL.tempCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.tempCounter_4C_net\,
            ce => \N__34965\,
            sr => \_gnd_net_\
        );

    \CONTROL.addrstack_addrstack_0_0_RNO_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57751\,
            lcout => \CONTROL.addrstack_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNII2KJ41_4_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__56415\,
            in1 => \N__59618\,
            in2 => \N__59902\,
            in3 => \N__56266\,
            lcout => \ALU.d_RNII2KJ41Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIR6J013_2_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__33744\,
            in1 => \N__56473\,
            in2 => \N__68932\,
            in3 => \N__69977\,
            lcout => \ALU.d_RNIR6J013Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_173_c_RNO_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__59884\,
            in1 => \N__59619\,
            in2 => \N__66029\,
            in3 => \N__66754\,
            lcout => \ALU.mult_173_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI68LSH_9_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62785\,
            in2 => \_gnd_net_\,
            in3 => \N__56414\,
            lcout => \ALU.d_RNI68LSHZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_173_c_RNIO8AO16_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__35236\,
            in1 => \N__35330\,
            in2 => \N__33707\,
            in3 => \_gnd_net_\,
            lcout => \ALU.mult_173_c_RNIO8AOZ0Z16\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \ALU.mult_19_c6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_432_c_RNI5DJ6A3_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33698\,
            in2 => \N__33689\,
            in3 => \N__33680\,
            lcout => \ALU.mult_19_7\,
            ltout => OPEN,
            carryin => \ALU.mult_19_c6\,
            carryout => \ALU.mult_19_c7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_435_c_RNIOA29R3_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33677\,
            in2 => \N__33665\,
            in3 => \N__33656\,
            lcout => \ALU.mult_19_8\,
            ltout => OPEN,
            carryin => \ALU.mult_19_c7\,
            carryout => \ALU.mult_19_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_438_c_RNIG9IJJ3_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33653\,
            in2 => \N__33644\,
            in3 => \N__33935\,
            lcout => \ALU.mult_19_9\,
            ltout => OPEN,
            carryin => \ALU.mult_19_c8\,
            carryout => \ALU.mult_19_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_441_c_RNIE942B3_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33932\,
            in2 => \N__33923\,
            in3 => \N__33914\,
            lcout => \ALU.mult_19_10\,
            ltout => OPEN,
            carryin => \ALU.mult_19_c9\,
            carryout => \ALU.mult_19_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_444_c_RNIOQ6GB3_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33911\,
            in2 => \N__33902\,
            in3 => \N__33890\,
            lcout => \ALU.mult_19_11\,
            ltout => OPEN,
            carryin => \ALU.mult_19_c10\,
            carryout => \ALU.mult_19_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_447_c_RNIE3M1A3_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33887\,
            in2 => \N__33881\,
            in3 => \N__33869\,
            lcout => \ALU.mult_19_12\,
            ltout => OPEN,
            carryin => \ALU.mult_19_c11\,
            carryout => \ALU.mult_19_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_450_c_RNIB3GKA3_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33866\,
            in2 => \N__33860\,
            in3 => \N__33845\,
            lcout => \ALU.mult_19_13\,
            ltout => OPEN,
            carryin => \ALU.mult_19_c12\,
            carryout => \ALU.mult_19_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_453_c_RNI9IGIB3_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33842\,
            in2 => \N__33836\,
            in3 => \N__33821\,
            lcout => \ALU.mult_19_14\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \ALU.mult_19_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_19_c14_THRU_LUT4_0_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33818\,
            lcout => \ALU.mult_19_c14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINP3HG_2_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000000000"
        )
    port map (
            in0 => \N__39101\,
            in1 => \N__53290\,
            in2 => \N__39047\,
            in3 => \N__66176\,
            lcout => \ALU.mult_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIMNQ8E1_12_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__65936\,
            in1 => \N__60953\,
            in2 => \N__61210\,
            in3 => \N__66753\,
            lcout => \ALU.mult_13_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_486_c_RNIPJD0I5_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58987\,
            in1 => \N__35252\,
            in2 => \_gnd_net_\,
            in3 => \N__51334\,
            lcout => OPEN,
            ltout => \ALU.mult_486_c_RNIPJD0IZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_4_c_RNI2R6596_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67065\,
            in2 => \N__34019\,
            in3 => \N__59369\,
            lcout => \ALU.addsub_cry_4_c_RNI2RZ0Z6596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5S4HI_5_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100110010100"
        )
    port map (
            in0 => \N__34011\,
            in1 => \N__74882\,
            in2 => \N__63302\,
            in3 => \N__59602\,
            lcout => \ALU.log_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICGRJG_1_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65522\,
            in2 => \_gnd_net_\,
            in3 => \N__55953\,
            lcout => \ALU.d_RNICGRJGZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_4_c_RNI5L6IQA_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34177\,
            in1 => \N__35594\,
            in2 => \_gnd_net_\,
            in3 => \N__33965\,
            lcout => \ALU.addsub_cry_4_c_RNI5L6IQAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBVMTL_5_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59601\,
            in2 => \_gnd_net_\,
            in3 => \N__68729\,
            lcout => \ALU.d_RNIBVMTLZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7ATTC1_8_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__65717\,
            in1 => \N__62820\,
            in2 => \N__62000\,
            in3 => \N__66629\,
            lcout => \ALU.mult_9_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIVMDLO_5_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59600\,
            in2 => \_gnd_net_\,
            in3 => \N__65716\,
            lcout => \ALU.d_RNIVMDLOZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9QA4D1_1_0_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__65718\,
            in1 => \N__60585\,
            in2 => \N__65564\,
            in3 => \N__66630\,
            lcout => \ALU.N_806_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNILV28R1_15_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__68727\,
            in1 => \N__65720\,
            in2 => \N__63670\,
            in3 => \N__66579\,
            lcout => \ALU.N_1030\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9QA4D1_0_0_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__66580\,
            in1 => \N__60575\,
            in2 => \N__65827\,
            in3 => \N__65527\,
            lcout => \ALU.rshift_3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIF6GEF1_12_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__60954\,
            in1 => \N__68721\,
            in2 => \N__65928\,
            in3 => \N__61170\,
            lcout => \ALU.c_RNIF6GEF1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN3QUB1_2_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__66175\,
            in1 => \N__65719\,
            in2 => \N__60205\,
            in3 => \N__66577\,
            lcout => \ALU.mult_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISLOMK_1_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__34095\,
            in1 => \N__34681\,
            in2 => \N__53301\,
            in3 => \N__34066\,
            lcout => \ALU.status_19_0\,
            ltout => \ALU.status_19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_95_c_RNO_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \N__60133\,
            in1 => \N__66174\,
            in2 => \N__34049\,
            in3 => \N__66581\,
            lcout => \ALU.mult_95_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID4IDO_0_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__66578\,
            in1 => \N__60574\,
            in2 => \_gnd_net_\,
            in3 => \N__65526\,
            lcout => \ALU.N_765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_388_c_RNIBULDP3_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101110"
        )
    port map (
            in0 => \N__34034\,
            in1 => \N__70184\,
            in2 => \N__59050\,
            in3 => \N__47936\,
            lcout => \ALU.mult_388_c_RNIBULDPZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_2_c_RNIUFTGN3_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__57231\,
            in1 => \N__59936\,
            in2 => \N__46508\,
            in3 => \N__67064\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_2_c_RNIUFTGNZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_388_c_RNIEAAJH7_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34133\,
            in2 => \N__34022\,
            in3 => \N__34253\,
            lcout => \ALU.mult_388_c_RNIEAAJHZ0Z7\,
            ltout => \ALU.mult_388_c_RNIEAAJHZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_388_c_RNIPGN6Q7_0_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__34241\,
            in1 => \N__57384\,
            in2 => \N__34247\,
            in3 => \N__69998\,
            lcout => \ALU.mult_388_c_RNIPGN6Q7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_388_c_RNIPGN6Q7_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__69999\,
            in1 => \N__34242\,
            in2 => \N__57405\,
            in3 => \N__34187\,
            lcout => \ALU.mult_388_c_RNIPGN6QZ0Z7\,
            ltout => \ALU.mult_388_c_RNIPGN6QZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_3_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__58740\,
            in1 => \_gnd_net_\,
            in2 => \N__34181\,
            in3 => \N__58665\,
            lcout => \ALU.aZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73145\,
            ce => \N__71189\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_d_s_5_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__59009\,
            in1 => \_gnd_net_\,
            in2 => \N__67115\,
            in3 => \N__70186\,
            lcout => \ALU.a_15_d_sZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a32_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__70185\,
            in1 => \N__67060\,
            in2 => \_gnd_net_\,
            in3 => \N__59005\,
            lcout => \ALU.aZ0Z32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_5_c_RNI6ET5D3_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__70089\,
            in1 => \N__59001\,
            in2 => \N__34157\,
            in3 => \N__34142\,
            lcout => \ALU.mult_5_c_RNI6ET5DZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_d_s_3_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__67052\,
            in1 => \_gnd_net_\,
            in2 => \N__59049\,
            in3 => \N__70090\,
            lcout => \ALU.a_15_d_sZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_1_c_RNI8FKPL3_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__57227\,
            in1 => \N__60290\,
            in2 => \N__43164\,
            in3 => \N__67053\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_1_c_RNI8FKPLZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_1_c_RNIJP8K37_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34132\,
            in2 => \N__34121\,
            in3 => \N__34118\,
            lcout => \ALU.addsub_cry_1_c_RNIJP8KZ0Z37\,
            ltout => \ALU.addsub_cry_1_c_RNIJP8KZ0Z37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_1_c_RNIICPEC7_0_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__57372\,
            in1 => \N__70000\,
            in2 => \N__34280\,
            in3 => \N__43574\,
            lcout => \ALU.addsub_cry_1_c_RNIICPEC7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_1_c_RNIICPEC7_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__43573\,
            in1 => \N__57371\,
            in2 => \N__70011\,
            in3 => \N__34277\,
            lcout => \ALU.addsub_cry_1_c_RNIICPECZ0Z7\,
            ltout => \ALU.addsub_cry_1_c_RNIICPECZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_2_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39603\,
            in2 => \N__34271\,
            in3 => \N__39514\,
            lcout => \ALU.aZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73150\,
            ce => \N__71213\,
            sr => \_gnd_net_\
        );

    \ALU.un1_operation_5_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__67051\,
            in1 => \_gnd_net_\,
            in2 => \N__59048\,
            in3 => \N__70088\,
            lcout => \ALU.un1_operation_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIG7RU_9_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__43553\,
            in1 => \N__47277\,
            in2 => \N__46211\,
            in3 => \N__54284\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI0FTR1_9_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__72353\,
            in1 => \N__46667\,
            in2 => \N__34268\,
            in3 => \N__47194\,
            lcout => \ALU.N_1094\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIID111_9_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__48833\,
            in1 => \N__47276\,
            in2 => \N__48991\,
            in3 => \N__54285\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4R9G1_9_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__37960\,
            in1 => \N__52745\,
            in2 => \N__34265\,
            in3 => \N__47195\,
            lcout => OPEN,
            ltout => \ALU.N_1142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7ELL3_9_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34262\,
            in2 => \N__34256\,
            in3 => \N__54134\,
            lcout => \aluOut_9\,
            ltout => \aluOut_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIN8NU4_9_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__53231\,
            in1 => \N__49577\,
            in2 => \N__34406\,
            in3 => \N__50153\,
            lcout => \ALU.d_RNIN8NU4Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIVLMT_2_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__36361\,
            in1 => \N__39415\,
            in2 => \N__35631\,
            in3 => \N__36317\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2RL91_2_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__34392\,
            in1 => \N__36073\,
            in2 => \N__34355\,
            in3 => \N__54234\,
            lcout => \ALU.N_1135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNITFGR_2_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__36362\,
            in1 => \N__34348\,
            in2 => \N__34333\,
            in3 => \N__36318\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNITB6K1_2_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__43896\,
            in1 => \N__35550\,
            in2 => \N__34310\,
            in3 => \N__35872\,
            lcout => OPEN,
            ltout => \ALU.N_1087_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2BA73_2_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54112\,
            in2 => \N__34307\,
            in3 => \N__34304\,
            lcout => \aluOut_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_RNIBQE03_0_0_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__54111\,
            in1 => \N__50152\,
            in2 => \N__49578\,
            in3 => \N__34297\,
            lcout => \CONTROL.operand1_ne_RNIBQE03_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m217_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000001000"
        )
    port map (
            in0 => \N__77315\,
            in1 => \N__75879\,
            in2 => \N__78863\,
            in3 => \N__78063\,
            lcout => \PROM.ROMDATA.m217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m238_am_1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111010100011"
        )
    port map (
            in0 => \N__75880\,
            in1 => \N__78849\,
            in2 => \N__76634\,
            in3 => \N__77316\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m238_am_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m238_am_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000100000"
        )
    port map (
            in0 => \N__78850\,
            in1 => \N__75881\,
            in2 => \N__34442\,
            in3 => \N__78064\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m238_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m244_ns_1_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010011101"
        )
    port map (
            in0 => \N__72693\,
            in1 => \N__45092\,
            in2 => \N__34439\,
            in3 => \N__45539\,
            lcout => \PROM.ROMDATA.m244_ns_1\,
            ltout => \PROM.ROMDATA.m244_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m244_ns_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001110"
        )
    port map (
            in0 => \N__72689\,
            in1 => \N__79420\,
            in2 => \N__34436\,
            in3 => \N__54355\,
            lcout => \PROM_ROMDATA_dintern_8ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_fast_ne_1_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100111010"
        )
    port map (
            in0 => \N__54358\,
            in1 => \N__34428\,
            in2 => \N__79489\,
            in3 => \N__72692\,
            lcout => \aluOperand1_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_fast_ne_1C_net\,
            ce => \N__36241\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_1_rep1_ne_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100001110"
        )
    port map (
            in0 => \N__72690\,
            in1 => \N__79421\,
            in2 => \N__34432\,
            in3 => \N__54356\,
            lcout => \aluOperand1_1_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_fast_ne_1C_net\,
            ce => \N__36241\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_1_rep2_ne_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100111010"
        )
    port map (
            in0 => \N__54357\,
            in1 => \N__34427\,
            in2 => \N__79488\,
            in3 => \N__72691\,
            lcout => \aluOperand1_1_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_fast_ne_1C_net\,
            ce => \N__36241\,
            sr => \_gnd_net_\
        );

    \ALU.b_RNI1OMT_3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__39866\,
            in1 => \N__36363\,
            in2 => \N__44242\,
            in3 => \N__36324\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6VL91_3_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__37850\,
            in1 => \N__58606\,
            in2 => \N__34409\,
            in3 => \N__54249\,
            lcout => \ALU.N_1136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIVHGR_3_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__37822\,
            in1 => \N__36364\,
            in2 => \N__37801\,
            in3 => \N__36325\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI1G6K1_3_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__37768\,
            in1 => \N__37741\,
            in2 => \N__34601\,
            in3 => \N__43897\,
            lcout => OPEN,
            ltout => \ALU.N_1088_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAJA73_3_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34598\,
            in2 => \N__34592\,
            in3 => \N__54041\,
            lcout => \aluOut_3\,
            ltout => \aluOut_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIH16V3_2_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49501\,
            in2 => \N__34589\,
            in3 => \N__50157\,
            lcout => \busState_1_RNIH16V3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI48EA1_13_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__57166\,
            in1 => \N__34559\,
            in2 => \N__52487\,
            in3 => \N__43919\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIAAVQ1_13_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__52358\,
            in1 => \N__67352\,
            in2 => \N__34571\,
            in3 => \N__47201\,
            lcout => \ALU.N_1098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI6GQI1_13_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__51548\,
            in1 => \N__34558\,
            in2 => \N__57638\,
            in3 => \N__43918\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIEQNB2_13_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__57892\,
            in1 => \N__65056\,
            in2 => \N__34511\,
            in3 => \N__47202\,
            lcout => OPEN,
            ltout => \ALU.N_1146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIR85G4_13_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34508\,
            in2 => \N__34502\,
            in3 => \N__54059\,
            lcout => \aluOut_13\,
            ltout => \aluOut_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIKLFS7_0_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__34499\,
            in1 => \N__34490\,
            in2 => \N__34460\,
            in3 => \N__49806\,
            lcout => \CONTROL.bus_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI4KP71_1_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__48409\,
            in1 => \N__46925\,
            in2 => \N__49177\,
            in3 => \N__46812\,
            lcout => \ALU.operand2_6_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJMOB4_0_1_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__53964\,
            in1 => \N__34652\,
            in2 => \N__71435\,
            in3 => \N__34645\,
            lcout => OPEN,
            ltout => \ALU.c_RNIJMOB4_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID42JA_1_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34661\,
            in2 => \N__34688\,
            in3 => \N__34634\,
            lcout => \ALU.d_RNID42JAZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7NGR1_1_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__46815\,
            in1 => \N__52166\,
            in2 => \N__37516\,
            in3 => \N__34667\,
            lcout => \ALU.N_1246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI2EJ51_1_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__37238\,
            in1 => \N__46926\,
            in2 => \N__46358\,
            in3 => \N__46813\,
            lcout => OPEN,
            ltout => \ALU.operand2_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3B472_1_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__46814\,
            in1 => \N__48943\,
            in2 => \N__34655\,
            in3 => \N__46463\,
            lcout => \ALU.N_1198\,
            ltout => \ALU.N_1198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJMOB4_1_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__34646\,
            in1 => \N__71380\,
            in2 => \N__34637\,
            in3 => \N__53963\,
            lcout => \ALU.c_RNIJMOB4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI7FBMHV_7_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__34628\,
            in1 => \N__34856\,
            in2 => \N__36263\,
            in3 => \N__34823\,
            lcout => \CONTROL.N_5\,
            ltout => \CONTROL.N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNIPON8992_3_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__34807\,
            in1 => \N__34739\,
            in2 => \N__34622\,
            in3 => \N__34816\,
            lcout => \CONTROL.addrstackptr_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI0GOJ_2_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34847\,
            in1 => \N__54814\,
            in2 => \_gnd_net_\,
            in3 => \N__49948\,
            lcout => \CONTROL.N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI060HM91_2_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38437\,
            in1 => \N__57792\,
            in2 => \N__60743\,
            in3 => \N__41923\,
            lcout => \CONTROL.un1_addrstackptr_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIO2O5VB_2_7_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111111"
        )
    port map (
            in0 => \N__41489\,
            in1 => \N__54661\,
            in2 => \N__71852\,
            in3 => \N__44712\,
            lcout => \CONTROL.g0_3_i_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_3_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__34817\,
            in1 => \N__34808\,
            in2 => \N__34753\,
            in3 => \N__34778\,
            lcout => \CONTROL.addrstackptrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.addrstackptr_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_ne_1_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__42196\,
            in1 => \N__71831\,
            in2 => \N__72305\,
            in3 => \N__54587\,
            lcout => \aluOperation_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluOperation_ne_1C_net\,
            ce => \N__38125\,
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState101_3_0_a2_308_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__72297\,
            in1 => \N__71830\,
            in2 => \_gnd_net_\,
            in3 => \N__42195\,
            lcout => \CONTROL.N_83_0\,
            ltout => \CONTROL.N_83_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m28_0_120_i_i_4_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__41258\,
            in1 => \N__34883\,
            in2 => \N__34715\,
            in3 => \N__34706\,
            lcout => \CONTROL.m28_0_120_i_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_12_i_o2_6_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__40958\,
            in1 => \N__41602\,
            in2 => \_gnd_net_\,
            in3 => \N__41257\,
            lcout => \CONTROL.N_75_0\,
            ltout => \CONTROL.N_75_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m38_i_2_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__41603\,
            in1 => \N__36797\,
            in2 => \N__34700\,
            in3 => \N__44749\,
            lcout => \CONTROL.m38_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_3_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__44748\,
            in1 => \N__44663\,
            in2 => \N__41696\,
            in3 => \N__44840\,
            lcout => \CONTROL.N_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState103_0_a2_2_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011111"
        )
    port map (
            in0 => \N__72264\,
            in1 => \_gnd_net_\,
            in2 => \N__42220\,
            in3 => \N__55444\,
            lcout => \CONTROL.N_219\,
            ltout => \CONTROL.N_219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m11_0_a2_1_0_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__54586\,
            in1 => \N__44662\,
            in2 => \N__34877\,
            in3 => \N__44839\,
            lcout => \CONTROL.N_350_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m38_i_a2_1_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__41650\,
            in1 => \N__38579\,
            in2 => \_gnd_net_\,
            in3 => \N__72293\,
            lcout => \CONTROL.N_246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m11_0_a2_2_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__54656\,
            in1 => \N__44866\,
            in2 => \N__44759\,
            in3 => \N__44703\,
            lcout => \CONTROL.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_0_0_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__41651\,
            in1 => \N__38580\,
            in2 => \_gnd_net_\,
            in3 => \N__55466\,
            lcout => OPEN,
            ltout => \CONTROL.m28_0_120_i_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNO_1_1_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38606\,
            in2 => \N__34874\,
            in3 => \N__54707\,
            lcout => OPEN,
            ltout => \CONTROL.busState_1_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNO_0_1_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__38624\,
            in1 => \_gnd_net_\,
            in2 => \N__34871\,
            in3 => \N__38633\,
            lcout => \CONTROL.busState_1_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_7_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101111111"
        )
    port map (
            in0 => \N__55465\,
            in1 => \N__42216\,
            in2 => \N__72317\,
            in3 => \N__54654\,
            lcout => \CONTROL.g0_3_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramWrite_5_m9_0_a2_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38581\,
            in2 => \_gnd_net_\,
            in3 => \N__35182\,
            lcout => \CONTROL.N_345\,
            ltout => \CONTROL.N_345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramWrite_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__35156\,
            in1 => \N__35134\,
            in2 => \N__35120\,
            in3 => \N__36817\,
            lcout => \ramWrite\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramWriteC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState114_1_0_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__54653\,
            in1 => \N__47043\,
            in2 => \N__36833\,
            in3 => \N__47015\,
            lcout => \CONTROL.un1_busState114_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_12_i_a2_6_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__44882\,
            in1 => \N__54652\,
            in2 => \N__41433\,
            in3 => \N__44700\,
            lcout => \CONTROL.N_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_10_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.dout_reto_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m1_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110101"
        )
    port map (
            in0 => \N__64747\,
            in1 => \N__64711\,
            in2 => \N__73661\,
            in3 => \N__77282\,
            lcout => \PROM.ROMDATA.m1\,
            ltout => \PROM.ROMDATA.m1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m312_am_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__78855\,
            in1 => \N__73857\,
            in2 => \N__34886\,
            in3 => \N__75906\,
            lcout => \PROM.ROMDATA.m312_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m298_am_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__75905\,
            in1 => \N__64877\,
            in2 => \N__73873\,
            in3 => \N__78856\,
            lcout => \PROM.ROMDATA.m298_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m2_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000100010"
        )
    port map (
            in0 => \N__77283\,
            in1 => \N__64748\,
            in2 => \N__64715\,
            in3 => \N__73627\,
            lcout => \PROM.ROMDATA.m2\,
            ltout => \PROM.ROMDATA.m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m451_am_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__75904\,
            in1 => \N__78996\,
            in2 => \N__35333\,
            in3 => \N__78854\,
            lcout => \PROM.ROMDATA.m451_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0OE8H_6_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__39086\,
            in1 => \N__62571\,
            in2 => \N__39044\,
            in3 => \N__53302\,
            lcout => \ALU.mult_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIG7E8H_4_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__39087\,
            in1 => \N__59898\,
            in2 => \N__39045\,
            in3 => \N__53303\,
            lcout => \ALU.mult_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_18_cry_0_c_RNO_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__39088\,
            in1 => \N__60624\,
            in2 => \N__39046\,
            in3 => \N__53304\,
            lcout => \ALU.status_18_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIDBF7E1_14_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__60994\,
            in1 => \N__65989\,
            in2 => \N__63854\,
            in3 => \N__66715\,
            lcout => \ALU.lshift_3_ns_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_391_c_RNIEC73T4_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__59124\,
            in1 => \N__35306\,
            in2 => \N__35297\,
            in3 => \N__51491\,
            lcout => \ALU.mult_391_c_RNIEC73TZ0Z4\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \ALU.mult_25_c4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_486_c_RNINTF5V4_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36986\,
            in2 => \N__35267\,
            in3 => \N__35246\,
            lcout => \ALU.mult_5\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c4\,
            carryout => \ALU.mult_25_c5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_489_c_RNIPFFTA9_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35243\,
            in2 => \N__35237\,
            in3 => \N__35216\,
            lcout => \ALU.mult_6\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c5\,
            carryout => \ALU.mult_25_c6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_492_c_RNION7CK6_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35213\,
            in2 => \N__35207\,
            in3 => \N__35192\,
            lcout => \ALU.mult_7\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c6\,
            carryout => \ALU.mult_25_c7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_495_c_RNI449047_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35516\,
            in2 => \N__35504\,
            in3 => \N__35495\,
            lcout => \ALU.mult_25_8\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c7\,
            carryout => \ALU.mult_25_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_498_c_RNI5QTSS6_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35492\,
            in2 => \N__35480\,
            in3 => \N__35471\,
            lcout => \ALU.mult_25_9\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c8\,
            carryout => \ALU.mult_25_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_501_c_RNII3J3L6_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35468\,
            in2 => \N__35462\,
            in3 => \N__35447\,
            lcout => \ALU.mult_25_10\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c9\,
            carryout => \ALU.mult_25_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_504_c_RNIA6C9P6_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35444\,
            in2 => \N__35432\,
            in3 => \N__35423\,
            lcout => \ALU.mult_25_11\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c10\,
            carryout => \ALU.mult_25_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_507_c_RNIBABOO6_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35420\,
            in2 => \N__35408\,
            in3 => \N__35399\,
            lcout => \ALU.mult_25_12\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \ALU.mult_25_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_510_c_RNIHTE1V6_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35396\,
            in2 => \N__35384\,
            in3 => \N__35375\,
            lcout => \ALU.mult_25_13\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c12\,
            carryout => \ALU.mult_25_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_513_c_RNIGEHOR6_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35372\,
            in2 => \N__35360\,
            in3 => \N__35351\,
            lcout => \ALU.mult_25_14\,
            ltout => OPEN,
            carryin => \ALU.mult_25_c13\,
            carryout => \ALU.mult_25_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_516_c_RNI98SKDC_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42347\,
            in1 => \N__35348\,
            in2 => \N__38894\,
            in3 => \N__35336\,
            lcout => \ALU.mult_516_c_RNI98SKDCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDR5C61_8_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__62859\,
            in1 => \N__68315\,
            in2 => \N__68908\,
            in3 => \N__61983\,
            lcout => \ALU.d_RNIDR5C61Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIUT8OG4_0_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__68845\,
            in1 => \N__48082\,
            in2 => \N__68460\,
            in3 => \N__48023\,
            lcout => \ALU.d_RNIUT8OG4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI8FSDB2_12_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__65755\,
            in1 => \N__61157\,
            in2 => \N__35588\,
            in3 => \N__61425\,
            lcout => OPEN,
            ltout => \ALU.N_646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIMNASS6_12_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__68846\,
            in1 => \N__68468\,
            in2 => \N__35576\,
            in3 => \N__39175\,
            lcout => OPEN,
            ltout => \ALU.lshift_15_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNICF0UCB_12_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__43166\,
            in1 => \N__43603\,
            in2 => \N__35573\,
            in3 => \N__68378\,
            lcout => \ALU.lshift_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINUT6P_13_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60938\,
            in2 => \_gnd_net_\,
            in3 => \N__65754\,
            lcout => \ALU.c_RNINUT6PZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_365_c_RNO_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__61156\,
            in1 => \N__65753\,
            in2 => \N__66717\,
            in3 => \N__60940\,
            lcout => \ALU.mult_365_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIS83N71_12_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__60939\,
            in1 => \N__68374\,
            in2 => \N__61194\,
            in3 => \N__68844\,
            lcout => \ALU.c_RNIS83N71Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.g_2_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39605\,
            in1 => \N__39531\,
            in2 => \_gnd_net_\,
            in3 => \N__39475\,
            lcout => g_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73140\,
            ce => \N__70994\,
            sr => \_gnd_net_\
        );

    \ALU.g_4_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57382\,
            in1 => \N__42536\,
            in2 => \_gnd_net_\,
            in3 => \N__39394\,
            lcout => g_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73140\,
            ce => \N__70994\,
            sr => \_gnd_net_\
        );

    \ALU.g_5_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57378\,
            in1 => \N__52628\,
            in2 => \_gnd_net_\,
            in3 => \N__39301\,
            lcout => g_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73140\,
            ce => \N__70994\,
            sr => \_gnd_net_\
        );

    \ALU.g_6_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43066\,
            in1 => \N__43120\,
            in2 => \_gnd_net_\,
            in3 => \N__42992\,
            lcout => g_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73140\,
            ce => \N__70994\,
            sr => \_gnd_net_\
        );

    \ALU.g_3_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__58679\,
            in1 => \N__58717\,
            in2 => \_gnd_net_\,
            in3 => \N__58816\,
            lcout => g_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73140\,
            ce => \N__70994\,
            sr => \_gnd_net_\
        );

    \ALU.g_10_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58526\,
            in1 => \N__58370\,
            in2 => \_gnd_net_\,
            in3 => \N__58284\,
            lcout => g_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73140\,
            ce => \N__70994\,
            sr => \_gnd_net_\
        );

    \ALU.g_11_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__58196\,
            in1 => \N__58110\,
            in2 => \_gnd_net_\,
            in3 => \N__58052\,
            lcout => g_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73140\,
            ce => \N__70994\,
            sr => \_gnd_net_\
        );

    \ALU.f_2_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39530\,
            in1 => \N__39607\,
            in2 => \_gnd_net_\,
            in3 => \N__39458\,
            lcout => f_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73142\,
            ce => \N__67871\,
            sr => \_gnd_net_\
        );

    \ALU.f_4_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57389\,
            in1 => \N__42547\,
            in2 => \_gnd_net_\,
            in3 => \N__39387\,
            lcout => f_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73142\,
            ce => \N__67871\,
            sr => \_gnd_net_\
        );

    \ALU.f_5_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57388\,
            in2 => \N__52636\,
            in3 => \N__39315\,
            lcout => f_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73142\,
            ce => \N__67871\,
            sr => \_gnd_net_\
        );

    \ALU.f_6_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43051\,
            in1 => \N__43119\,
            in2 => \_gnd_net_\,
            in3 => \N__42983\,
            lcout => f_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73142\,
            ce => \N__67871\,
            sr => \_gnd_net_\
        );

    \ALU.f_3_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__58739\,
            in1 => \N__58663\,
            in2 => \_gnd_net_\,
            in3 => \N__58800\,
            lcout => f_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73142\,
            ce => \N__67871\,
            sr => \_gnd_net_\
        );

    \ALU.f_10_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58494\,
            in1 => \N__58366\,
            in2 => \_gnd_net_\,
            in3 => \N__58294\,
            lcout => f_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73142\,
            ce => \N__67871\,
            sr => \_gnd_net_\
        );

    \ALU.f_11_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__58118\,
            in1 => \N__58188\,
            in2 => \_gnd_net_\,
            in3 => \N__58049\,
            lcout => f_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73142\,
            ce => \N__67871\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ZERO_LUT4_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ZERO_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_2_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39515\,
            in1 => \N__39599\,
            in2 => \_gnd_net_\,
            in3 => \N__39455\,
            lcout => \ALU.cZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73144\,
            ce => \N__71554\,
            sr => \_gnd_net_\
        );

    \ALU.c_4_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__42546\,
            in1 => \_gnd_net_\,
            in2 => \N__57383\,
            in3 => \N__39392\,
            lcout => \ALU.cZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73144\,
            ce => \N__71554\,
            sr => \_gnd_net_\
        );

    \ALU.c_5_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52612\,
            in1 => \N__39314\,
            in2 => \_gnd_net_\,
            in3 => \N__57351\,
            lcout => \ALU.cZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73144\,
            ce => \N__71554\,
            sr => \_gnd_net_\
        );

    \ALU.c_6_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43041\,
            in1 => \N__43105\,
            in2 => \_gnd_net_\,
            in3 => \N__42978\,
            lcout => \ALU.cZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73144\,
            ce => \N__71554\,
            sr => \_gnd_net_\
        );

    \ALU.c_3_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__58741\,
            in1 => \N__58664\,
            in2 => \_gnd_net_\,
            in3 => \N__58801\,
            lcout => \ALU.cZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73144\,
            ce => \N__71554\,
            sr => \_gnd_net_\
        );

    \ALU.c_10_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58495\,
            in2 => \N__58373\,
            in3 => \N__58295\,
            lcout => \ALU.cZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73144\,
            ce => \N__71554\,
            sr => \_gnd_net_\
        );

    \ALU.c_11_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__58109\,
            in1 => \N__58189\,
            in2 => \_gnd_net_\,
            in3 => \N__58051\,
            lcout => \ALU.cZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73144\,
            ce => \N__71554\,
            sr => \_gnd_net_\
        );

    \ALU.d_2_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39598\,
            in1 => \N__39517\,
            in2 => \_gnd_net_\,
            in3 => \N__39457\,
            lcout => \ALU.dZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73147\,
            ce => \N__70249\,
            sr => \_gnd_net_\
        );

    \ALU.d_4_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42548\,
            in1 => \N__57396\,
            in2 => \_gnd_net_\,
            in3 => \N__39393\,
            lcout => \ALU.dZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73147\,
            ce => \N__70249\,
            sr => \_gnd_net_\
        );

    \ALU.d_5_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__52623\,
            in1 => \_gnd_net_\,
            in2 => \N__57412\,
            in3 => \N__39321\,
            lcout => \ALU.dZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73147\,
            ce => \N__70249\,
            sr => \_gnd_net_\
        );

    \ALU.d_6_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43065\,
            in1 => \N__43118\,
            in2 => \_gnd_net_\,
            in3 => \N__42982\,
            lcout => \ALU.dZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73147\,
            ce => \N__70249\,
            sr => \_gnd_net_\
        );

    \ALU.d_3_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58752\,
            in1 => \N__58808\,
            in2 => \_gnd_net_\,
            in3 => \N__58676\,
            lcout => \ALU.dZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73147\,
            ce => \N__70249\,
            sr => \_gnd_net_\
        );

    \ALU.d_10_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58525\,
            in1 => \N__58365\,
            in2 => \_gnd_net_\,
            in3 => \N__58299\,
            lcout => \ALU.dZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73147\,
            ce => \N__70249\,
            sr => \_gnd_net_\
        );

    \ALU.d_11_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__58119\,
            in1 => \N__58190\,
            in2 => \_gnd_net_\,
            in3 => \N__58057\,
            lcout => \ALU.dZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73147\,
            ce => \N__70249\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_fast_ne_2_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__44497\,
            in1 => \N__40297\,
            in2 => \N__40925\,
            in3 => \N__79507\,
            lcout => \aluOperand2_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_fast_ne_2C_net\,
            ce => \N__40647\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_ne_2_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__40296\,
            in1 => \N__40920\,
            in2 => \N__79527\,
            in3 => \N__44498\,
            lcout => \aluOperand2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_fast_ne_2C_net\,
            ce => \N__40647\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI6DCT_11_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__57997\,
            in1 => \N__36184\,
            in2 => \_gnd_net_\,
            in3 => \N__43237\,
            lcout => \ALU.d_RNI6DCTZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNICJCT_14_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43238\,
            in1 => \N__57852\,
            in2 => \_gnd_net_\,
            in3 => \N__67783\,
            lcout => \ALU.d_RNICJCTZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_ne_0_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__72694\,
            in1 => \N__44927\,
            in2 => \N__41072\,
            in3 => \N__50720\,
            lcout => \aluOperand2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_fast_ne_2C_net\,
            ce => \N__40647\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI02EVNB_4_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36158\,
            in1 => \N__39251\,
            in2 => \_gnd_net_\,
            in3 => \N__68516\,
            lcout => \ALU.d_RNI02EVNBZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIG2L52_15_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__46684\,
            in1 => \N__36146\,
            in2 => \N__50404\,
            in3 => \N__53425\,
            lcout => \ALU.N_1212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI7F2G1_15_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__46549\,
            in1 => \N__53574\,
            in2 => \N__46237\,
            in3 => \N__53477\,
            lcout => \ALU.operand2_3_ns_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI5PJ21_15_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__46550\,
            in1 => \N__36371\,
            in2 => \N__46238\,
            in3 => \N__36326\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNID2PE1_15_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__43903\,
            in1 => \N__50400\,
            in2 => \N__36140\,
            in3 => \N__46685\,
            lcout => \ALU.N_1100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI710B1_15_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__53612\,
            in1 => \N__36370\,
            in2 => \N__53530\,
            in3 => \N__36327\,
            lcout => \ALU.dout_6_ns_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIE4B6N4_15_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__37637\,
            in1 => \N__63615\,
            in2 => \N__69168\,
            in3 => \N__50351\,
            lcout => \ALU.c_RNIE4B6N4Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_16_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__38248\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63463\,
            lcout => \CONTROL.increment28lto5_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_11_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63462\,
            in2 => \_gnd_net_\,
            in3 => \N__38249\,
            lcout => OPEN,
            ltout => \CONTROL.increment28lto5_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_a7_4_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__48468\,
            in1 => \N__40826\,
            in2 => \N__36266\,
            in3 => \N__38209\,
            lcout => \CONTROL.g0_3_i_a7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m221cf1_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001111"
        )
    port map (
            in0 => \N__36206\,
            in1 => \N__74038\,
            in2 => \N__73412\,
            in3 => \N__72688\,
            lcout => \PROM.ROMDATA.m221cf1\,
            ltout => \PROM.ROMDATA.m221cf1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m221_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45238\,
            in1 => \_gnd_net_\,
            in2 => \N__36251\,
            in3 => \N__36196\,
            lcout => \PROM_ROMDATA_dintern_7ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand1_ne_0_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36197\,
            in1 => \N__36248\,
            in2 => \_gnd_net_\,
            in3 => \N__45239\,
            lcout => \aluOperand1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand1_ne_0C_net\,
            ce => \N__36242\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m221cf0_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__74037\,
            in1 => \N__36205\,
            in2 => \N__72742\,
            in3 => \N__73433\,
            lcout => \PROM.ROMDATA.m221cf0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_7_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63461\,
            in2 => \_gnd_net_\,
            in3 => \N__38247\,
            lcout => \CONTROL.increment28lto5_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState103_0_a2_1_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__54584\,
            in1 => \N__36878\,
            in2 => \N__36397\,
            in3 => \N__41210\,
            lcout => OPEN,
            ltout => \CONTROL.N_320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState103_0_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__36452\,
            in1 => \N__36377\,
            in2 => \N__36410\,
            in3 => \N__41201\,
            lcout => \CONTROL.un1_busState103_0_0\,
            ltout => \CONTROL.un1_busState103_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_1_0_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__63030\,
            in1 => \N__36713\,
            in2 => \N__36407\,
            in3 => \N__41582\,
            lcout => \aluParams_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluParams_1_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState103_0_o2_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71820\,
            in2 => \_gnd_net_\,
            in3 => \N__44661\,
            lcout => \CONTROL.N_95_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState103_0_a2_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__54583\,
            in1 => \N__41396\,
            in2 => \N__41235\,
            in3 => \N__44871\,
            lcout => \CONTROL.N_318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNITJ3GK_12_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001101000"
        )
    port map (
            in0 => \N__56910\,
            in1 => \N__74682\,
            in2 => \N__63076\,
            in3 => \N__61151\,
            lcout => \ALU.N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNITVOEK_12_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__61152\,
            in1 => \N__63026\,
            in2 => \_gnd_net_\,
            in3 => \N__56909\,
            lcout => \ALU.c_RNITVOEKZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA7CLH_8_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001101000"
        )
    port map (
            in0 => \N__55812\,
            in1 => \N__74681\,
            in2 => \N__63075\,
            in3 => \N__61930\,
            lcout => \ALU.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_1_ne_RNO_0_1_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100010011"
        )
    port map (
            in0 => \N__44656\,
            in1 => \N__74815\,
            in2 => \N__41357\,
            in3 => \N__44869\,
            lcout => OPEN,
            ltout => \CONTROL.N_340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_1_ne_1_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001011"
        )
    port map (
            in0 => \N__44870\,
            in1 => \N__54585\,
            in2 => \N__36533\,
            in3 => \N__44657\,
            lcout => \aluParams_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluParams_1_ne_1C_net\,
            ce => \N__36530\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAJ1KH_8_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__61931\,
            in1 => \N__63022\,
            in2 => \_gnd_net_\,
            in3 => \N__55811\,
            lcout => \ALU.d_RNIAJ1KHZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState114_2_0_0_x1_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__44867\,
            in1 => \N__41305\,
            in2 => \N__54651\,
            in3 => \N__44654\,
            lcout => \CONTROL.un1_busState114_2_0_0_xZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState114_2_0_0_x0_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111010"
        )
    port map (
            in0 => \N__44655\,
            in1 => \N__54579\,
            in2 => \N__41356\,
            in3 => \N__44868\,
            lcout => OPEN,
            ltout => \CONTROL.un1_busState114_2_0_0_xZ0Z0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState114_2_0_0_ns_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71745\,
            in2 => \N__36518\,
            in3 => \N__36515\,
            lcout => \CONTROL.un1_busState114_2_0_0_0\,
            ltout => \CONTROL.un1_busState114_2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState114_2_0_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__47033\,
            in1 => \N__46984\,
            in2 => \N__36509\,
            in3 => \N__54580\,
            lcout => \CONTROL.un1_busState114_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_4_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__38127\,
            in1 => \N__41203\,
            in2 => \N__69885\,
            in3 => \N__41394\,
            lcout => \aluOperation_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluOperation_4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_1_sqmuxa_0_a2_2_0_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__55451\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54539\,
            lcout => \CONTROL.aluReadBus_1_sqmuxa_0_a2_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState96_1_i_2_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001010001"
        )
    port map (
            in0 => \N__40963\,
            in1 => \N__41575\,
            in2 => \N__36487\,
            in3 => \N__41202\,
            lcout => \CONTROL.N_48_0\,
            ltout => \CONTROL.N_48_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_2_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__41576\,
            in1 => \N__70054\,
            in2 => \N__36635\,
            in3 => \N__36632\,
            lcout => \aluOperation_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluOperation_4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_RNO_0_2_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__54541\,
            in1 => \N__41393\,
            in2 => \N__71853\,
            in3 => \N__44650\,
            lcout => \CONTROL.un1_controlWord_14_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluReadBus_RNO_1_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110011"
        )
    port map (
            in0 => \N__41392\,
            in1 => \N__38699\,
            in2 => \N__36625\,
            in3 => \N__38623\,
            lcout => \CONTROL.un1_busState97_1_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment_5_0__m6_i_0_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__54540\,
            in1 => \N__42221\,
            in2 => \N__72316\,
            in3 => \N__55452\,
            lcout => \CONTROL.un1_busState114_2_0_o2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNII6GE_7_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__73319\,
            in1 => \N__36566\,
            in2 => \_gnd_net_\,
            in3 => \N__45145\,
            lcout => OPEN,
            ltout => \CONTROL.N_422_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNII9UU_7_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__36554\,
            in1 => \_gnd_net_\,
            in2 => \N__36539\,
            in3 => \N__73677\,
            lcout => \progRomAddress_7\,
            ltout => \progRomAddress_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_2_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__72263\,
            in1 => \N__41008\,
            in2 => \N__36536\,
            in3 => \N__45766\,
            lcout => \CONTROL.ctrlOut_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_2C_net\,
            ce => \N__44396\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m90_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110110011100"
        )
    port map (
            in0 => \N__77862\,
            in1 => \N__78779\,
            in2 => \N__75984\,
            in3 => \N__77174\,
            lcout => \PROM.ROMDATA.m90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_3dflt_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001010"
        )
    port map (
            in0 => \N__72262\,
            in1 => \N__41834\,
            in2 => \N__72606\,
            in3 => \N__64397\,
            lcout => \controlWord_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIE2GE_5_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45146\,
            in1 => \N__45662\,
            in2 => \_gnd_net_\,
            in3 => \N__41723\,
            lcout => OPEN,
            ltout => \CONTROL.N_420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIC3UU_5_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__73679\,
            in1 => \_gnd_net_\,
            in2 => \N__36746\,
            in3 => \N__41771\,
            lcout => \CONTROL.programCounter_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_1_cry_0_c_RNO_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47407\,
            in1 => \N__73678\,
            in2 => \_gnd_net_\,
            in3 => \N__50962\,
            lcout => \CONTROL.programCounter_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_1_RNO_0_0_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__41108\,
            in1 => \N__41424\,
            in2 => \N__72626\,
            in3 => \N__41810\,
            lcout => \CONTROL.N_105_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI1CMQ_12_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__42070\,
            in1 => \N__36755\,
            in2 => \_gnd_net_\,
            in3 => \N__38753\,
            lcout => \CONTROL.N_427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m177_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47309\,
            in1 => \N__72503\,
            in2 => \_gnd_net_\,
            in3 => \N__64900\,
            lcout => \PROM_ROMDATA_dintern_5ro\,
            ltout => \PROM_ROMDATA_dintern_5ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState111_0_202_a2_0_o2_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__71802\,
            in1 => \_gnd_net_\,
            in2 => \N__36692\,
            in3 => \N__72226\,
            lcout => \CONTROL.N_80_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_0_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__72227\,
            in1 => \N__42208\,
            in2 => \_gnd_net_\,
            in3 => \N__71803\,
            lcout => \CONTROL.N_98_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_1_i_3_1_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000001000"
        )
    port map (
            in0 => \N__71804\,
            in1 => \N__54573\,
            in2 => \N__42235\,
            in3 => \N__44639\,
            lcout => \CONTROL.g0_1_i_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState114_1_0_a2_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__44640\,
            in1 => \N__42212\,
            in2 => \_gnd_net_\,
            in3 => \N__71805\,
            lcout => OPEN,
            ltout => \CONTROL.N_209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState114_1_0_0_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36879\,
            in2 => \N__36836\,
            in3 => \N__54574\,
            lcout => \CONTROL.un1_busState114_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m38_i_a2_0_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__41423\,
            in1 => \N__54632\,
            in2 => \N__38582\,
            in3 => \N__44884\,
            lcout => OPEN,
            ltout => \CONTROL.N_349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m38_i_1_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36788\,
            in2 => \N__36824\,
            in3 => \N__36813\,
            lcout => \CONTROL.m38_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m38_i_a2_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110101"
        )
    port map (
            in0 => \N__51065\,
            in1 => \N__45343\,
            in2 => \N__72698\,
            in3 => \N__44883\,
            lcout => \CONTROL.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_12_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36782\,
            lcout => \CONTROL.programCounter_1_reto_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState_0_sqmuxa_i_a2_2_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41655\,
            in2 => \_gnd_net_\,
            in3 => \N__38567\,
            lcout => \CONTROL.N_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_1dflt_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__72608\,
            in1 => \N__51064\,
            in2 => \N__45344\,
            in3 => \N__72224\,
            lcout => \controlWord_1\,
            ltout => \controlWord_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState_1_sqmuxa_i_a2_1_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__72225\,
            in1 => \_gnd_net_\,
            in2 => \N__36749\,
            in3 => \N__38566\,
            lcout => \CONTROL.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState97_i_i_o2_0_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001001"
        )
    port map (
            in0 => \N__41580\,
            in1 => \N__41256\,
            in2 => \N__40962\,
            in3 => \N__41434\,
            lcout => \CONTROL.N_136_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m506_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__74487\,
            in1 => \N__76600\,
            in2 => \N__65029\,
            in3 => \N__75907\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m508_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__79503\,
            in2 => \N__36953\,
            in3 => \N__79897\,
            lcout => \PROM.ROMDATA.N_571_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI64MA6_0_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__71471\,
            in1 => \N__36932\,
            in2 => \_gnd_net_\,
            in3 => \N__37874\,
            lcout => \ALU.d_RNI64MA6Z0Z_0\,
            ltout => \ALU.d_RNI64MA6Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_21_0_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39040\,
            in2 => \N__36899\,
            in3 => \N__53298\,
            lcout => OPEN,
            ltout => \ALU.log_1_3_ns_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_17_0_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63254\,
            in2 => \N__36896\,
            in3 => \N__60616\,
            lcout => OPEN,
            ltout => \ALU.log_1_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_11_0_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010010101100"
        )
    port map (
            in0 => \N__63255\,
            in1 => \N__74895\,
            in2 => \N__36893\,
            in3 => \N__66716\,
            lcout => OPEN,
            ltout => \ALU.log_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_5_0_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__63256\,
            in1 => \N__37193\,
            in2 => \N__36890\,
            in3 => \N__37373\,
            lcout => OPEN,
            ltout => \ALU.status_8_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_2_0_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__48176\,
            in1 => \N__51458\,
            in2 => \N__36887\,
            in3 => \N__51203\,
            lcout => \ALU.status_RNO_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_365_c_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37052\,
            in2 => \N__37385\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \ALU.mult_13_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_365_c_RNINK1M82_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37040\,
            in2 => \N__37028\,
            in3 => \N__37016\,
            lcout => \ALU.mult_13_14\,
            ltout => OPEN,
            carryin => \ALU.mult_13_c13\,
            carryout => \ALU.mult_13_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_371_c_RNIAJLO71_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37013\,
            in2 => \_gnd_net_\,
            in3 => \N__37004\,
            lcout => \ALU.mult_13_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_365_c_RNI8ALO96_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__63835\,
            in1 => \N__38821\,
            in2 => \N__42377\,
            in3 => \N__66714\,
            lcout => \ALU.mult_365_c_RNI8ALOZ0Z96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIL4PC21_6_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__62232\,
            in1 => \N__55958\,
            in2 => \N__56130\,
            in3 => \N__62558\,
            lcout => \ALU.d_RNIL4PC21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9VEDD1_4_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__59620\,
            in1 => \N__65990\,
            in2 => \N__59912\,
            in3 => \N__66713\,
            lcout => \ALU.mult_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_546_c_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48790\,
            in2 => \N__48772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \ALU.mult_29_c8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_546_c_RNIUNL1A8_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36980\,
            in2 => \N__36968\,
            in3 => \N__36959\,
            lcout => \ALU.mult_9\,
            ltout => OPEN,
            carryin => \ALU.mult_29_c8\,
            carryout => \ALU.mult_29_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_549_c_RNIV9413G_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42437\,
            in2 => \N__42463\,
            in3 => \N__36956\,
            lcout => \ALU.mult_10\,
            ltout => OPEN,
            carryin => \ALU.mult_29_c9\,
            carryout => \ALU.mult_29_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_552_c_RNIK1H74A_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42416\,
            in2 => \N__37172\,
            in3 => \N__37163\,
            lcout => \ALU.mult_11\,
            ltout => OPEN,
            carryin => \ALU.mult_29_c10\,
            carryout => \ALU.mult_29_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_555_c_RNI9QLKVH_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38957\,
            in2 => \N__38977\,
            in3 => \N__37160\,
            lcout => \ALU.mult_12\,
            ltout => OPEN,
            carryin => \ALU.mult_29_c11\,
            carryout => \ALU.mult_29_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_558_c_RNIN3VB2C_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37157\,
            in2 => \N__38930\,
            in3 => \N__37151\,
            lcout => \ALU.mult_13\,
            ltout => OPEN,
            carryin => \ALU.mult_29_c12\,
            carryout => \ALU.mult_29_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_561_c_RNIL4S0IG_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37148\,
            in2 => \N__38909\,
            in3 => \N__37142\,
            lcout => \ALU.mult_14\,
            ltout => OPEN,
            carryin => \ALU.mult_29_c13\,
            carryout => \ALU.mult_29_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_564_c_RNIRTQTDC_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37139\,
            in2 => \_gnd_net_\,
            in3 => \N__37133\,
            lcout => \ALU.mult_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_9_c_RNI0ALKH7_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110100011"
        )
    port map (
            in0 => \N__39244\,
            in1 => \N__61505\,
            in2 => \N__66902\,
            in3 => \N__68459\,
            lcout => \ALU.a_15_am_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_549_c_RNIB6TIDG_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__59044\,
            in1 => \N__37130\,
            in2 => \_gnd_net_\,
            in3 => \N__37094\,
            lcout => OPEN,
            ltout => \ALU.mult_549_c_RNIB6TIDGZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_549_c_RNIE7260O_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101001010100"
        )
    port map (
            in0 => \N__66901\,
            in1 => \N__67047\,
            in2 => \N__37088\,
            in3 => \N__37085\,
            lcout => \ALU.mult_549_c_RNIE7260OZ0\,
            ltout => \ALU.mult_549_c_RNIE7260OZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_10_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__58455\,
            in1 => \_gnd_net_\,
            in2 => \N__37079\,
            in3 => \N__58343\,
            lcout => \ALU.aZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73141\,
            ce => \N__71211\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_m3_s_13_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59043\,
            in2 => \_gnd_net_\,
            in3 => \N__59295\,
            lcout => \ALU.a_15_m3_sZ0Z_13\,
            ltout => \ALU.a_15_m3_sZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_s_13_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__67046\,
            in1 => \_gnd_net_\,
            in2 => \N__37244\,
            in3 => \_gnd_net_\,
            lcout => \ALU.a_15_sZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a32_0_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59042\,
            in2 => \_gnd_net_\,
            in3 => \N__67045\,
            lcout => \ALU.a32Z0Z_0\,
            ltout => \ALU.a32Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_1_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__59296\,
            in1 => \N__52205\,
            in2 => \N__37241\,
            in3 => \N__69014\,
            lcout => \ALU.aZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73141\,
            ce => \N__71211\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNICUA7B5_0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011111101"
        )
    port map (
            in0 => \N__70168\,
            in1 => \N__37178\,
            in2 => \N__59139\,
            in3 => \N__40175\,
            lcout => OPEN,
            ltout => \ALU.d_RNICUA7B5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_0_c_RNI43EE86_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67044\,
            in2 => \N__37208\,
            in3 => \N__60326\,
            lcout => \ALU.a_15_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIL3JT71_0_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__56929\,
            in1 => \N__65556\,
            in2 => \N__56804\,
            in3 => \N__60602\,
            lcout => \ALU.d_RNIL3JT71Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5A8KO_1_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010001000"
        )
    port map (
            in0 => \N__74853\,
            in1 => \N__65551\,
            in2 => \_gnd_net_\,
            in3 => \N__65926\,
            lcout => \ALU.N_556\,
            ltout => \ALU.N_556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3MGBH1_1_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__70167\,
            in1 => \N__63291\,
            in2 => \N__37181\,
            in3 => \N__37369\,
            lcout => \ALU.d_RNI3MGBH1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_39_c_RNO_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__60965\,
            in1 => \N__56787\,
            in2 => \N__61216\,
            in3 => \N__56928\,
            lcout => \ALU.status_17_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_365_c_RNO_0_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60964\,
            in2 => \_gnd_net_\,
            in3 => \N__66582\,
            lcout => \ALU.mult_365_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5A8KO_0_1_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111101110"
        )
    port map (
            in0 => \N__74854\,
            in1 => \N__65552\,
            in2 => \_gnd_net_\,
            in3 => \N__65927\,
            lcout => \ALU.N_572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_10_c_RNISV0175_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69944\,
            in1 => \N__61276\,
            in2 => \N__69679\,
            in3 => \N__37292\,
            lcout => \ALU.a_15_am_rn_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_552_c_RNI70R9DA_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37341\,
            in1 => \N__69645\,
            in2 => \_gnd_net_\,
            in3 => \N__37304\,
            lcout => \ALU.mult_552_c_RNI70R9DAZ0\,
            ltout => \ALU.mult_552_c_RNI70R9DAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_552_c_RNIOT7VLF_0_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__37285\,
            in1 => \N__43037\,
            in2 => \N__37295\,
            in3 => \N__37532\,
            lcout => \ALU.mult_552_c_RNIOT7VLFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIP0VNF4_15_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__43184\,
            in1 => \N__68464\,
            in2 => \N__42872\,
            in3 => \N__68809\,
            lcout => \ALU.rshift_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_552_c_RNIOT7VLF_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011011100"
        )
    port map (
            in0 => \N__37531\,
            in1 => \N__43038\,
            in2 => \N__37286\,
            in3 => \N__37274\,
            lcout => \ALU.mult_552_c_RNIOT7VLFZ0\,
            ltout => \ALU.mult_552_c_RNIOT7VLFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_11_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58165\,
            in2 => \N__37268\,
            in3 => \N__58111\,
            lcout => \ALU.aZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73146\,
            ce => \N__71216\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_am_sn_11_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__69641\,
            in1 => \N__67043\,
            in2 => \_gnd_net_\,
            in3 => \N__69943\,
            lcout => \ALU.a_15_am_snZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_1_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__59298\,
            in1 => \N__52223\,
            in2 => \N__69666\,
            in3 => \N__69013\,
            lcout => h_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73151\,
            ce => \N__69453\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_s_11_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__69646\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59297\,
            lcout => \ALU.a_15_sZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_489_c_RNIGEUL1A_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__67042\,
            in1 => \N__62345\,
            in2 => \_gnd_net_\,
            in3 => \N__37478\,
            lcout => \ALU.mult_489_c_RNIGEUL1AZ0\,
            ltout => \ALU.mult_489_c_RNIGEUL1AZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_489_c_RNIPGBQMC_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__69647\,
            in1 => \N__52678\,
            in2 => \N__37466\,
            in3 => \N__63319\,
            lcout => \ALU.mult_489_c_RNIPGBQMCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_489_c_RNIPGBQMC_0_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__52679\,
            in1 => \N__63320\,
            in2 => \N__69680\,
            in3 => \N__37463\,
            lcout => OPEN,
            ltout => \ALU.mult_489_c_RNIPGBQMCZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_489_c_RNI1J3GCU_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__39209\,
            in1 => \_gnd_net_\,
            in2 => \N__37457\,
            in3 => \N__37454\,
            lcout => \ALU.mult_489_c_RNI1J3GCUZ0\,
            ltout => \ALU.mult_489_c_RNI1J3GCUZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_6_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43039\,
            in2 => \N__37448\,
            in3 => \N__43104\,
            lcout => h_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73151\,
            ce => \N__69453\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4HL061_0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__66685\,
            in1 => \N__60365\,
            in2 => \N__67204\,
            in3 => \N__60566\,
            lcout => \ALU.d_RNI4HL061Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA4TMK_0_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110111010100"
        )
    port map (
            in0 => \N__50541\,
            in1 => \N__60572\,
            in2 => \N__74832\,
            in3 => \N__66686\,
            lcout => OPEN,
            ltout => \ALU.a_15_m2_d_d_ns_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4D6E01_0_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__59282\,
            in1 => \N__50542\,
            in2 => \N__37691\,
            in3 => \N__37659\,
            lcout => OPEN,
            ltout => \ALU.d_RNI4D6E01Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQQ9O83_0_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__59328\,
            in1 => \N__37636\,
            in2 => \N__37604\,
            in3 => \N__60573\,
            lcout => OPEN,
            ltout => \ALU.d_RNIQQ9O83Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINUGCF4_0_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69651\,
            in2 => \N__37601\,
            in3 => \N__37598\,
            lcout => \ALU.d_RNINUGCF4Z0Z_0\,
            ltout => \ALU.d_RNINUGCF4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_0_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__69160\,
            in1 => \N__69627\,
            in2 => \N__37592\,
            in3 => \N__52055\,
            lcout => \ALU.aZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73154\,
            ce => \N__71193\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_s_15_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__59281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__70139\,
            lcout => \ALU.a_15_m2_sZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI933S_0_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46325\,
            in1 => \N__37579\,
            in2 => \_gnd_net_\,
            in3 => \N__53572\,
            lcout => \ALU.e_RNI933SZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_0_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__52080\,
            in1 => \N__69161\,
            in2 => \N__69689\,
            in3 => \N__52054\,
            lcout => h_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73160\,
            ce => \N__69450\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0G5D_0_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43983\,
            in1 => \N__37548\,
            in2 => \_gnd_net_\,
            in3 => \N__51967\,
            lcout => \ALU.d_RNI0G5DZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIDFF01_0_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48901\,
            in1 => \N__46429\,
            in2 => \_gnd_net_\,
            in3 => \N__53573\,
            lcout => OPEN,
            ltout => \ALU.c_RNIDFF01Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNITEVO2_0_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__53859\,
            in1 => \N__37898\,
            in2 => \N__37892\,
            in3 => \N__53410\,
            lcout => \ALU.operand2_7_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIS3PO_0_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49131\,
            in1 => \N__48380\,
            in2 => \_gnd_net_\,
            in3 => \N__43982\,
            lcout => OPEN,
            ltout => \ALU.b_RNIS3POZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITCRC4_0_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__53860\,
            in1 => \N__37889\,
            in2 => \N__37883\,
            in3 => \N__37880\,
            lcout => \ALU.operand2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNICGJM_9_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46207\,
            in1 => \N__43552\,
            in2 => \_gnd_net_\,
            in3 => \N__43981\,
            lcout => \ALU.e_RNICGJMZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI3E5B1_3_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__39862\,
            in1 => \N__53570\,
            in2 => \N__44235\,
            in3 => \N__53466\,
            lcout => OPEN,
            ltout => \ALU.operand2_6_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI8SEV1_3_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__37843\,
            in1 => \N__58602\,
            in2 => \N__37829\,
            in3 => \N__53405\,
            lcout => \ALU.N_1248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI18V81_3_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__37826\,
            in1 => \N__53571\,
            in2 => \N__37802\,
            in3 => \N__53467\,
            lcout => OPEN,
            ltout => \ALU.operand2_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI4G2B2_3_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__37769\,
            in1 => \N__37737\,
            in2 => \N__37694\,
            in3 => \N__53406\,
            lcout => OPEN,
            ltout => \ALU.N_1200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGMEO4_3_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53861\,
            in2 => \N__38093\,
            in3 => \N__38090\,
            lcout => OPEN,
            ltout => \ALU.d_RNIGMEO4Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2CUG6_3_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71400\,
            in2 => \N__38084\,
            in3 => \N__38081\,
            lcout => \ALU.d_RNI2CUG6Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNI4KOJ_4_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38027\,
            in1 => \N__55334\,
            in2 => \_gnd_net_\,
            in3 => \N__50168\,
            lcout => \CONTROL.N_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_9_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__66845\,
            in1 => \N__58498\,
            in2 => \N__52889\,
            in3 => \N__52808\,
            lcout => h_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73181\,
            ce => \N__69454\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKKNJ_9_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43242\,
            in1 => \N__37941\,
            in2 => \_gnd_net_\,
            in3 => \N__52744\,
            lcout => \ALU.d_RNIKKNJZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIG8BV_9_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48832\,
            in1 => \N__48981\,
            in2 => \_gnd_net_\,
            in3 => \N__43243\,
            lcout => \ALU.b_RNIG8BVZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI65HE2_9_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__37925\,
            in1 => \N__43415\,
            in2 => \N__53940\,
            in3 => \N__46782\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIECHF4_9_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__37916\,
            in1 => \N__53898\,
            in2 => \N__37910\,
            in3 => \N__37907\,
            lcout => OPEN,
            ltout => \ALU.operand2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4K8P6_9_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100111"
        )
    port map (
            in0 => \N__71401\,
            in1 => \N__40400\,
            in2 => \N__37901\,
            in3 => \N__49825\,
            lcout => \ALU.combOperand2_0_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_0_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__56573\,
            in1 => \N__38303\,
            in2 => \N__38285\,
            in3 => \N__48425\,
            lcout => \aluStatus_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_0_0_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100110011"
        )
    port map (
            in0 => \N__56532\,
            in1 => \N__48463\,
            in2 => \N__71504\,
            in3 => \N__69318\,
            lcout => \ALU.status_e_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69317\,
            in2 => \_gnd_net_\,
            in3 => \N__71500\,
            lcout => \ALU.un1_a41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment28lto5_1_1_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63459\,
            in2 => \_gnd_net_\,
            in3 => \N__38264\,
            lcout => OPEN,
            ltout => \CONTROL.increment28lto5_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment28lto5_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001010101"
        )
    port map (
            in0 => \N__72252\,
            in1 => \N__41018\,
            in2 => \N__38276\,
            in3 => \N__38160\,
            lcout => \CONTROL.N_361_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_14_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63460\,
            in2 => \_gnd_net_\,
            in3 => \N__38265\,
            lcout => OPEN,
            ltout => \CONTROL.increment28lto5_1_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_2_i_a7_3_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__38205\,
            in1 => \N__40819\,
            in2 => \N__38219\,
            in3 => \N__48453\,
            lcout => \CONTROL.g0_2_i_a7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment28lto5_1_2_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100110011001"
        )
    port map (
            in0 => \N__72251\,
            in1 => \N__40818\,
            in2 => \N__48464\,
            in3 => \N__38204\,
            lcout => \CONTROL.increment28lto5_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_ne_5_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__44660\,
            in1 => \N__54582\,
            in2 => \N__41397\,
            in3 => \N__44901\,
            lcout => \aluOperation_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluOperation_ne_5C_net\,
            ce => \N__38126\,
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState96_1_i_i_a2_0_1_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__41689\,
            in1 => \N__38584\,
            in2 => \_gnd_net_\,
            in3 => \N__55456\,
            lcout => \CONTROL.un1_busState96_1_i_i_a2_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState96_1_i_i_o2_0_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__55455\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44658\,
            lcout => \CONTROL.N_140_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_6dflt_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72273\,
            in2 => \_gnd_net_\,
            in3 => \N__55454\,
            lcout => \controlWord_6\,
            ltout => \controlWord_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState96_1_i_i_a2_1_1_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__38583\,
            in1 => \N__41688\,
            in2 => \N__38354\,
            in3 => \N__44659\,
            lcout => OPEN,
            ltout => \CONTROL.un1_busState96_1_i_i_a2_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState96_1_i_i_0_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100111111"
        )
    port map (
            in0 => \N__38351\,
            in1 => \N__54719\,
            in2 => \N__38345\,
            in3 => \N__54581\,
            lcout => OPEN,
            ltout => \CONTROL.un1_busState96_1_i_iZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI41SBR02_7_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__38330\,
            in1 => \N__38342\,
            in2 => \N__38336\,
            in3 => \N__41117\,
            lcout => \CONTROL.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_5dflt_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__47305\,
            in1 => \N__72272\,
            in2 => \N__72607\,
            in3 => \N__64904\,
            lcout => \controlWord_5\,
            ltout => \controlWord_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState96_1_i_i_o2_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100100011"
        )
    port map (
            in0 => \N__44635\,
            in1 => \N__54571\,
            in2 => \N__38333\,
            in3 => \N__44862\,
            lcout => \CONTROL.N_134_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState_0_sqmuxa_i_a2_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__44769\,
            in1 => \N__44863\,
            in2 => \N__38528\,
            in3 => \N__44636\,
            lcout => \CONTROL.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_2_i_a7_2_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__53627\,
            in1 => \N__45401\,
            in2 => \N__45479\,
            in3 => \N__54572\,
            lcout => \CONTROL.g0_2_i_a7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_22_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__54569\,
            in1 => \N__71758\,
            in2 => \_gnd_net_\,
            in3 => \N__44634\,
            lcout => \CONTROL.N_133_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m126_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__72504\,
            in1 => \N__64396\,
            in2 => \_gnd_net_\,
            in3 => \N__41833\,
            lcout => \PROM_ROMDATA_dintern_3ro\,
            ltout => \PROM_ROMDATA_dintern_3ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_6_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54568\,
            in2 => \N__38504\,
            in3 => \N__44632\,
            lcout => \CONTROL.N_133_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIO2O5VB_1_7_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__44633\,
            in1 => \N__41464\,
            in2 => \N__71819\,
            in3 => \N__54570\,
            lcout => \CONTROL.g0_3_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIO2O5VB_7_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111111"
        )
    port map (
            in0 => \N__41463\,
            in1 => \N__54575\,
            in2 => \N__71821\,
            in3 => \N__44649\,
            lcout => OPEN,
            ltout => \CONTROL.g0_2_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI7FBMHV_0_7_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__38486\,
            in1 => \N__38477\,
            in2 => \N__38471\,
            in3 => \N__42149\,
            lcout => \CONTROL.N_5_0\,
            ltout => \CONTROL.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNIJQC4JV_1_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111110101"
        )
    port map (
            in0 => \N__38468\,
            in1 => \N__38444\,
            in2 => \N__38375\,
            in3 => \N__57820\,
            lcout => \CONTROL.g0_12_1\,
            ltout => \CONTROL.g0_12_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNITKBIQ83_2_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011110001011"
        )
    port map (
            in0 => \N__60682\,
            in1 => \N__38734\,
            in2 => \N__38372\,
            in3 => \N__41958\,
            lcout => \CONTROL.addrstackptr_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_2dflt_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__41100\,
            in1 => \N__72261\,
            in2 => \N__72672\,
            in3 => \N__41805\,
            lcout => \controlWord_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_4dflt_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__72260\,
            in1 => \N__72563\,
            in2 => \N__54389\,
            in3 => \N__74138\,
            lcout => \controlWord_4\,
            ltout => \controlWord_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIQ59BL4_7_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__41101\,
            in1 => \N__72618\,
            in2 => \N__38738\,
            in3 => \N__41806\,
            lcout => \CONTROL.N_249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_2_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001001110110001"
        )
    port map (
            in0 => \N__38735\,
            in1 => \N__38723\,
            in2 => \N__60701\,
            in3 => \N__41959\,
            lcout => \CONTROL.addrstackptrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.addrstackptr_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m28_0_120_i_i_0_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110111"
        )
    port map (
            in0 => \N__41233\,
            in1 => \N__38678\,
            in2 => \N__38810\,
            in3 => \N__38644\,
            lcout => \CONTROL.m28_0_120_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState97_1_0_a2_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001100"
        )
    port map (
            in0 => \N__44865\,
            in1 => \N__41581\,
            in2 => \N__41415\,
            in3 => \N__41234\,
            lcout => \CONTROL.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m28_0_120_i_i_a2_2_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__54543\,
            in1 => \N__41372\,
            in2 => \N__41670\,
            in3 => \N__44864\,
            lcout => \CONTROL.N_338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment_5_0__m6_i_x2_0_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001011010"
        )
    port map (
            in0 => \N__44638\,
            in1 => \_gnd_net_\,
            in2 => \N__41416\,
            in3 => \N__71806\,
            lcout => \CONTROL.N_114_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m42_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__72511\,
            in1 => \N__74011\,
            in2 => \N__45554\,
            in3 => \N__47702\,
            lcout => \PROM_ROMDATA_dintern_0ro\,
            ltout => \PROM_ROMDATA_dintern_0ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState_0_sqmuxa_i_a2_0_0_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38531\,
            in3 => \N__54542\,
            lcout => \CONTROL.un1_busState_0_sqmuxa_i_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m28_0_120_i_i_o2_1_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__55453\,
            in1 => \N__41371\,
            in2 => \N__72320\,
            in3 => \N__44637\,
            lcout => \CONTROL.N_304_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m433_ns_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38744\,
            in1 => \N__47798\,
            in2 => \_gnd_net_\,
            in3 => \N__79845\,
            lcout => \PROM.ROMDATA.m433_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m294_bm_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__78838\,
            in1 => \N__74129\,
            in2 => \N__75967\,
            in3 => \N__78059\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m294_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m294_ns_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41081\,
            in1 => \_gnd_net_\,
            in2 => \N__38780\,
            in3 => \N__76592\,
            lcout => \PROM.ROMDATA.m294_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m31_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__78836\,
            in1 => \N__78055\,
            in2 => \_gnd_net_\,
            in3 => \N__77280\,
            lcout => \PROM.ROMDATA.m31\,
            ltout => \PROM.ROMDATA.m31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m353_bm_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41819\,
            in2 => \N__38777\,
            in3 => \N__75846\,
            lcout => \PROM.ROMDATA.m353_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_12_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38774\,
            lcout => \CONTROL.dout_reto_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73234\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m391_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001000001"
        )
    port map (
            in0 => \N__77281\,
            in1 => \N__75847\,
            in2 => \N__78071\,
            in3 => \N__78837\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m391_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m433_bm_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76591\,
            in2 => \N__38747\,
            in3 => \N__74246\,
            lcout => \PROM.ROMDATA.m433_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m382_ns_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__79342\,
            in1 => \N__42137\,
            in2 => \N__47363\,
            in3 => \N__42119\,
            lcout => \PROM.ROMDATA.m382_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI27KBD_0_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100111100"
        )
    port map (
            in0 => \N__39024\,
            in1 => \N__39089\,
            in2 => \N__63275\,
            in3 => \N__53292\,
            lcout => \ALU.d_RNI27KBDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA3Q1H_0_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000010000"
        )
    port map (
            in0 => \N__53294\,
            in1 => \N__39100\,
            in2 => \N__60627\,
            in3 => \N__39025\,
            lcout => \ALU.N_794_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI6USD6_2_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__49604\,
            in1 => \N__50218\,
            in2 => \N__60626\,
            in3 => \N__38855\,
            lcout => \N_225_0\,
            ltout => \N_225_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNISBUGH_14_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__63843\,
            in1 => \N__39091\,
            in2 => \N__38834\,
            in3 => \N__53295\,
            lcout => OPEN,
            ltout => \ALU.mult_15_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_371_c_RNIHIRFF5_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__39200\,
            in1 => \N__38831\,
            in2 => \N__38825\,
            in3 => \N__38822\,
            lcout => \ALU.mult_23_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIIRAJH_10_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011000000"
        )
    port map (
            in0 => \N__39023\,
            in1 => \N__39090\,
            in2 => \N__61715\,
            in3 => \N__53293\,
            lcout => \ALU.mult_11_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIA5S1H_8_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010100000"
        )
    port map (
            in0 => \N__39095\,
            in1 => \N__39027\,
            in2 => \N__62022\,
            in3 => \N__53296\,
            lcout => \ALU.mult_9_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIRFM5I_11_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011101000"
        )
    port map (
            in0 => \N__63112\,
            in1 => \N__61466\,
            in2 => \N__74894\,
            in3 => \N__57046\,
            lcout => \ALU.log_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIKU5GD1_0_14_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__66027\,
            in1 => \N__63669\,
            in2 => \N__63853\,
            in3 => \N__66764\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIR6KVA2_12_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__61012\,
            in1 => \N__61203\,
            in2 => \N__39104\,
            in3 => \N__66028\,
            lcout => \ALU.N_647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI5O9IH_12_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010100000"
        )
    port map (
            in0 => \N__39096\,
            in1 => \N__39026\,
            in2 => \N__61217\,
            in3 => \N__53297\,
            lcout => \ALU.mult_13_12\,
            ltout => \ALU.mult_13_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_467_c_RNICRDK6B_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__38981\,
            in1 => \_gnd_net_\,
            in2 => \N__38960\,
            in3 => \N__42400\,
            lcout => \ALU.mult_467_c_RNICRDK6BZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_526_c_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42401\,
            in2 => \N__38951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \ALU.mult_27_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_526_c_RNIHBG235_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42386\,
            in2 => \N__38942\,
            in3 => \N__38921\,
            lcout => \ALU.mult_27_13\,
            ltout => OPEN,
            carryin => \ALU.mult_27_c12\,
            carryout => \ALU.mult_27_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_529_c_RNIM6FVL9_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42370\,
            in2 => \N__38918\,
            in3 => \N__38900\,
            lcout => \ALU.mult_27_14\,
            ltout => OPEN,
            carryin => \ALU.mult_27_c13\,
            carryout => \ALU.mult_27_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_27_c14_THRU_LUT4_0_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38897\,
            lcout => \ALU.mult_27_c14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_546_c_RNIG1E6I8_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59144\,
            in2 => \N__38882\,
            in3 => \N__40353\,
            lcout => \ALU.mult_546_c_RNIG1E6IZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINMQ0E1_10_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011000000"
        )
    port map (
            in0 => \N__61465\,
            in1 => \N__65935\,
            in2 => \N__61716\,
            in3 => \N__66697\,
            lcout => \ALU.mult_11_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_558_c_RNIB3E8DC_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__59145\,
            in1 => \N__39656\,
            in2 => \_gnd_net_\,
            in3 => \N__39182\,
            lcout => \ALU.mult_558_c_RNIB3E8DCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFCNKL_9_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62818\,
            in2 => \_gnd_net_\,
            in3 => \N__68841\,
            lcout => \ALU.d_RNIFCNKLZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIG61LG_9_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__62819\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68439\,
            lcout => \ALU.d_RNIG61LGZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIULN025_0_2_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__68440\,
            in1 => \N__43599\,
            in2 => \N__43165\,
            in3 => \N__68842\,
            lcout => \ALU.d_RNIULN025_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIULN025_2_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110101"
        )
    port map (
            in0 => \N__68843\,
            in1 => \N__43160\,
            in2 => \N__43604\,
            in3 => \N__68441\,
            lcout => OPEN,
            ltout => \ALU.d_RNIULN025Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPTFHMD_2_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39176\,
            in2 => \N__39152\,
            in3 => \N__39149\,
            lcout => OPEN,
            ltout => \ALU.lshift_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIO0KOKE_10_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__70191\,
            in2 => \N__39143\,
            in3 => \N__51296\,
            lcout => \ALU.c_RNIO0KOKEZ0Z_10\,
            ltout => \ALU.c_RNIO0KOKEZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_10_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58456\,
            in2 => \N__39140\,
            in3 => \N__58283\,
            lcout => \ALU.bZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73143\,
            ce => \N__67938\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNI8TL4B6_12_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__42787\,
            in1 => \N__42794\,
            in2 => \_gnd_net_\,
            in3 => \N__39188\,
            lcout => \ALU.N_1025\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIHOSI72_12_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__65903\,
            in1 => \N__42811\,
            in2 => \_gnd_net_\,
            in3 => \N__42788\,
            lcout => OPEN,
            ltout => \ALU.N_965_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFHCRU4_2_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__39233\,
            in1 => \_gnd_net_\,
            in2 => \N__39212\,
            in3 => \N__68920\,
            lcout => \ALU.d_RNIFHCRU4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBN2FN8_11_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__70187\,
            in1 => \N__51322\,
            in2 => \_gnd_net_\,
            in3 => \N__42821\,
            lcout => \ALU.c_RNIBN2FN8Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINMQ0E1_0_10_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__61439\,
            in1 => \N__65904\,
            in2 => \N__61717\,
            in3 => \N__66699\,
            lcout => \ALU.lshift_3_ns_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIKU5GD1_14_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__66698\,
            in1 => \N__63644\,
            in2 => \N__63842\,
            in3 => \N__65902\,
            lcout => \ALU.mult_15_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINT9PO2_10_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__68919\,
            in1 => \N__42810\,
            in2 => \N__62656\,
            in3 => \N__65905\,
            lcout => \ALU.c_RNINT9PO2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI61KC1_13_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51541\,
            in1 => \N__57631\,
            in2 => \_gnd_net_\,
            in3 => \N__43295\,
            lcout => \ALU.b_RNI61KC1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAHCT_13_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43294\,
            in1 => \N__57891\,
            in2 => \_gnd_net_\,
            in3 => \N__65060\,
            lcout => \ALU.d_RNIAHCTZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI890L_13_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52350\,
            in1 => \N__67348\,
            in2 => \_gnd_net_\,
            in3 => \N__43293\,
            lcout => \ALU.c_RNI890LZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI4P741_13_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43296\,
            in1 => \N__52477\,
            in2 => \_gnd_net_\,
            in3 => \N__57170\,
            lcout => OPEN,
            ltout => \ALU.a_RNI4P741Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNILN2L2_13_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__39698\,
            in1 => \N__53951\,
            in2 => \N__39692\,
            in3 => \N__46811\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9K0D5_13_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__53952\,
            in1 => \N__39689\,
            in2 => \N__39683\,
            in3 => \N__39680\,
            lcout => \ALU.operand2_13\,
            ltout => \ALU.operand2_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINGV4G_13_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39652\,
            in2 => \N__39614\,
            in3 => \N__71467\,
            lcout => \ALU.N_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJAJOO_10_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__61697\,
            in1 => \N__62811\,
            in2 => \_gnd_net_\,
            in3 => \N__66721\,
            lcout => \ALU.N_837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_2_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39606\,
            in1 => \N__39535\,
            in2 => \_gnd_net_\,
            in3 => \N__39468\,
            lcout => \ALU.bZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73155\,
            ce => \N__67943\,
            sr => \_gnd_net_\
        );

    \ALU.b_4_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42529\,
            in1 => \N__57350\,
            in2 => \_gnd_net_\,
            in3 => \N__39395\,
            lcout => \ALU.bZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73155\,
            ce => \N__67943\,
            sr => \_gnd_net_\
        );

    \ALU.b_5_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57349\,
            in1 => \N__52619\,
            in2 => \_gnd_net_\,
            in3 => \N__39320\,
            lcout => \ALU.bZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73155\,
            ce => \N__67943\,
            sr => \_gnd_net_\
        );

    \ALU.b_6_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43040\,
            in1 => \N__43086\,
            in2 => \_gnd_net_\,
            in3 => \N__42977\,
            lcout => \ALU.bZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73155\,
            ce => \N__67943\,
            sr => \_gnd_net_\
        );

    \ALU.b_3_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__58812\,
            in1 => \N__58745\,
            in2 => \_gnd_net_\,
            in3 => \N__58678\,
            lcout => \ALU.bZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73155\,
            ce => \N__67943\,
            sr => \_gnd_net_\
        );

    \ALU.b_11_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__58184\,
            in1 => \N__58108\,
            in2 => \_gnd_net_\,
            in3 => \N__58050\,
            lcout => \ALU.bZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73155\,
            ce => \N__67943\,
            sr => \_gnd_net_\
        );

    \ALU.b_12_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67757\,
            in2 => \N__67622\,
            in3 => \N__67691\,
            lcout => \ALU.bZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73155\,
            ce => \N__67943\,
            sr => \_gnd_net_\
        );

    \CONTROL.g3_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__53720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53668\,
            lcout => \CONTROL.gZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDC6LJ1_2_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__65957\,
            in1 => \N__39764\,
            in2 => \_gnd_net_\,
            in3 => \N__68515\,
            lcout => \ALU.lshift_15_0_1\,
            ltout => \ALU.lshift_15_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNITNPJL2_14_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__39732\,
            in1 => \N__69928\,
            in2 => \N__39707\,
            in3 => \N__39704\,
            lcout => \ALU.a_15_m0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI6KIQO_14_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001010000"
        )
    port map (
            in0 => \N__63802\,
            in1 => \N__63668\,
            in2 => \N__69965\,
            in3 => \N__66682\,
            lcout => \ALU.a_15_m0_sx_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI34ECO_9_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62764\,
            in2 => \_gnd_net_\,
            in3 => \N__65955\,
            lcout => \ALU.d_RNI34ECOZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9QA4D1_0_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010001000"
        )
    port map (
            in0 => \N__65958\,
            in1 => \N__60568\,
            in2 => \N__65575\,
            in3 => \N__66683\,
            lcout => OPEN,
            ltout => \ALU.mult_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI05SGP3_0_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__59066\,
            in1 => \N__40184\,
            in2 => \N__40178\,
            in3 => \N__47986\,
            lcout => \ALU.a_15_m3_d_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJOQE21_0_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__65569\,
            in1 => \N__60567\,
            in2 => \N__56141\,
            in3 => \N__55875\,
            lcout => \ALU.d_RNIJOQE21Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_293_c_RNO_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__66684\,
            in1 => \N__62765\,
            in2 => \N__61982\,
            in3 => \N__65956\,
            lcout => \ALU.mult_293_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI8KVQ_5_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40134\,
            in1 => \N__40090\,
            in2 => \_gnd_net_\,
            in3 => \N__43974\,
            lcout => \ALU.c_RNI8KVQZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNI48JM_5_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43975\,
            in1 => \N__40069\,
            in2 => \_gnd_net_\,
            in3 => \N__40043\,
            lcout => OPEN,
            ltout => \ALU.e_RNI48JMZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNILHDD2_5_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__53887\,
            in1 => \N__40013\,
            in2 => \N__40007\,
            in3 => \N__46779\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBAG34_5_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__40196\,
            in1 => \N__39905\,
            in2 => \N__40004\,
            in3 => \N__53888\,
            lcout => \ALU.operand2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI7HSP_5_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39973\,
            in1 => \_gnd_net_\,
            in2 => \N__46922\,
            in3 => \N__39922\,
            lcout => \ALU.b_RNI7HSPZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBT8E_5_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46892\,
            in2 => \N__40267\,
            in3 => \N__40219\,
            lcout => \ALU.d_RNIBT8EZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_2_rep1_ne_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__79411\,
            in1 => \N__40916\,
            in2 => \N__40298\,
            in3 => \N__44495\,
            lcout => \aluOperand2_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_2_rep1_neC_net\,
            ce => \N__40657\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_2_rep2_ne_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__44496\,
            in1 => \N__40292\,
            in2 => \N__40924\,
            in3 => \N__79412\,
            lcout => \aluOperand2_2_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_2_rep1_neC_net\,
            ce => \N__40657\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m407_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__74492\,
            in1 => \N__76583\,
            in2 => \N__45805\,
            in3 => \N__75815\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m418_ns_1_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__79879\,
            in1 => \N__40796\,
            in2 => \N__40190\,
            in3 => \N__72727\,
            lcout => \PROM.ROMDATA.m418_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m134_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__78851\,
            in1 => \N__78050\,
            in2 => \_gnd_net_\,
            in3 => \N__77312\,
            lcout => \PROM.ROMDATA.m134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_fast_ne_1_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__79880\,
            in1 => \N__40800\,
            in2 => \N__79495\,
            in3 => \N__72729\,
            lcout => \aluOperand2_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_fast_ne_1C_net\,
            ce => \N__40658\,
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_1_rep1_ne_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__72728\,
            in1 => \N__79433\,
            in2 => \N__40802\,
            in3 => \N__79882\,
            lcout => \aluOperand2_1_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_fast_ne_1C_net\,
            ce => \N__40658\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m488_ns_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100011000"
        )
    port map (
            in0 => \N__77313\,
            in1 => \N__74087\,
            in2 => \N__78070\,
            in3 => \N__78852\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m488_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m500_ns_1_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__64298\,
            in1 => \N__79432\,
            in2 => \N__40187\,
            in3 => \N__79878\,
            lcout => \PROM.ROMDATA.m500_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.operand2_ne_1_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__79881\,
            in1 => \N__40801\,
            in2 => \N__79496\,
            in3 => \N__72730\,
            lcout => \aluOperand2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.operand2_fast_ne_1C_net\,
            ce => \N__40658\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJP1AE_0_9_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__40601\,
            in1 => \N__40541\,
            in2 => \N__40499\,
            in3 => \N__40513\,
            lcout => \ALU.combOperand2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI27JA5_1_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__50156\,
            in1 => \N__40498\,
            in2 => \N__62886\,
            in3 => \N__50342\,
            lcout => \CONTROL.N_202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_RNIEUOJ_9_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40463\,
            in1 => \N__40309\,
            in2 => \_gnd_net_\,
            in3 => \N__50154\,
            lcout => OPEN,
            ltout => \CONTROL.N_170_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIDRGO1_2_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__50155\,
            in1 => \N__40433\,
            in2 => \N__40403\,
            in3 => \N__49575\,
            lcout => \N_186\,
            ltout => \N_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNILFVQ7_0_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__49576\,
            in1 => \N__40394\,
            in2 => \N__40388\,
            in3 => \N__49818\,
            lcout => bus_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_9_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__72300\,
            in1 => \N__72380\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.ctrlOut_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_9C_net\,
            ce => \N__44398\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m284_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__50759\,
            in1 => \N__43714\,
            in2 => \N__79861\,
            in3 => \N__78956\,
            lcout => \PROM.ROMDATA.m284\,
            ltout => \PROM.ROMDATA.m284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_12dflt_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__79298\,
            in1 => \N__40913\,
            in2 => \N__40832\,
            in3 => \N__44478\,
            lcout => \controlWord_12\,
            ltout => \controlWord_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment28lto5_0_ns_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40775\,
            in2 => \N__40829\,
            in3 => \N__40769\,
            lcout => \CONTROL.increment28lto5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m273_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__78955\,
            in1 => \N__75619\,
            in2 => \N__76619\,
            in3 => \N__78753\,
            lcout => \PROM.ROMDATA.m273\,
            ltout => \PROM.ROMDATA.m273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m276_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__72683\,
            in1 => \N__79297\,
            in2 => \N__40781\,
            in3 => \N__79783\,
            lcout => \PROM_ROMDATA_dintern_11ro\,
            ltout => \PROM_ROMDATA_dintern_11ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment28lto5_0_x1_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__72249\,
            in1 => \N__40750\,
            in2 => \N__40778\,
            in3 => \N__56656\,
            lcout => \CONTROL.increment28lto5_0_xZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment28lto5_0_x0_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__40749\,
            in1 => \N__72250\,
            in2 => \_gnd_net_\,
            in3 => \N__40762\,
            lcout => \CONTROL.increment28lto5_0_xZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_1_i_a6_0_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__40763\,
            in1 => \N__56657\,
            in2 => \N__40754\,
            in3 => \N__40715\,
            lcout => \CONTROL.g0_1_i_a6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_1_i_a6_1_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__53662\,
            in1 => \N__45509\,
            in2 => \N__53717\,
            in3 => \N__45392\,
            lcout => \CONTROL.g0_1_i_a6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_a7_0_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__45391\,
            in1 => \N__53705\,
            in2 => \N__45516\,
            in3 => \N__53661\,
            lcout => \CONTROL.g0_3_i_a7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m271_1_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111110101"
        )
    port map (
            in0 => \N__79210\,
            in1 => \N__47524\,
            in2 => \N__72726\,
            in3 => \N__47537\,
            lcout => \PROM.ROMDATA.m271_1\,
            ltout => \PROM.ROMDATA.m271_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m271_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__72655\,
            in1 => \N__44920\,
            in2 => \N__41057\,
            in3 => \N__50713\,
            lcout => \PROM_ROMDATA_dintern_10ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m258_ns_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__79818\,
            in1 => \N__45194\,
            in2 => \_gnd_net_\,
            in3 => \N__45356\,
            lcout => \PROM.ROMDATA.m258_ns\,
            ltout => \PROM.ROMDATA.m258_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m260_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011000110010"
        )
    port map (
            in0 => \N__72656\,
            in1 => \N__45031\,
            in2 => \N__41024\,
            in3 => \N__50470\,
            lcout => \PROM_ROMDATA_dintern_9ro\,
            ltout => \PROM_ROMDATA_dintern_9ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment28lto5_1_0_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__53704\,
            in1 => \N__45505\,
            in2 => \N__41021\,
            in3 => \N__45390\,
            lcout => \CONTROL.increment28lto5_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m404_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__79299\,
            in1 => \N__64246\,
            in2 => \N__47528\,
            in3 => \N__75708\,
            lcout => \PROM.ROMDATA.N_566_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m470_bm_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__64245\,
            in1 => \N__76470\,
            in2 => \N__69359\,
            in3 => \N__75598\,
            lcout => \PROM.ROMDATA.m470_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_RNO_0_6_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__41194\,
            in1 => \N__54766\,
            in2 => \N__40967\,
            in3 => \N__41559\,
            lcout => \CONTROL.aluOperation_12_i_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState97_i_i_o2_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__41558\,
            in1 => \N__41192\,
            in2 => \N__41395\,
            in3 => \N__44903\,
            lcout => \CONTROL.N_86_0\,
            ltout => \CONTROL.N_86_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_cnst_2_0__m38_i_m2_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__41193\,
            in1 => \_gnd_net_\,
            in2 => \N__41705\,
            in3 => \N__41697\,
            lcout => \CONTROL.N_135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m444_am_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__64870\,
            in1 => \N__78712\,
            in2 => \_gnd_net_\,
            in3 => \N__75597\,
            lcout => \PROM.ROMDATA.m444_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluParams_7_f0_163_0_o2_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54544\,
            in2 => \_gnd_net_\,
            in3 => \N__44631\,
            lcout => \CONTROL.N_74_0\,
            ltout => \CONTROL.N_74_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIUBNO8E_7_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__41476\,
            in1 => \N__41391\,
            in2 => \N__41264\,
            in3 => \N__44902\,
            lcout => OPEN,
            ltout => \CONTROL.un1_busState96_1_i_i_232_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNINU4NAR_7_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__41191\,
            in1 => \_gnd_net_\,
            in2 => \N__41120\,
            in3 => \N__47002\,
            lcout => \CONTROL.programCounter_ret_36_RNINU4NARZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_RNIT3IG_5_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45658\,
            in1 => \N__64595\,
            in2 => \_gnd_net_\,
            in3 => \N__41764\,
            lcout => \CONTROL.programCounter_ret_19_RNIT3IGZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m23_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__77865\,
            in1 => \_gnd_net_\,
            in2 => \N__78845\,
            in3 => \N__77182\,
            lcout => \PROM.ROMDATA.m23\,
            ltout => \PROM.ROMDATA.m23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m97_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001010"
        )
    port map (
            in0 => \N__73997\,
            in1 => \N__73491\,
            in2 => \N__41111\,
            in3 => \N__75852\,
            lcout => \PROM_ROMDATA_dintern_31_0__N_556_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m294_am_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001001000"
        )
    port map (
            in0 => \N__77866\,
            in1 => \N__78787\,
            in2 => \N__75968\,
            in3 => \N__77183\,
            lcout => \PROM.ROMDATA.m294_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m16_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100000000"
        )
    port map (
            in0 => \N__73572\,
            in1 => \N__73808\,
            in2 => \N__73719\,
            in3 => \N__77863\,
            lcout => \PROM.ROMDATA.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m125_e_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__79142\,
            in1 => \N__79613\,
            in2 => \N__76462\,
            in3 => \_gnd_net_\,
            lcout => m125_e,
            ltout => \m125_e_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m125_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__41846\,
            in1 => \N__50572\,
            in2 => \N__41837\,
            in3 => \N__75851\,
            lcout => \PROM.ROMDATA.N_557_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m77_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011010"
        )
    port map (
            in0 => \N__77864\,
            in1 => \_gnd_net_\,
            in2 => \N__78844\,
            in3 => \N__77181\,
            lcout => \PROM.ROMDATA.m77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m93_ns_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__54968\,
            in1 => \N__51107\,
            in2 => \N__79417\,
            in3 => \N__51047\,
            lcout => m93_ns,
            ltout => \m93_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNI257R22_7_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__74007\,
            in1 => \N__50561\,
            in2 => \N__41792\,
            in3 => \N__72695\,
            lcout => \CONTROL.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_5_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41789\,
            lcout => \CONTROL.addrstack_reto_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI4MHF_5_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41716\,
            in1 => \N__64594\,
            in2 => \_gnd_net_\,
            in3 => \N__41763\,
            lcout => \CONTROL.programCounter_ret_1_RNI4MHFZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_5_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_35_rep2_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__50872\,
            in1 => \_gnd_net_\,
            in2 => \N__50842\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL_programCounter11_reto_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_rep1_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50830\,
            in2 => \_gnd_net_\,
            in3 => \N__50871\,
            lcout => \CONTROL.un1_programCounter9_reto_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m48_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110010101"
        )
    port map (
            in0 => \N__78746\,
            in1 => \N__77995\,
            in2 => \N__75966\,
            in3 => \N__77258\,
            lcout => \PROM.ROMDATA.m48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_2_1_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101111111"
        )
    port map (
            in0 => \N__55421\,
            in1 => \N__72307\,
            in2 => \N__42262\,
            in3 => \N__54633\,
            lcout => \CONTROL.g0_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_4_2_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__72311\,
            in1 => \N__42026\,
            in2 => \_gnd_net_\,
            in3 => \N__55423\,
            lcout => \CONTROL.g0_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment_0_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__47010\,
            in1 => \N__42017\,
            in2 => \N__44713\,
            in3 => \N__47050\,
            lcout => \CONTROL.incrementZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.increment_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNIF0HGO91_7_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__60653\,
            in1 => \N__42280\,
            in2 => \N__42011\,
            in3 => \N__41976\,
            lcout => \CONTROL.g1_1\,
            ltout => \CONTROL.g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNIF61SK42_7_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__42334\,
            in1 => \N__42304\,
            in2 => \N__41888\,
            in3 => \N__41852\,
            lcout => \CONTROL.addrstackptr_N_7_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIEO2I4H_7_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001000110"
        )
    port map (
            in0 => \N__54635\,
            in1 => \N__42249\,
            in2 => \N__41864\,
            in3 => \N__47009\,
            lcout => \CONTROL.g0_i_m2_1\,
            ltout => \CONTROL.g0_i_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_7_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__42335\,
            in1 => \N__42305\,
            in2 => \N__42296\,
            in3 => \N__42293\,
            lcout => \CONTROL.addrstackptrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.increment_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_2_i_1_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111111111111"
        )
    port map (
            in0 => \N__54634\,
            in1 => \N__42248\,
            in2 => \N__72319\,
            in3 => \N__55422\,
            lcout => \CONTROL.g0_2_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m381_am_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__74410\,
            in1 => \N__76609\,
            in2 => \N__47885\,
            in3 => \N__75856\,
            lcout => \PROM.ROMDATA.m381_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m382_ns_1_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__42131\,
            in1 => \N__79341\,
            in2 => \N__47897\,
            in3 => \N__79846\,
            lcout => \PROM.ROMDATA.m382_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIHEO982_2_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__60187\,
            in1 => \N__66240\,
            in2 => \N__42113\,
            in3 => \N__66047\,
            lcout => OPEN,
            ltout => \ALU.N_858_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7RHUG5_2_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__68931\,
            in1 => \N__42575\,
            in2 => \N__42095\,
            in3 => \N__68526\,
            lcout => OPEN,
            ltout => \ALU.rshift_15_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0V48BA_2_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__68527\,
            in1 => \N__56474\,
            in2 => \N__42092\,
            in3 => \N__56491\,
            lcout => \ALU.rshift_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9VEDD1_0_4_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__59637\,
            in1 => \N__66045\,
            in2 => \N__59911\,
            in3 => \N__66768\,
            lcout => OPEN,
            ltout => \ALU.rshift_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5MBM92_6_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__66046\,
            in1 => \N__62587\,
            in2 => \N__42089\,
            in3 => \N__62233\,
            lcout => \ALU.N_862\,
            ltout => \ALU.N_862_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFVCT15_6_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56490\,
            in2 => \N__42569\,
            in3 => \N__68930\,
            lcout => OPEN,
            ltout => \ALU.N_922_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI1AHUF8_2_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52684\,
            in2 => \N__42566\,
            in3 => \N__42563\,
            lcout => \ALU.d_RNI1AHUF8Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_293_c_RNIOCJMD9_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__42464\,
            in1 => \N__42710\,
            in2 => \N__42446\,
            in3 => \_gnd_net_\,
            lcout => \ALU.mult_293_c_RNIOCJMDZ0Z9\,
            ltout => OPEN,
            carryin => \bfn_19_9_0_\,
            carryout => \ALU.mult_21_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_464_c_RNIRCBMA3_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42683\,
            in2 => \N__42425\,
            in3 => \N__42404\,
            lcout => \ALU.mult_21_11\,
            ltout => OPEN,
            carryin => \ALU.mult_21_c10\,
            carryout => \ALU.mult_21_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_467_c_RNISOO9S3_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42665\,
            in2 => \N__45902\,
            in3 => \N__42389\,
            lcout => \ALU.mult_21_12\,
            ltout => OPEN,
            carryin => \ALU.mult_21_c11\,
            carryout => \ALU.mult_21_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_470_c_RNIB61LK3_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42641\,
            in2 => \N__45869\,
            in3 => \N__42380\,
            lcout => \ALU.mult_21_13\,
            ltout => OPEN,
            carryin => \ALU.mult_21_c12\,
            carryout => \ALU.mult_21_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_473_c_RNIR822C3_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42602\,
            in2 => \N__45836\,
            in3 => \N__42359\,
            lcout => \ALU.mult_21_14\,
            ltout => OPEN,
            carryin => \ALU.mult_21_c13\,
            carryout => \ALU.mult_21_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_476_c_RNIFLP0O7_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__42854\,
            in1 => \N__42356\,
            in2 => \_gnd_net_\,
            in3 => \N__42350\,
            lcout => \ALU.mult_476_c_RNIFLP0OZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2BV762_8_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42815\,
            in1 => \N__42776\,
            in2 => \_gnd_net_\,
            in3 => \N__66026\,
            lcout => \ALU.N_866\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_293_c_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42881\,
            in2 => \N__42755\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_10_0_\,
            carryout => \ALU.mult_9_c9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_293_c_RNIKDLV62_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42740\,
            in2 => \N__42728\,
            in3 => \N__42704\,
            lcout => \ALU.mult_9_10\,
            ltout => OPEN,
            carryin => \ALU.mult_9_c9\,
            carryout => \ALU.mult_9_c10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_299_c_RNIJ4OGS1_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42701\,
            in2 => \N__42695\,
            in3 => \N__42677\,
            lcout => \ALU.mult_9_11\,
            ltout => OPEN,
            carryin => \ALU.mult_9_c10\,
            carryout => \ALU.mult_9_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_305_c_RNIVQ5JJ1_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45947\,
            in2 => \N__42674\,
            in3 => \N__42659\,
            lcout => \ALU.mult_9_12\,
            ltout => OPEN,
            carryin => \ALU.mult_9_c11\,
            carryout => \ALU.mult_9_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_311_c_RNIUDNBM1_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42848\,
            in2 => \N__42656\,
            in3 => \N__42635\,
            lcout => \ALU.mult_9_13\,
            ltout => OPEN,
            carryin => \ALU.mult_9_c12\,
            carryout => \ALU.mult_9_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_317_c_RNID87GM1_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42632\,
            in2 => \N__42617\,
            in3 => \N__42596\,
            lcout => \ALU.mult_9_14\,
            ltout => OPEN,
            carryin => \ALU.mult_9_c13\,
            carryout => \ALU.mult_9_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_323_c_RNIAA0B82_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42593\,
            in1 => \N__45821\,
            in2 => \N__45938\,
            in3 => \N__42578\,
            lcout => \ALU.mult_323_c_RNIAA0BZ0Z82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGD2441_8_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__56413\,
            in1 => \N__62871\,
            in2 => \N__62021\,
            in3 => \N__56259\,
            lcout => \ALU.d_RNIGD2441Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIOFVO52_4_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__65968\,
            in1 => \_gnd_net_\,
            in2 => \N__45740\,
            in3 => \N__48059\,
            lcout => \ALU.N_639\,
            ltout => \ALU.N_639_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFVCT15_8_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__68923\,
            in1 => \_gnd_net_\,
            in2 => \N__42842\,
            in3 => \N__46163\,
            lcout => OPEN,
            ltout => \ALU.d_RNIFVCT15Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4U6858_2_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42839\,
            in2 => \N__42824\,
            in3 => \N__68458\,
            lcout => \ALU.lshift_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIR02AP_10_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__61703\,
            in1 => \N__61460\,
            in2 => \_gnd_net_\,
            in3 => \N__66704\,
            lcout => \ALU.N_851\,
            ltout => \ALU.N_851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINT9PO2_0_10_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__65967\,
            in1 => \N__62648\,
            in2 => \N__42797\,
            in3 => \N__68922\,
            lcout => \ALU.c_RNINT9PO2_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_335_c_RNO_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__61702\,
            in1 => \N__65966\,
            in2 => \N__66773\,
            in3 => \N__61461\,
            lcout => \ALU.mult_335_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIQ12IP_12_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__66701\,
            in1 => \N__60990\,
            in2 => \_gnd_net_\,
            in3 => \N__61211\,
            lcout => \ALU.N_978\,
            ltout => \ALU.N_978_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIE08272_12_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62655\,
            in2 => \N__42779\,
            in3 => \N__66013\,
            lcout => \ALU.N_967\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIEOKO_1_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__65557\,
            in1 => \N__63150\,
            in2 => \_gnd_net_\,
            in3 => \N__42899\,
            lcout => \ALU.d_RNIIEOKOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI48CC42_2_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45724\,
            in1 => \N__47978\,
            in2 => \_gnd_net_\,
            in3 => \N__66014\,
            lcout => \ALU.N_635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI2HF0A9_8_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46052\,
            in1 => \N__42887\,
            in2 => \_gnd_net_\,
            in3 => \N__68528\,
            lcout => \ALU.rshift_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIO8DPO_14_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__63809\,
            in1 => \N__63645\,
            in2 => \_gnd_net_\,
            in3 => \N__66700\,
            lcout => \ALU.N_980\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIG8JO24_15_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__68790\,
            in1 => \N__42868\,
            in2 => \_gnd_net_\,
            in3 => \N__43183\,
            lcout => \ALU.N_1026\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_293_c_RNO_0_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62805\,
            in2 => \_gnd_net_\,
            in3 => \N__66718\,
            lcout => \ALU.mult_293_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIN266M_11_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__61434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68789\,
            lcout => \ALU.c_RNIN266MZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNITTCO62_10_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66080\,
            in2 => \N__46117\,
            in3 => \N__46066\,
            lcout => \ALU.N_867\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNID11991_15_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__63658\,
            in1 => \N__66082\,
            in2 => \_gnd_net_\,
            in3 => \N__66720\,
            lcout => \ALU.N_1011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIET09P_12_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__66719\,
            in1 => \N__61435\,
            in2 => \_gnd_net_\,
            in3 => \N__61212\,
            lcout => \ALU.N_852\,
            ltout => \ALU.N_852_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIR8GG72_12_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__53332\,
            in1 => \_gnd_net_\,
            in2 => \N__43187\,
            in3 => \N__66081\,
            lcout => \ALU.N_966\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQQRSN_2_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__65565\,
            in1 => \_gnd_net_\,
            in2 => \N__66767\,
            in3 => \N__66287\,
            lcout => \ALU.N_766\,
            ltout => \ALU.N_766_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0KELT1_2_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__66079\,
            in1 => \_gnd_net_\,
            in2 => \N__43169\,
            in3 => \N__48583\,
            lcout => \ALU.N_634\,
            ltout => \ALU.N_634_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILTB1L4_2_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43590\,
            in2 => \N__43127\,
            in3 => \N__68921\,
            lcout => OPEN,
            ltout => \ALU.N_811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIK8M6K5_6_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__70197\,
            in1 => \N__51262\,
            in2 => \N__43124\,
            in3 => \N__68529\,
            lcout => \ALU.d_RNIK8M6K5Z0Z_6\,
            ltout => \ALU.d_RNIK8M6K5Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_6_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__43055\,
            in1 => \_gnd_net_\,
            in2 => \N__42995\,
            in3 => \N__42990\,
            lcout => \ALU.aZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73161\,
            ce => \N__71199\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKRBVN_0_4_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__60237\,
            in1 => \N__59849\,
            in2 => \_gnd_net_\,
            in3 => \N__66746\,
            lcout => \ALU.N_606\,
            ltout => \ALU.N_606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIAC0J42_2_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42908\,
            in2 => \N__42902\,
            in3 => \N__66077\,
            lcout => \ALU.N_636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDBRC52_4_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__66078\,
            in1 => \N__48672\,
            in2 => \_gnd_net_\,
            in3 => \N__43610\,
            lcout => \ALU.N_638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m0_am_2_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__43531\,
            in1 => \N__49830\,
            in2 => \_gnd_net_\,
            in3 => \N__43507\,
            lcout => \ALU.a_15_m0_amZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGE45L7_9_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51437\,
            in1 => \N__48002\,
            in2 => \_gnd_net_\,
            in3 => \N__70117\,
            lcout => \ALU.a_15_m1_9\,
            ltout => \ALU.a_15_m1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_9_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__66844\,
            in1 => \N__58552\,
            in2 => \N__43556\,
            in3 => \N__52805\,
            lcout => \ALU.aZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73172\,
            ce => \N__71198\,
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIV0F38_0_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001110010"
        )
    port map (
            in0 => \N__49831\,
            in1 => \N__43532\,
            in2 => \N__43511\,
            in3 => \_gnd_net_\,
            lcout => bus_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI5FSP_4_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46897\,
            in1 => \N__44139\,
            in2 => \_gnd_net_\,
            in3 => \N__43444\,
            lcout => \ALU.b_RNI5FSPZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIHV2S_9_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__72348\,
            in1 => \N__46654\,
            in2 => \_gnd_net_\,
            in3 => \N__46898\,
            lcout => \ALU.c_RNIHV2SZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9R8E_4_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46896\,
            in1 => \N__43402\,
            in2 => \_gnd_net_\,
            in3 => \N__43349\,
            lcout => \ALU.d_RNI9R8EZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI83KC1_14_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__57582\,
            in1 => \N__67964\,
            in2 => \_gnd_net_\,
            in3 => \N__43303\,
            lcout => \ALU.b_RNI83KC1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_7_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101011000"
        )
    port map (
            in0 => \N__58886\,
            in1 => \N__51931\,
            in2 => \N__67242\,
            in3 => \N__51853\,
            lcout => h_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73183\,
            ce => \N__69449\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIO7K62_7_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__46402\,
            in1 => \N__43937\,
            in2 => \N__48867\,
            in3 => \N__46780\,
            lcout => \ALU.N_1204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISJ0R1_7_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__46781\,
            in1 => \N__51806\,
            in2 => \N__43822\,
            in3 => \N__43616\,
            lcout => OPEN,
            ltout => \ALU.N_1252_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO5IF4_7_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53889\,
            in2 => \N__43649\,
            in3 => \N__43646\,
            lcout => OPEN,
            ltout => \ALU.d_RNIO5IF4Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIM3JB6_7_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__71436\,
            in2 => \N__43640\,
            in3 => \N__43637\,
            lcout => OPEN,
            ltout => \ALU.d_RNIM3JB6Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3GMNC_7_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__53305\,
            in1 => \N__49580\,
            in2 => \N__43622\,
            in3 => \N__43759\,
            lcout => \ALU.status_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIB0OT_7_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__46610\,
            in1 => \N__43915\,
            in2 => \N__46298\,
            in3 => \N__47273\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIN3QQ1_7_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__46403\,
            in1 => \N__48871\,
            in2 => \N__43619\,
            in3 => \N__47190\,
            lcout => \ALU.N_1092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNID4971_7_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__53401\,
            in1 => \N__48346\,
            in2 => \N__49081\,
            in3 => \N__43979\,
            lcout => \ALU.operand2_6_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_RNIBU251_7_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__43980\,
            in1 => \N__46294\,
            in2 => \N__46609\,
            in3 => \N__53400\,
            lcout => \ALU.operand2_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNID6UV_7_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__48347\,
            in1 => \N__43914\,
            in2 => \N__49080\,
            in3 => \N__47272\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRF6F1_7_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__43815\,
            in1 => \N__51805\,
            in2 => \N__43799\,
            in3 => \N__47191\,
            lcout => OPEN,
            ltout => \ALU.N_1140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNILNEJ3_7_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54118\,
            in2 => \N__43796\,
            in3 => \N__43793\,
            lcout => \aluOut_7\,
            ltout => \aluOut_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIG8VE5_1_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__50305\,
            in1 => \N__43787\,
            in2 => \N__43772\,
            in3 => \N__50213\,
            lcout => \N_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m267_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__78769\,
            in1 => \N__78026\,
            in2 => \N__75993\,
            in3 => \N__77295\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m442_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__44307\,
            in1 => \N__79788\,
            in2 => \N__43748\,
            in3 => \N__76585\,
            lcout => \PROM.ROMDATA.m442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m282_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__78766\,
            in1 => \N__78023\,
            in2 => \N__75990\,
            in3 => \N__77292\,
            lcout => \PROM.ROMDATA.m282\,
            ltout => \PROM.ROMDATA.m282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.dout_13_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__44308\,
            in1 => \N__43703\,
            in2 => \N__43679\,
            in3 => \N__76586\,
            lcout => \CONTROL.ctrlOut_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.dout_13C_net\,
            ce => \N__44397\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m444_bm_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000111"
        )
    port map (
            in0 => \N__78767\,
            in1 => \N__78024\,
            in2 => \N__75991\,
            in3 => \N__77293\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m444_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m447_ns_1_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__44336\,
            in1 => \N__79787\,
            in2 => \N__44327\,
            in3 => \N__76584\,
            lcout => \PROM.ROMDATA.m447_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m289_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001000"
        )
    port map (
            in0 => \N__78768\,
            in1 => \N__78025\,
            in2 => \N__75992\,
            in3 => \N__77294\,
            lcout => \PROM.ROMDATA.m289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m418_ns_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__64169\,
            in1 => \N__72684\,
            in2 => \N__44294\,
            in3 => \N__79300\,
            lcout => \PROM_ROMDATA_dintern_19ro\,
            ltout => \PROM_ROMDATA_dintern_19ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_19dflt_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44258\,
            in3 => \N__72256\,
            lcout => \controlWord_19\,
            ltout => \controlWord_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_3_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__70549\,
            in1 => \N__44243\,
            in2 => \N__44195\,
            in3 => \N__70790\,
            lcout => \A3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_3C_net\,
            ce => \N__70330\,
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_4_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__44192\,
            in1 => \N__70789\,
            in2 => \N__44162\,
            in3 => \N__70551\,
            lcout => \A4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_3C_net\,
            ce => \N__70330\,
            sr => \_gnd_net_\
        );

    \RAM.un1_WR_105_0_7_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44101\,
            in1 => \N__44059\,
            in2 => \N__44962\,
            in3 => \N__44032\,
            lcout => \RAM.un1_WR_105_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_15_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__45020\,
            in1 => \N__70788\,
            in2 => \N__53534\,
            in3 => \N__70550\,
            lcout => \A15_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_3C_net\,
            ce => \N__70330\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m266_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111011111111"
        )
    port map (
            in0 => \N__78731\,
            in1 => \N__77199\,
            in2 => \N__75614\,
            in3 => \N__77909\,
            lcout => \PROM.ROMDATA.m266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m446_bm_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__64007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__75304\,
            lcout => \PROM.ROMDATA.m446_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m157_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__78732\,
            in1 => \N__77200\,
            in2 => \_gnd_net_\,
            in3 => \N__77910\,
            lcout => \PROM.ROMDATA.m157\,
            ltout => \PROM.ROMDATA.m157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m268_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100010001"
        )
    port map (
            in0 => \N__44945\,
            in1 => \N__76603\,
            in2 => \N__44939\,
            in3 => \N__75299\,
            lcout => \PROM.ROMDATA.m268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m265_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__78733\,
            in1 => \N__77201\,
            in2 => \N__75615\,
            in3 => \N__77911\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m270_bm_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__79714\,
            in1 => \_gnd_net_\,
            in2 => \N__44936\,
            in3 => \N__44933\,
            lcout => \PROM.ROMDATA.m270_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.aluOperation_6_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__44909\,
            in1 => \N__44900\,
            in2 => \N__44774\,
            in3 => \N__44704\,
            lcout => \aluOperation_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.aluOperation_6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m278_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__64235\,
            in1 => \N__76604\,
            in2 => \N__79830\,
            in3 => \N__75303\,
            lcout => \PROM.ROMDATA.N_544_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_RNIUD971_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45144\,
            in1 => \N__45641\,
            in2 => \_gnd_net_\,
            in3 => \N__45296\,
            lcout => \progRomAddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m258_bm_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__75306\,
            in1 => \N__64105\,
            in2 => \N__76579\,
            in3 => \N__47708\,
            lcout => \PROM.ROMDATA.m258_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_1_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_RNIQ9971_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45161\,
            in1 => \N__45155\,
            in2 => \_gnd_net_\,
            in3 => \N__45143\,
            lcout => \progRomAddress_5\,
            ltout => \progRomAddress_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m243_1_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__79248\,
            in1 => \N__76463\,
            in2 => \N__45098\,
            in3 => \N__75305\,
            lcout => \PROM.ROMDATA.m243_1\,
            ltout => \PROM.ROMDATA.m243_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m244_ns_1_1_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110111011"
        )
    port map (
            in0 => \N__72648\,
            in1 => \N__79751\,
            in2 => \N__45095\,
            in3 => \N__64106\,
            lcout => \PROM.ROMDATA.m244_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_0_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45080\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.dout_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m260_1_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001111110011"
        )
    port map (
            in0 => \N__45065\,
            in1 => \N__79249\,
            in2 => \N__72725\,
            in3 => \N__64107\,
            lcout => \PROM.ROMDATA.m260_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNILC5J_2_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55077\,
            in1 => \N__54803\,
            in2 => \_gnd_net_\,
            in3 => \N__47564\,
            lcout => \N_417\,
            ltout => \N_417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m27_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__64597\,
            in1 => \N__64694\,
            in2 => \N__45326\,
            in3 => \N__77175\,
            lcout => \PROM.ROMDATA.N_28_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_2_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNI6OHF_6_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__64596\,
            in1 => \_gnd_net_\,
            in2 => \N__47816\,
            in3 => \N__45614\,
            lcout => \CONTROL.programCounter_ret_1_RNI6OHFZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_3_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45290\,
            lcout => \CONTROL.dout_reto_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_4_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m215_ns_1_N_2L1_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101011111"
        )
    port map (
            in0 => \N__75307\,
            in1 => \N__78943\,
            in2 => \N__64871\,
            in3 => \N__78634\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m215_ns_1_N_2L1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m215_ns_1_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110010"
        )
    port map (
            in0 => \N__79207\,
            in1 => \N__47714\,
            in2 => \N__45242\,
            in3 => \N__76500\,
            lcout => \PROM.ROMDATA.m215_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_3_i_a7_1_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110111"
        )
    port map (
            in0 => \N__53718\,
            in1 => \N__53666\,
            in2 => \N__45523\,
            in3 => \N__45402\,
            lcout => \CONTROL.g0_3_i_a7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_2_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45206\,
            lcout => \CONTROL_addrstack_reto_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m36_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__47570\,
            in1 => \N__54935\,
            in2 => \_gnd_net_\,
            in3 => \N__79286\,
            lcout => \PROM.ROMDATA.m36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m235_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111001011000"
        )
    port map (
            in0 => \N__77185\,
            in1 => \N__78806\,
            in2 => \N__75914\,
            in3 => \N__77878\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.N_526_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m238_bm_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__76534\,
            in1 => \N__64108\,
            in2 => \N__45542\,
            in3 => \N__75736\,
            lcout => \PROM.ROMDATA.m238_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m30_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011111100"
        )
    port map (
            in0 => \N__77186\,
            in1 => \N__78807\,
            in2 => \N__75915\,
            in3 => \N__77879\,
            lcout => \PROM.ROMDATA.m30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g0_5_0_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110111"
        )
    port map (
            in0 => \N__53719\,
            in1 => \N__53667\,
            in2 => \N__45524\,
            in3 => \N__45403\,
            lcout => \CONTROL.g0_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m258_am_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47687\,
            in1 => \N__47693\,
            in2 => \_gnd_net_\,
            in3 => \N__76535\,
            lcout => \PROM.ROMDATA.m258_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNINE5J_3_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55078\,
            in1 => \N__51125\,
            in2 => \_gnd_net_\,
            in3 => \N__47639\,
            lcout => \N_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m69_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64340\,
            in2 => \_gnd_net_\,
            in3 => \N__74023\,
            lcout => \PROM_ROMDATA_dintern_31_0__N_555_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m53_am_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__45566\,
            in1 => \N__51368\,
            in2 => \_gnd_net_\,
            in3 => \N__76605\,
            lcout => \PROM.ROMDATA.m53_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_5_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45680\,
            lcout => \CONTROL.dout_reto_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_RNIV5IG_6_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45572\,
            in1 => \N__45613\,
            in2 => \_gnd_net_\,
            in3 => \N__64598\,
            lcout => \CONTROL.programCounter_ret_19_RNIV5IGZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_6_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45632\,
            lcout => \CONTROL.addrstack_reto_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m53_bm_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__47804\,
            in1 => \N__45599\,
            in2 => \_gnd_net_\,
            in3 => \N__76606\,
            lcout => \PROM.ROMDATA.m53_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_6_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45593\,
            lcout => \CONTROL.dout_reto_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m7_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001100001"
        )
    port map (
            in0 => \N__77875\,
            in1 => \N__78831\,
            in2 => \N__75916\,
            in3 => \N__77187\,
            lcout => \PROM.ROMDATA.m7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m392_bm_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000001001"
        )
    port map (
            in0 => \N__77188\,
            in1 => \N__78808\,
            in2 => \N__76002\,
            in3 => \N__77876\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m392_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m392_ns_LC_19_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47552\,
            in2 => \N__45560\,
            in3 => \N__76607\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m392_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m401_ns_1_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__79418\,
            in1 => \N__47855\,
            in2 => \N__45557\,
            in3 => \N__79808\,
            lcout => \PROM.ROMDATA.m401_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m396_bm_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000010"
        )
    port map (
            in0 => \N__77877\,
            in1 => \N__78832\,
            in2 => \N__75917\,
            in3 => \N__77189\,
            lcout => \PROM.ROMDATA.m396_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m396_am_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__78995\,
            in1 => \N__45809\,
            in2 => \_gnd_net_\,
            in3 => \N__75746\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m396_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m396_ns_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45785\,
            in2 => \N__45779\,
            in3 => \N__76608\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m396_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m401_ns_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__79419\,
            in1 => \N__47771\,
            in2 => \N__45776\,
            in3 => \N__45773\,
            lcout => \PROM.ROMDATA.m401_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBQSTO_11_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61470\,
            in2 => \_gnd_net_\,
            in3 => \N__66049\,
            lcout => \ALU.c_RNIBQSTOZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNID9MMO_4_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__59910\,
            in1 => \N__59638\,
            in2 => \_gnd_net_\,
            in3 => \N__66763\,
            lcout => \ALU.N_607\,
            ltout => \ALU.N_607_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4DGL42_4_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45728\,
            in2 => \N__45683\,
            in3 => \N__66050\,
            lcout => \ALU.N_637\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIG5G6F1_10_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__61471\,
            in1 => \N__61636\,
            in2 => \N__66083\,
            in3 => \N__68909\,
            lcout => \ALU.c_RNIG5G6F1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIT73F71_10_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__68910\,
            in1 => \N__61472\,
            in2 => \N__61675\,
            in3 => \N__68507\,
            lcout => \ALU.c_RNIT73F71Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFHB5A2_8_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100100110001"
        )
    port map (
            in0 => \N__66051\,
            in1 => \N__45962\,
            in2 => \N__62026\,
            in3 => \N__62883\,
            lcout => \ALU.N_643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4N3K21_8_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__62884\,
            in1 => \N__56416\,
            in2 => \N__68530\,
            in3 => \N__62010\,
            lcout => \ALU.d_RNI4N3K21Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIH8D821_8_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110010100000"
        )
    port map (
            in0 => \N__55949\,
            in1 => \N__62882\,
            in2 => \N__62025\,
            in3 => \N__56120\,
            lcout => \ALU.d_RNIH8D821Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_335_c_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46127\,
            in2 => \N__45929\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_10_0_\,
            carryout => \ALU.mult_11_c11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_335_c_RNI96NH82_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45917\,
            in2 => \N__45911\,
            in3 => \N__45893\,
            lcout => \ALU.mult_11_12\,
            ltout => OPEN,
            carryin => \ALU.mult_11_c11\,
            carryout => \ALU.mult_11_c12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_341_c_RNIVBI3U1_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45890\,
            in2 => \N__45878\,
            in3 => \N__45860\,
            lcout => \ALU.mult_11_13\,
            ltout => OPEN,
            carryin => \ALU.mult_11_c12\,
            carryout => \ALU.mult_11_c13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_347_c_RNITD0CL1_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45815\,
            in2 => \N__45857\,
            in3 => \N__45827\,
            lcout => \ALU.mult_11_14\,
            ltout => OPEN,
            carryin => \ALU.mult_11_c13\,
            carryout => \ALU.mult_11_c14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_11_c14_THRU_LUT4_0_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45824\,
            lcout => \ALU.mult_11_c14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIOSF6H_11_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__61473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__68395\,
            lcout => \ALU.c_RNIOSF6HZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_335_c_RNO_0_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61446\,
            in2 => \_gnd_net_\,
            in3 => \N__66702\,
            lcout => \ALU.mult_335_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPTT4O_8_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__66703\,
            in1 => \N__62017\,
            in2 => \_gnd_net_\,
            in3 => \N__62209\,
            lcout => \ALU.N_835\,
            ltout => \ALU.N_835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGSBJN2_8_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__66059\,
            in1 => \N__68929\,
            in2 => \N__46121\,
            in3 => \N__46075\,
            lcout => OPEN,
            ltout => \ALU.rshift_7_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIND5CS4_12_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__46118\,
            in1 => \N__53333\,
            in2 => \N__46100\,
            in3 => \N__68926\,
            lcout => OPEN,
            ltout => \ALU.N_925_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIEPHJC7_12_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52685\,
            in2 => \N__46097\,
            in3 => \N__45968\,
            lcout => \ALU.a_15_m0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIL9TBN2_6_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__65276\,
            in1 => \N__68924\,
            in2 => \N__46094\,
            in3 => \N__66058\,
            lcout => OPEN,
            ltout => \ALU.rshift_7_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI9GG8Q4_8_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__68925\,
            in1 => \N__46076\,
            in2 => \N__46055\,
            in3 => \N__52705\,
            lcout => \ALU.N_921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI08R632_15_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__70007\,
            in1 => \N__46032\,
            in2 => \_gnd_net_\,
            in3 => \N__45983\,
            lcout => \ALU.c_RNI08R632Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_1_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__59290\,
            in1 => \N__69748\,
            in2 => \N__52246\,
            in3 => \N__69012\,
            lcout => \ALU.eZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73156\,
            ce => \N__69243\,
            sr => \_gnd_net_\
        );

    \ALU.e_0_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69170\,
            in1 => \N__52123\,
            in2 => \N__69752\,
            in3 => \N__52033\,
            lcout => \ALU.eZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73156\,
            ce => \N__69243\,
            sr => \_gnd_net_\
        );

    \ALU.e_7_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101011000"
        )
    port map (
            in0 => \N__58877\,
            in1 => \N__51904\,
            in2 => \N__67266\,
            in3 => \N__51858\,
            lcout => \ALU.eZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73156\,
            ce => \N__69243\,
            sr => \_gnd_net_\
        );

    \ALU.e_8_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__51727\,
            in1 => \N__67226\,
            in2 => \N__51788\,
            in3 => \N__51638\,
            lcout => \ALU.eZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73156\,
            ce => \N__69243\,
            sr => \_gnd_net_\
        );

    \ALU.e_15_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__67225\,
            in1 => \N__52933\,
            in2 => \N__59176\,
            in3 => \N__53006\,
            lcout => \ALU.eZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73156\,
            ce => \N__69243\,
            sr => \_gnd_net_\
        );

    \ALU.e_9_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__52871\,
            in1 => \N__66843\,
            in2 => \N__58547\,
            in3 => \N__52787\,
            lcout => \ALU.eZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73156\,
            ce => \N__69243\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIIM1475_12_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__68812\,
            in1 => \N__46178\,
            in2 => \_gnd_net_\,
            in3 => \N__46159\,
            lcout => \ALU.N_707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_14_c_RNI134CV5_0_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__46523\,
            in1 => \N__63524\,
            in2 => \N__67255\,
            in3 => \N__68483\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_14_c_RNI134CV5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_14_c_RNIKS9S5H_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46139\,
            in2 => \N__46133\,
            in3 => \N__46514\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_14_c_RNIKS9S5HZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI3NTFTL_15_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000011111"
        )
    port map (
            in0 => \N__59338\,
            in1 => \N__67219\,
            in2 => \N__46130\,
            in3 => \N__46565\,
            lcout => \ALU.a_15_1_15\,
            ltout => \ALU.a_15_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100001101"
        )
    port map (
            in0 => \N__59169\,
            in1 => \N__67212\,
            in2 => \N__46553\,
            in3 => \N__52987\,
            lcout => \ALU.aZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73162\,
            ce => \N__71207\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4MD4S4_2_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46477\,
            in1 => \N__46500\,
            in2 => \_gnd_net_\,
            in3 => \N__68810\,
            lcout => \ALU.N_812\,
            ltout => \ALU.N_812_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_14_c_RNI134CV5_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110101"
        )
    port map (
            in0 => \N__68482\,
            in1 => \N__63523\,
            in2 => \N__46517\,
            in3 => \N__67208\,
            lcout => \ALU.addsub_cry_14_c_RNI134CVZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIDEP395_2_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__46501\,
            in1 => \N__68481\,
            in2 => \N__46481\,
            in3 => \N__68811\,
            lcout => \ALU.lshift_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_1_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__59248\,
            in1 => \N__52236\,
            in2 => \N__69678\,
            in3 => \N__69009\,
            lcout => \ALU.cZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73173\,
            ce => \N__71558\,
            sr => \_gnd_net_\
        );

    \ALU.c_0_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69149\,
            in1 => \N__52122\,
            in2 => \N__69747\,
            in3 => \N__52049\,
            lcout => \ALU.cZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73173\,
            ce => \N__71558\,
            sr => \_gnd_net_\
        );

    \ALU.c_7_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101100100"
        )
    port map (
            in0 => \N__58889\,
            in1 => \N__67273\,
            in2 => \N__51933\,
            in3 => \N__51851\,
            lcout => \ALU.cZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73173\,
            ce => \N__71558\,
            sr => \_gnd_net_\
        );

    \ALU.c_8_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67271\,
            in1 => \N__51776\,
            in2 => \N__51728\,
            in3 => \N__51633\,
            lcout => \ALU.cZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73173\,
            ce => \N__71558\,
            sr => \_gnd_net_\
        );

    \ALU.c_15_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101000101"
        )
    port map (
            in0 => \N__52931\,
            in1 => \N__67272\,
            in2 => \N__59177\,
            in3 => \N__53009\,
            lcout => \ALU.cZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73173\,
            ce => \N__71558\,
            sr => \_gnd_net_\
        );

    \ALU.c_9_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__58524\,
            in1 => \N__52879\,
            in2 => \N__52807\,
            in3 => \N__66833\,
            lcout => \ALU.cZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73173\,
            ce => \N__71558\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNI500DG_7_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__55886\,
            in1 => \N__63217\,
            in2 => \_gnd_net_\,
            in3 => \N__62158\,
            lcout => \ALU.d_RNI500DGZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI5KAEG_7_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011101000"
        )
    port map (
            in0 => \N__62157\,
            in1 => \N__74778\,
            in2 => \N__63273\,
            in3 => \N__55887\,
            lcout => \ALU.log_1_7\,
            ltout => \ALU.log_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_492_c_RNIQ5B457_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59100\,
            in2 => \N__46643\,
            in3 => \N__46640\,
            lcout => OPEN,
            ltout => \ALU.mult_492_c_RNIQ5BZ0Z457_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_492_c_RNIGN2JEC_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__59101\,
            in1 => \N__70096\,
            in2 => \N__46625\,
            in3 => \N__46622\,
            lcout => \ALU.mult_492_c_RNIGN2JECZ0\,
            ltout => \ALU.mult_492_c_RNIGN2JECZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_7_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011000110010"
        )
    port map (
            in0 => \N__67230\,
            in1 => \N__58887\,
            in2 => \N__46613\,
            in3 => \N__51932\,
            lcout => \ALU.aZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73184\,
            ce => \N__71176\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO75BG_7_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__62156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55885\,
            lcout => \ALU.d_RNIO75BGZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_d_d_s_0_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__70095\,
            in1 => \N__69790\,
            in2 => \_gnd_net_\,
            in3 => \N__63218\,
            lcout => \ALU.a_15_m2_d_d_sZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2s2_i_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69789\,
            in2 => \_gnd_net_\,
            in3 => \N__70094\,
            lcout => \ALU.a_15_sm0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI9SHF_14_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52291\,
            in1 => \N__67312\,
            in2 => \_gnd_net_\,
            in3 => \N__46923\,
            lcout => \ALU.c_RNI9SHFZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m2_s_1_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__69972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59262\,
            lcout => \ALU.a_15_m2_sZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPNGFE_14_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__53306\,
            in1 => \N__47062\,
            in2 => \N__46697\,
            in3 => \N__49581\,
            lcout => \ALU.status_19_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI5CPU_14_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52447\,
            in1 => \N__57454\,
            in2 => \_gnd_net_\,
            in3 => \N__46924\,
            lcout => OPEN,
            ltout => \ALU.a_RNI5CPUZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINT5A2_14_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__46850\,
            in1 => \N__53938\,
            in2 => \N__46844\,
            in3 => \N__46827\,
            lcout => OPEN,
            ltout => \ALU.operand2_7_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIFU325_14_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__53939\,
            in1 => \N__46733\,
            in2 => \N__46724\,
            in3 => \N__46721\,
            lcout => OPEN,
            ltout => \ALU.operand2_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNINISC7_14_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46712\,
            in2 => \N__46700\,
            in3 => \N__71454\,
            lcout => \ALU.d_RNINISC7Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_RNI80U51_14_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__57458\,
            in1 => \N__47275\,
            in2 => \N__52451\,
            in3 => \N__54298\,
            lcout => OPEN,
            ltout => \ALU.dout_3_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIG4FM1_14_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__67313\,
            in1 => \N__52284\,
            in2 => \N__46688\,
            in3 => \N__47192\,
            lcout => \ALU.N_1099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNIA8AE1_14_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__67963\,
            in1 => \N__47274\,
            in2 => \N__57586\,
            in3 => \N__54299\,
            lcout => OPEN,
            ltout => \ALU.dout_6_ns_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKK772_14_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__67784\,
            in1 => \N__57859\,
            in2 => \N__47216\,
            in3 => \N__47193\,
            lcout => OPEN,
            ltout => \ALU.N_1147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI7T474_14_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47099\,
            in2 => \N__47093\,
            in3 => \N__54139\,
            lcout => \aluOut_14\,
            ltout => \aluOut_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI51G56_1_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__47090\,
            in1 => \N__50325\,
            in2 => \N__47075\,
            in3 => \N__50214\,
            lcout => \N_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.increment_1_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__47051\,
            in1 => \N__47011\,
            in2 => \N__46964\,
            in3 => \N__54686\,
            lcout => \CONTROL.incrementZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.increment_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIH85J_0_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55079\,
            in1 => \N__50990\,
            in2 => \_gnd_net_\,
            in3 => \N__47615\,
            lcout => \N_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m399_bm_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000100"
        )
    port map (
            in0 => \N__78027\,
            in1 => \N__78823\,
            in2 => \N__75994\,
            in3 => \N__77296\,
            lcout => \PROM.ROMDATA.m399_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m422_am_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000100100"
        )
    port map (
            in0 => \N__77297\,
            in1 => \N__75938\,
            in2 => \N__78862\,
            in3 => \N__78028\,
            lcout => \PROM.ROMDATA.m422_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m422_bm_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__75939\,
            in1 => \N__64863\,
            in2 => \_gnd_net_\,
            in3 => \N__78827\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m422_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m422_ns_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47372\,
            in2 => \N__47366\,
            in3 => \N__76587\,
            lcout => \PROM.ROMDATA.m422_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m381_bm_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__75940\,
            in1 => \N__50447\,
            in2 => \N__76623\,
            in3 => \N__64254\,
            lcout => \PROM.ROMDATA.m381_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m482_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__78828\,
            in1 => \N__47514\,
            in2 => \N__64875\,
            in3 => \N__75941\,
            lcout => \PROM.ROMDATA.N_551_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m298_ns_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47345\,
            in1 => \N__64031\,
            in2 => \_gnd_net_\,
            in3 => \N__76483\,
            lcout => \PROM.ROMDATA.m298_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_RNIMGJ31_4_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__73721\,
            in1 => \_gnd_net_\,
            in2 => \N__47681\,
            in3 => \N__55168\,
            lcout => \CONTROL.programCounter_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m35_1_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__76482\,
            in1 => \N__47726\,
            in2 => \N__50645\,
            in3 => \N__79761\,
            lcout => \PROM.ROMDATA.m35_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m498_bm_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011010111"
        )
    port map (
            in0 => \N__78830\,
            in1 => \N__77932\,
            in2 => \N__77314\,
            in3 => \N__75934\,
            lcout => \PROM.ROMDATA.m498_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m124_e_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__73720\,
            in1 => \N__79762\,
            in2 => \N__47680\,
            in3 => \N__55167\,
            lcout => \PROM.ROMDATA.N_543_mux_2\,
            ltout => \PROM.ROMDATA.N_543_mux_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m176_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__64323\,
            in1 => \N__79293\,
            in2 => \N__47312\,
            in3 => \N__75932\,
            lcout => \PROM.ROMDATA.N_559_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m392_am_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__75933\,
            in1 => \N__78829\,
            in2 => \N__64324\,
            in3 => \N__78980\,
            lcout => \PROM.ROMDATA.m392_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m163_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__77198\,
            in1 => \_gnd_net_\,
            in2 => \N__77994\,
            in3 => \N__78730\,
            lcout => \PROM.ROMDATA.m163\,
            ltout => \PROM.ROMDATA.m163_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m176_x_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__75247\,
            in1 => \_gnd_net_\,
            in2 => \N__47540\,
            in3 => \N__79208\,
            lcout => \PROM.ROMDATA.m176_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m474_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__79209\,
            in1 => \N__75248\,
            in2 => \N__47523\,
            in3 => \N__64965\,
            lcout => \PROM.ROMDATA.N_569_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m109_am_1_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000101000110"
        )
    port map (
            in0 => \N__78727\,
            in1 => \N__77842\,
            in2 => \N__75539\,
            in3 => \N__77196\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m109_am_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m109_am_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101101111"
        )
    port map (
            in0 => \N__76479\,
            in1 => \N__75243\,
            in2 => \N__47429\,
            in3 => \N__78729\,
            lcout => \PROM.ROMDATA.m109_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m11_am_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110110011110"
        )
    port map (
            in0 => \N__78728\,
            in1 => \N__77843\,
            in2 => \N__75540\,
            in3 => \N__77197\,
            lcout => \PROM.ROMDATA.m11_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_0_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47426\,
            lcout => \CONTROL_addrstack_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73225\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_0_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__47403\,
            in1 => \N__73712\,
            in2 => \_gnd_net_\,
            in3 => \N__50955\,
            lcout => \CONTROL.programCounter_1_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73225\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIPG5J_4_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55057\,
            in1 => \N__55183\,
            in2 => \_gnd_net_\,
            in3 => \N__55301\,
            lcout => \N_419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_1_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47660\,
            lcout => \CONTROL_addrstack_reto_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_RNIEO8J_3_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55120\,
            in1 => \N__47635\,
            in2 => \_gnd_net_\,
            in3 => \N__64465\,
            lcout => \CONTROL.programCounter_ret_19_RNIEO8JZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNILA8I_3_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__64466\,
            in1 => \N__51121\,
            in2 => \_gnd_net_\,
            in3 => \N__55119\,
            lcout => OPEN,
            ltout => \CONTROL.programCounter_ret_1_RNILA8IZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_fast_RNI93CH1_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55056\,
            in1 => \_gnd_net_\,
            in2 => \N__47624\,
            in3 => \N__47621\,
            lcout => \progRomAddress_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIF48I_0_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47611\,
            in1 => \N__55118\,
            in2 => \_gnd_net_\,
            in3 => \N__50947\,
            lcout => \CONTROL.programCounter_ret_1_RNIF48IZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_3_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47600\,
            lcout => \CONTROL_addrstack_reto_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m35_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__47588\,
            in1 => \N__47582\,
            in2 => \N__54923\,
            in3 => \N__79715\,
            lcout => \PROM.ROMDATA.m35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIJ88I_2_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47563\,
            in1 => \N__64692\,
            in2 => \_gnd_net_\,
            in3 => \N__55123\,
            lcout => \CONTROL.programCounter_ret_1_RNIJ88IZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_1_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__75291\,
            in1 => \N__78625\,
            in2 => \_gnd_net_\,
            in3 => \N__77613\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m215_ns_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m215_ns_1_1_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101111001"
        )
    port map (
            in0 => \N__77114\,
            in1 => \N__76499\,
            in2 => \N__47717\,
            in3 => \N__75292\,
            lcout => \PROM.ROMDATA.m215_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m178_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__78636\,
            in1 => \N__77615\,
            in2 => \_gnd_net_\,
            in3 => \N__77116\,
            lcout => \PROM.ROMDATA.m178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_RNICM8J_2_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__54802\,
            in1 => \N__64693\,
            in2 => \_gnd_net_\,
            in3 => \N__55124\,
            lcout => \CONTROL.programCounter_ret_19_RNICM8JZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m256_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000110010"
        )
    port map (
            in0 => \N__78635\,
            in1 => \N__77614\,
            in2 => \N__75613\,
            in3 => \N__77115\,
            lcout => \PROM.ROMDATA.m256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_35_fast_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50834\,
            in2 => \_gnd_net_\,
            in3 => \N__50898\,
            lcout => \CONTROL.programCounter11_reto_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m38_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101101010"
        )
    port map (
            in0 => \N__77620\,
            in1 => \N__78688\,
            in2 => \N__75919\,
            in3 => \N__76937\,
            lcout => \PROM.ROMDATA.m38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m251_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100111000"
        )
    port map (
            in0 => \N__76933\,
            in1 => \N__78692\,
            in2 => \N__75912\,
            in3 => \N__77618\,
            lcout => \PROM.ROMDATA.m251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m253_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000101010"
        )
    port map (
            in0 => \N__77617\,
            in1 => \N__75726\,
            in2 => \N__78833\,
            in3 => \N__76934\,
            lcout => \PROM.ROMDATA.m253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m389_bm_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000010"
        )
    port map (
            in0 => \N__76936\,
            in1 => \N__78693\,
            in2 => \N__75913\,
            in3 => \N__77619\,
            lcout => \PROM.ROMDATA.m389_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m20_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__64741\,
            in1 => \N__64698\,
            in2 => \N__64641\,
            in3 => \N__76932\,
            lcout => \PROM.ROMDATA.m20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_6_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47846\,
            lcout => \CONTROL.programCounter_1_reto_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m51_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110110001"
        )
    port map (
            in0 => \N__77616\,
            in1 => \N__78687\,
            in2 => \N__75918\,
            in3 => \N__76935\,
            lcout => \PROM.ROMDATA.m51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m433_am_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__76528\,
            in1 => \N__74447\,
            in2 => \N__73373\,
            in3 => \N__75750\,
            lcout => \PROM.ROMDATA.m433_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m399_am_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010001"
        )
    port map (
            in0 => \N__77874\,
            in1 => \N__75383\,
            in2 => \N__64861\,
            in3 => \N__78639\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m399_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m399_ns_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76529\,
            in2 => \N__47786\,
            in3 => \N__47783\,
            lcout => \PROM.ROMDATA.m399_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m461_ns_1_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000111"
        )
    port map (
            in0 => \N__64199\,
            in1 => \N__79391\,
            in2 => \N__47906\,
            in3 => \N__79850\,
            lcout => \PROM.ROMDATA.m461_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_36_4_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47744\,
            lcout => \CONTROL_addrstack_reto_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m22_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000010011"
        )
    port map (
            in0 => \N__78638\,
            in1 => \N__77873\,
            in2 => \N__75676\,
            in3 => \N__77184\,
            lcout => \PROM.ROMDATA.m22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m451_bm_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__64837\,
            in1 => \N__75384\,
            in2 => \N__73892\,
            in3 => \N__78640\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m451_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m451_ns_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76530\,
            in2 => \N__47918\,
            in3 => \N__47915\,
            lcout => \PROM.ROMDATA.m451_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m375_bm_LC_20_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__47873\,
            in1 => \N__76527\,
            in2 => \N__74285\,
            in3 => \N__75790\,
            lcout => \PROM.ROMDATA.m375_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m280_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__78994\,
            in1 => \N__75791\,
            in2 => \N__76602\,
            in3 => \N__78695\,
            lcout => \PROM.ROMDATA.m280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m376_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001010010000"
        )
    port map (
            in0 => \N__77882\,
            in1 => \N__75789\,
            in2 => \N__78835\,
            in3 => \N__77192\,
            lcout => \PROM.ROMDATA.m376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m255_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__77881\,
            in1 => \_gnd_net_\,
            in2 => \N__78834\,
            in3 => \N__77190\,
            lcout => \PROM.ROMDATA.N_256_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m389_am_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__78993\,
            in1 => \N__78696\,
            in2 => \N__75950\,
            in3 => \N__77880\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m389_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m389_ns_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47867\,
            in2 => \N__47858\,
            in3 => \N__76526\,
            lcout => \PROM.ROMDATA.m389_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m103_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__77191\,
            in1 => \N__78700\,
            in2 => \_gnd_net_\,
            in3 => \N__77883\,
            lcout => \PROM.ROMDATA.m103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIMNQ8E1_0_12_LC_21_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__61010\,
            in1 => \N__66063\,
            in2 => \N__61225\,
            in3 => \N__66757\,
            lcout => OPEN,
            ltout => \ALU.lshift_3_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIUU8GB2_10_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__66064\,
            in1 => \N__61640\,
            in2 => \N__48092\,
            in3 => \N__61474\,
            lcout => OPEN,
            ltout => \ALU.N_645_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI5G4OF5_10_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__68918\,
            in1 => \N__68511\,
            in2 => \N__48089\,
            in3 => \N__48032\,
            lcout => OPEN,
            ltout => \ALU.a_15_m1_am_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIRFBHE9_0_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__48016\,
            in1 => \N__48086\,
            in2 => \N__48065\,
            in3 => \N__68510\,
            lcout => \ALU.d_RNIRFBHE9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBK47O_0_8_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__62023\,
            in1 => \N__62885\,
            in2 => \_gnd_net_\,
            in3 => \N__66756\,
            lcout => OPEN,
            ltout => \ALU.N_611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMQD952_8_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__66062\,
            in1 => \_gnd_net_\,
            in2 => \N__48062\,
            in3 => \N__48058\,
            lcout => \ALU.N_641\,
            ltout => \ALU.N_641_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNITG2137_0_LC_21_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__68509\,
            in1 => \N__47942\,
            in2 => \N__48026\,
            in3 => \N__48015\,
            lcout => \ALU.d_RNITG2137Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIQGO2C2_0_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110011"
        )
    port map (
            in0 => \N__66061\,
            in1 => \N__68508\,
            in2 => \N__47990\,
            in3 => \N__68917\,
            lcout => \ALU.a_15_m1_am_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0OR9G_3_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100010111"
        )
    port map (
            in0 => \N__63253\,
            in1 => \N__60260\,
            in2 => \N__74816\,
            in3 => \N__68490\,
            lcout => \ALU.a_15_m3_d_d_0_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBRG4Q9_0_12_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__58497\,
            in1 => \N__70171\,
            in2 => \N__48188\,
            in3 => \N__48175\,
            lcout => \ALU.c_RNIBRG4Q9_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_555_c_RNIJF56AM_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__69640\,
            in1 => \N__48290\,
            in2 => \_gnd_net_\,
            in3 => \N__48506\,
            lcout => \ALU.mult_555_c_RNIJF56AMZ0\,
            ltout => \ALU.mult_555_c_RNIJF56AMZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_12_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67742\,
            in2 => \N__48272\,
            in3 => \N__67654\,
            lcout => \ALU.aZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73157\,
            ce => \N__71197\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNI5SENO2_12_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__48236\,
            in1 => \N__68927\,
            in2 => \N__48212\,
            in3 => \N__66060\,
            lcout => OPEN,
            ltout => \ALU.lshift_7_ns_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI3I5IR4_8_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__68928\,
            in1 => \N__48677\,
            in2 => \N__48194\,
            in3 => \N__48710\,
            lcout => OPEN,
            ltout => \ALU.N_704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGNBT49_8_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__70169\,
            in1 => \N__48535\,
            in2 => \N__48191\,
            in3 => \N__68484\,
            lcout => \ALU.d_RNIGNBT49Z0Z_8\,
            ltout => \ALU.d_RNIGNBT49Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIBRG4Q9_12_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__58496\,
            in1 => \N__70170\,
            in2 => \N__48179\,
            in3 => \N__48174\,
            lcout => \ALU.c_RNIBRG4Q9Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_8_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67231\,
            in1 => \N__51784\,
            in2 => \N__51723\,
            in3 => \N__51637\,
            lcout => h_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73163\,
            ce => \N__69452\,
            sr => \_gnd_net_\
        );

    \ALU.h_15_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__67207\,
            in1 => \N__52934\,
            in2 => \N__59140\,
            in3 => \N__53012\,
            lcout => h_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73163\,
            ce => \N__69452\,
            sr => \_gnd_net_\
        );

    \ALU.mult_555_c_RNI5VJUOI_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__61042\,
            in1 => \N__67205\,
            in2 => \_gnd_net_\,
            in3 => \N__48518\,
            lcout => \ALU.mult_555_c_RNI5VJUOIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_546_c_RNIJOT4J8_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__66896\,
            in1 => \N__67206\,
            in2 => \_gnd_net_\,
            in3 => \N__48500\,
            lcout => \ALU.mult_546_c_RNIJOT4JZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_3_0_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__61277\,
            in1 => \N__60839\,
            in2 => \N__53360\,
            in3 => \N__61043\,
            lcout => OPEN,
            ltout => \ALU.status_14_12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_1_0_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__69512\,
            in1 => \N__48487\,
            in2 => \N__48428\,
            in3 => \N__53342\,
            lcout => \ALU.status_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_1_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111000001111"
        )
    port map (
            in0 => \N__59306\,
            in1 => \N__69002\,
            in2 => \N__52245\,
            in3 => \N__69729\,
            lcout => \ALU.bZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73174\,
            ce => \N__67931\,
            sr => \_gnd_net_\
        );

    \ALU.b_0_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69169\,
            in1 => \N__52118\,
            in2 => \N__69744\,
            in3 => \N__52050\,
            lcout => \ALU.bZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73174\,
            ce => \N__67931\,
            sr => \_gnd_net_\
        );

    \ALU.b_7_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011001010100"
        )
    port map (
            in0 => \N__58888\,
            in1 => \N__67218\,
            in2 => \N__51863\,
            in3 => \N__51930\,
            lcout => \ALU.bZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73174\,
            ce => \N__67931\,
            sr => \_gnd_net_\
        );

    \ALU.b_8_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67217\,
            in1 => \N__51775\,
            in2 => \N__51720\,
            in3 => \N__51632\,
            lcout => \ALU.bZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73174\,
            ce => \N__67931\,
            sr => \_gnd_net_\
        );

    \ALU.b_15_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110100011"
        )
    port map (
            in0 => \N__53007\,
            in1 => \N__52932\,
            in2 => \N__59141\,
            in3 => \N__67216\,
            lcout => \ALU.bZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73174\,
            ce => \N__67931\,
            sr => \_gnd_net_\
        );

    \ALU.b_9_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__52878\,
            in1 => \N__66827\,
            in2 => \N__58565\,
            in3 => \N__52786\,
            lcout => \ALU.bZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73174\,
            ce => \N__67931\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIS1QRR6_0_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__68480\,
            in1 => \N__48626\,
            in2 => \N__48719\,
            in3 => \N__48611\,
            lcout => \ALU.lshift_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_495_c_RNIKOB51J_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101100"
        )
    port map (
            in0 => \N__57065\,
            in1 => \N__57134\,
            in2 => \N__48806\,
            in3 => \N__48779\,
            lcout => \ALU.mult_495_c_RNIKOB51JZ0\,
            ltout => \ALU.mult_495_c_RNIKOB51JZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_8_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__67214\,
            in1 => \N__51704\,
            in2 => \N__48755\,
            in3 => \N__51779\,
            lcout => \ALU.aZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73185\,
            ce => \N__71163\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNINF0N42_0_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110011"
        )
    port map (
            in0 => \N__66066\,
            in1 => \N__68479\,
            in2 => \N__48596\,
            in3 => \N__68895\,
            lcout => \ALU.lshift_15_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIIDDI52_8_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48709\,
            in1 => \N__48673\,
            in2 => \_gnd_net_\,
            in3 => \N__66067\,
            lcout => \ALU.N_640\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_7_c_RNIDLTN71_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__61760\,
            in1 => \N__67213\,
            in2 => \_gnd_net_\,
            in3 => \N__51238\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_7_c_RNIDLTNZ0Z71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_7_c_RNIHPLU38_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__70159\,
            in1 => \N__67215\,
            in2 => \N__48620\,
            in3 => \N__48617\,
            lcout => \ALU.addsub_cry_7_c_RNIHPLUZ0Z38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIO3LAS3_0_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__66065\,
            in1 => \N__48610\,
            in2 => \N__48595\,
            in3 => \N__68894\,
            lcout => \ALU.N_809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_1_LC_21_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__59249\,
            in1 => \N__52241\,
            in2 => \N__69698\,
            in3 => \N__69010\,
            lcout => f_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73192\,
            ce => \N__67860\,
            sr => \_gnd_net_\
        );

    \ALU.f_0_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69117\,
            in1 => \N__52096\,
            in2 => \N__69699\,
            in3 => \N__52051\,
            lcout => f_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73192\,
            ce => \N__67860\,
            sr => \_gnd_net_\
        );

    \ALU.f_7_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101011000"
        )
    port map (
            in0 => \N__58884\,
            in1 => \N__51929\,
            in2 => \N__67286\,
            in3 => \N__51857\,
            lcout => f_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73192\,
            ce => \N__67860\,
            sr => \_gnd_net_\
        );

    \ALU.f_8_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67269\,
            in1 => \N__51777\,
            in2 => \N__51721\,
            in3 => \N__51634\,
            lcout => f_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73192\,
            ce => \N__67860\,
            sr => \_gnd_net_\
        );

    \ALU.f_15_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__67282\,
            in1 => \N__52936\,
            in2 => \N__59143\,
            in3 => \N__53010\,
            lcout => f_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73192\,
            ce => \N__67860\,
            sr => \_gnd_net_\
        );

    \ALU.f_9_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__52856\,
            in1 => \N__66831\,
            in2 => \N__58563\,
            in3 => \N__52801\,
            lcout => f_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73192\,
            ce => \N__67860\,
            sr => \_gnd_net_\
        );

    \ALU.g_1_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101000101"
        )
    port map (
            in0 => \N__52240\,
            in1 => \N__59291\,
            in2 => \N__69746\,
            in3 => \N__69011\,
            lcout => g_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73199\,
            ce => \N__70986\,
            sr => \_gnd_net_\
        );

    \ALU.g_0_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__52117\,
            in1 => \N__69106\,
            in2 => \N__69745\,
            in3 => \N__52052\,
            lcout => g_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73199\,
            ce => \N__70986\,
            sr => \_gnd_net_\
        );

    \ALU.g_7_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101011000"
        )
    port map (
            in0 => \N__58885\,
            in1 => \N__51937\,
            in2 => \N__67267\,
            in3 => \N__51852\,
            lcout => g_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73199\,
            ce => \N__70986\,
            sr => \_gnd_net_\
        );

    \ALU.g_8_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__51703\,
            in1 => \N__51783\,
            in2 => \N__67268\,
            in3 => \N__51636\,
            lcout => g_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73199\,
            ce => \N__70986\,
            sr => \_gnd_net_\
        );

    \ALU.g_15_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001100100011"
        )
    port map (
            in0 => \N__67232\,
            in1 => \N__52937\,
            in2 => \N__59120\,
            in3 => \N__53011\,
            lcout => g_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73199\,
            ce => \N__70986\,
            sr => \_gnd_net_\
        );

    \ALU.g_9_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__52866\,
            in1 => \N__66832\,
            in2 => \N__58551\,
            in3 => \N__52806\,
            lcout => g_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73199\,
            ce => \N__70986\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNID85GQ_0_15_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__59267\,
            in1 => \N__49194\,
            in2 => \N__50543\,
            in3 => \N__50513\,
            lcout => OPEN,
            ltout => \ALU.c_RNID85GQ_0Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI9DCRE2_15_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74524\,
            in2 => \N__50354\,
            in3 => \N__50504\,
            lcout => \ALU.c_RNI9DCRE2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNI117N5_1_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__63592\,
            in1 => \N__50326\,
            in2 => \N__50243\,
            in3 => \N__50215\,
            lcout => \N_208\,
            ltout => \N_208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIH202E_15_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__53757\,
            in1 => \N__53299\,
            in2 => \N__49844\,
            in3 => \N__49592\,
            lcout => \ALU.status_19_14\,
            ltout => \ALU.status_19_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJI6SH_15_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100000"
        )
    port map (
            in0 => \N__63594\,
            in1 => \_gnd_net_\,
            in2 => \N__49841\,
            in3 => \N__74833\,
            lcout => \ALU.c_RNIJI6SHZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.busState_1_RNIRLED8_0_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110001011"
        )
    port map (
            in0 => \N__49838\,
            in1 => \N__49832\,
            in2 => \N__49628\,
            in3 => \N__49593\,
            lcout => bus_15,
            ltout => \bus_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNID85GQ_15_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__50537\,
            in1 => \N__59266\,
            in2 => \N__50516\,
            in3 => \N__50512\,
            lcout => \ALU.c_RNID85GQZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIU5NNB_15_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__53758\,
            in1 => \N__63593\,
            in2 => \_gnd_net_\,
            in3 => \N__53300\,
            lcout => \ALU.un14_log_0_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m248_ns_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001111"
        )
    port map (
            in0 => \N__55221\,
            in1 => \N__76648\,
            in2 => \N__50921\,
            in3 => \N__76471\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m248_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m249_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__76472\,
            in1 => \N__79873\,
            in2 => \N__50498\,
            in3 => \N__50591\,
            lcout => \PROM.ROMDATA.m249\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m410_am_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__77956\,
            in1 => \N__78818\,
            in2 => \N__75814\,
            in3 => \N__77273\,
            lcout => \PROM.ROMDATA.m410_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m359_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__77272\,
            in1 => \_gnd_net_\,
            in2 => \N__78860\,
            in3 => \N__77955\,
            lcout => \PROM.ROMDATA.m359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m304_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000001000"
        )
    port map (
            in0 => \N__77274\,
            in1 => \N__75534\,
            in2 => \N__78861\,
            in3 => \N__77957\,
            lcout => \PROM.ROMDATA.m304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m71_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__77954\,
            in1 => \N__78814\,
            in2 => \_gnd_net_\,
            in3 => \N__77271\,
            lcout => \PROM.ROMDATA.N_72_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m413_bm_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__78819\,
            in1 => \N__75533\,
            in2 => \_gnd_net_\,
            in3 => \N__78984\,
            lcout => \PROM.ROMDATA.m413_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m150_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011111010"
        )
    port map (
            in0 => \N__77142\,
            in1 => \_gnd_net_\,
            in2 => \N__78038\,
            in3 => \N__78810\,
            lcout => \PROM.ROMDATA.m150\,
            ltout => \PROM.ROMDATA.m150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m195_am_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000101"
        )
    port map (
            in0 => \N__75529\,
            in1 => \N__50693\,
            in2 => \N__50651\,
            in3 => \N__76480\,
            lcout => \PROM.ROMDATA.m195_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m228_am_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001100001000"
        )
    port map (
            in0 => \N__77143\,
            in1 => \N__75528\,
            in2 => \N__78040\,
            in3 => \N__78812\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m228_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m229_1_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__50590\,
            in1 => \_gnd_net_\,
            in2 => \N__50648\,
            in3 => \N__76481\,
            lcout => \PROM.ROMDATA.m229_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m25_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001001"
        )
    port map (
            in0 => \N__77140\,
            in1 => \N__75526\,
            in2 => \N__78037\,
            in3 => \N__78809\,
            lcout => \PROM.ROMDATA.m25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m438_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__54863\,
            in1 => \N__50633\,
            in2 => \_gnd_net_\,
            in3 => \N__79843\,
            lcout => \PROM.ROMDATA.m438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m173_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__77141\,
            in1 => \N__75527\,
            in2 => \N__78039\,
            in3 => \N__78811\,
            lcout => \PROM.ROMDATA.m173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m246_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011011101"
        )
    port map (
            in0 => \N__78813\,
            in1 => \N__77953\,
            in2 => \_gnd_net_\,
            in3 => \N__77144\,
            lcout => \PROM.ROMDATA.m246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__g1_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__75659\,
            in1 => \N__73503\,
            in2 => \_gnd_net_\,
            in3 => \N__50579\,
            lcout => \PROM_ROMDATA_dintern_31_0__g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m145_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010001001"
        )
    port map (
            in0 => \N__77805\,
            in1 => \N__75653\,
            in2 => \N__78543\,
            in3 => \N__77123\,
            lcout => \PROM.ROMDATA.m145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m169_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__77125\,
            in1 => \N__78320\,
            in2 => \N__75890\,
            in3 => \N__77808\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m169_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m270_am_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__76485\,
            in1 => \N__79862\,
            in2 => \N__50723\,
            in3 => \N__50678\,
            lcout => \PROM.ROMDATA.m270_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m13_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__77124\,
            in1 => \N__78319\,
            in2 => \_gnd_net_\,
            in3 => \N__77806\,
            lcout => \PROM.ROMDATA.m13\,
            ltout => \PROM.ROMDATA.m13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m18_am_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__77807\,
            in1 => \N__75654\,
            in2 => \N__50696\,
            in3 => \N__78362\,
            lcout => \PROM.ROMDATA.m18_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m188_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101001010"
        )
    port map (
            in0 => \N__77122\,
            in1 => \N__78315\,
            in2 => \N__75889\,
            in3 => \N__77804\,
            lcout => \PROM.ROMDATA.m188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m263_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001001000000"
        )
    port map (
            in0 => \N__76484\,
            in1 => \N__75655\,
            in2 => \N__50687\,
            in3 => \N__64964\,
            lcout => \PROM.ROMDATA.m263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_RNIAK8J_1_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__54901\,
            in1 => \N__73766\,
            in2 => \_gnd_net_\,
            in3 => \N__55122\,
            lcout => \CONTROL.programCounter_ret_19_RNIAK8JZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_1_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50672\,
            lcout => \CONTROL.dout_reto_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_RNI8I8J_0_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__50986\,
            in1 => \N__55121\,
            in2 => \_gnd_net_\,
            in3 => \N__50948\,
            lcout => \CONTROL.programCounter_ret_19_RNI8I8JZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m74_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001111001"
        )
    port map (
            in0 => \N__77611\,
            in1 => \N__76966\,
            in2 => \N__75611\,
            in3 => \N__78468\,
            lcout => \PROM.ROMDATA.m74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m248_ns_1_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100111101"
        )
    port map (
            in0 => \N__78472\,
            in1 => \N__75287\,
            in2 => \N__76454\,
            in3 => \N__77612\,
            lcout => \PROM.ROMDATA.m248_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_fast_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__50899\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50835\,
            lcout => \CONTROL.un1_programCounter9_reto_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m104_ns_1_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000011000"
        )
    port map (
            in0 => \N__76965\,
            in1 => \N__75283\,
            in2 => \N__78704\,
            in3 => \_gnd_net_\,
            lcout => \PROM.ROMDATA.m104_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m284_1_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__78569\,
            in1 => \N__79747\,
            in2 => \N__75612\,
            in3 => \N__76268\,
            lcout => \PROM.ROMDATA.m284_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_fast_RNITMBH1_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55053\,
            in1 => \N__50747\,
            in2 => \_gnd_net_\,
            in3 => \N__50741\,
            lcout => \progRomAddress_0\,
            ltout => \progRomAddress_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m143_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001111010010"
        )
    port map (
            in0 => \N__77688\,
            in1 => \N__75236\,
            in2 => \N__50735\,
            in3 => \N__78327\,
            lcout => \PROM.ROMDATA.m143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m72_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111011111001"
        )
    port map (
            in0 => \N__78328\,
            in1 => \N__77689\,
            in2 => \N__75538\,
            in3 => \N__76927\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m80_am_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76273\,
            in2 => \N__50732\,
            in3 => \N__50729\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m80_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m93_ns_1_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__79314\,
            in1 => \N__79839\,
            in2 => \N__51050\,
            in3 => \N__64757\,
            lcout => \PROM.ROMDATA.m93_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m179_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000111001"
        )
    port map (
            in0 => \N__76925\,
            in1 => \N__75234\,
            in2 => \N__77893\,
            in3 => \N__78325\,
            lcout => \PROM.ROMDATA.m179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_fast_RNI5VBH1_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55054\,
            in1 => \N__51035\,
            in2 => \_gnd_net_\,
            in3 => \N__51029\,
            lcout => \progRomAddress_2\,
            ltout => \progRomAddress_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m127_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011011"
        )
    port map (
            in0 => \N__76926\,
            in1 => \N__75235\,
            in2 => \N__51023\,
            in3 => \N__78326\,
            lcout => \PROM.ROMDATA.m127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m196_ns_1_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__79844\,
            in1 => \N__55253\,
            in2 => \N__79413\,
            in3 => \N__50996\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m196_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m196_ns_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__51164\,
            in1 => \N__51020\,
            in2 => \N__51008\,
            in3 => \N__79318\,
            lcout => \PROM.ROMDATA.m196_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m185_am_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__51005\,
            in1 => \N__76269\,
            in2 => \_gnd_net_\,
            in3 => \N__74185\,
            lcout => \PROM.ROMDATA.m185_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m193_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000001"
        )
    port map (
            in0 => \N__77608\,
            in1 => \N__76977\,
            in2 => \N__75886\,
            in3 => \N__78677\,
            lcout => \PROM.ROMDATA.m193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m191_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111011111010"
        )
    port map (
            in0 => \N__76978\,
            in1 => \N__78679\,
            in2 => \N__75960\,
            in3 => \N__77609\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m195_bm_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__76270\,
            in1 => \_gnd_net_\,
            in2 => \N__51173\,
            in3 => \N__51170\,
            lcout => \PROM.ROMDATA.m195_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_3_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51158\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.programCounter_1_reto_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73267\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m92_am_LC_21_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000110100001"
        )
    port map (
            in0 => \N__77610\,
            in1 => \N__75821\,
            in2 => \N__55205\,
            in3 => \N__78678\,
            lcout => \PROM.ROMDATA.m92_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m62_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001011011100"
        )
    port map (
            in0 => \N__77794\,
            in1 => \N__78694\,
            in2 => \N__75903\,
            in3 => \N__77151\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m64_bm_LC_21_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__54922\,
            in1 => \_gnd_net_\,
            in2 => \N__51098\,
            in3 => \N__76322\,
            lcout => \PROM.ROMDATA.m64_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m65_ns_1_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__79319\,
            in1 => \N__51095\,
            in2 => \N__51086\,
            in3 => \N__79840\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m65_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m65_ns_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__51074\,
            in1 => \N__51374\,
            in2 => \N__51068\,
            in3 => \N__79320\,
            lcout => m65_ns,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_RNIGQ8J_4_LC_21_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__55294\,
            in1 => \N__55155\,
            in2 => \_gnd_net_\,
            in3 => \N__55138\,
            lcout => \CONTROL.programCounter_ret_19_RNIGQ8JZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m58_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001101101"
        )
    port map (
            in0 => \N__77150\,
            in1 => \N__78686\,
            in2 => \N__75962\,
            in3 => \N__77795\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m64_am_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__76321\,
            in1 => \_gnd_net_\,
            in2 => \N__51377\,
            in3 => \N__55196\,
            lcout => \PROM.ROMDATA.m64_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m45_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101110001"
        )
    port map (
            in0 => \N__77149\,
            in1 => \N__78685\,
            in2 => \N__75961\,
            in3 => \N__77793\,
            lcout => \PROM.ROMDATA.m45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNID1RPI_14_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011101000"
        )
    port map (
            in0 => \N__63116\,
            in1 => \N__74860\,
            in2 => \N__63848\,
            in3 => \N__56741\,
            lcout => \ALU.log_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_20_0_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011101000"
        )
    port map (
            in0 => \N__63114\,
            in1 => \N__66314\,
            in2 => \N__74886\,
            in3 => \N__68943\,
            lcout => \ALU.status_8_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_14_0_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__51359\,
            in1 => \N__51344\,
            in2 => \N__51323\,
            in3 => \N__51295\,
            lcout => OPEN,
            ltout => \ALU.status_8_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_7_0_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__51263\,
            in1 => \N__51242\,
            in2 => \N__51206\,
            in3 => \N__51179\,
            lcout => \ALU.status_8_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_19_0_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110110010"
        )
    port map (
            in0 => \N__63115\,
            in1 => \N__53048\,
            in2 => \N__74887\,
            in3 => \N__74607\,
            lcout => OPEN,
            ltout => \ALU.log_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_15_0_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__57248\,
            in1 => \N__51188\,
            in2 => \N__51182\,
            in3 => \N__57514\,
            lcout => \ALU.status_8_13_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIV5AOK_13_LC_22_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011101000"
        )
    port map (
            in0 => \N__63301\,
            in1 => \N__61009\,
            in2 => \N__74826\,
            in3 => \N__56829\,
            lcout => \ALU.c_RNIV5AOKZ0Z_13\,
            ltout => \ALU.c_RNIV5AOKZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIO5N04A_0_13_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__70198\,
            in1 => \N__58533\,
            in2 => \N__51554\,
            in3 => \N__51502\,
            lcout => \ALU.c_RNIO5N04A_0Z0Z_13\,
            ltout => \ALU.c_RNIO5N04A_0Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_13_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67432\,
            in2 => \N__51551\,
            in3 => \N__67388\,
            lcout => \ALU.bZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73158\,
            ce => \N__67942\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNIO5N04A_13_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__70199\,
            in1 => \N__51515\,
            in2 => \N__51509\,
            in3 => \N__58534\,
            lcout => \ALU.c_RNIO5N04AZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_13_0_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011101000"
        )
    port map (
            in0 => \N__63299\,
            in1 => \N__61008\,
            in2 => \N__74825\,
            in3 => \N__56828\,
            lcout => OPEN,
            ltout => \ALU.N_16_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_6_0_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__51490\,
            in1 => \_gnd_net_\,
            in2 => \N__51461\,
            in3 => \N__51443\,
            lcout => \ALU.status_8_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_12_0_LC_22_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101110010010"
        )
    port map (
            in0 => \N__63298\,
            in1 => \N__62939\,
            in2 => \N__74824\,
            in3 => \N__62887\,
            lcout => \ALU.log_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI7KS2I_9_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001110000110"
        )
    port map (
            in0 => \N__62888\,
            in1 => \N__74771\,
            in2 => \N__62949\,
            in3 => \N__63300\,
            lcout => \ALU.d_RNI7KS2IZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.e_12_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__67743\,
            in2 => \N__67602\,
            in3 => \N__67655\,
            lcout => \ALU.eZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73164\,
            ce => \N__69245\,
            sr => \_gnd_net_\
        );

    \ALU.e_13_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__67494\,
            in1 => \N__67442\,
            in2 => \_gnd_net_\,
            in3 => \N__67392\,
            lcout => \ALU.eZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73164\,
            ce => \N__69245\,
            sr => \_gnd_net_\
        );

    \ALU.e_14_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__68137\,
            in1 => \N__68057\,
            in2 => \_gnd_net_\,
            in3 => \N__68004\,
            lcout => \ALU.eZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73164\,
            ce => \N__69245\,
            sr => \_gnd_net_\
        );

    \ALU.g_12_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67741\,
            in1 => \N__67668\,
            in2 => \_gnd_net_\,
            in3 => \N__67595\,
            lcout => g_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73175\,
            ce => \N__70993\,
            sr => \_gnd_net_\
        );

    \ALU.g_13_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67455\,
            in1 => \N__67512\,
            in2 => \_gnd_net_\,
            in3 => \N__67400\,
            lcout => g_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73175\,
            ce => \N__70993\,
            sr => \_gnd_net_\
        );

    \ALU.g_14_LC_22_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__68138\,
            in1 => \N__68086\,
            in2 => \_gnd_net_\,
            in3 => \N__68001\,
            lcout => g_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73175\,
            ce => \N__70993\,
            sr => \_gnd_net_\
        );

    \ALU.d_1_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__59305\,
            in1 => \N__69690\,
            in2 => \N__52247\,
            in3 => \N__68989\,
            lcout => \ALU.dZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73186\,
            ce => \N__70250\,
            sr => \_gnd_net_\
        );

    \ALU.d_0_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__69156\,
            in1 => \N__52124\,
            in2 => \N__69715\,
            in3 => \N__52053\,
            lcout => \ALU.dZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73186\,
            ce => \N__70250\,
            sr => \_gnd_net_\
        );

    \ALU.d_7_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010101100100"
        )
    port map (
            in0 => \N__58864\,
            in1 => \N__67254\,
            in2 => \N__51938\,
            in3 => \N__51862\,
            lcout => \ALU.dZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73186\,
            ce => \N__70250\,
            sr => \_gnd_net_\
        );

    \ALU.d_8_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67252\,
            in1 => \N__51778\,
            in2 => \N__51722\,
            in3 => \N__51635\,
            lcout => \ALU.dZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73186\,
            ce => \N__70250\,
            sr => \_gnd_net_\
        );

    \ALU.d_15_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000011101111"
        )
    port map (
            in0 => \N__53008\,
            in1 => \N__67253\,
            in2 => \N__59142\,
            in3 => \N__52935\,
            lcout => \ALU.dZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73186\,
            ce => \N__70250\,
            sr => \_gnd_net_\
        );

    \ALU.d_9_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__52870\,
            in1 => \N__66806\,
            in2 => \N__58564\,
            in3 => \N__52788\,
            lcout => \ALU.dZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73186\,
            ce => \N__70250\,
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPFFDD1_0_6_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__66766\,
            in1 => \N__62583\,
            in2 => \N__59645\,
            in3 => \N__66074\,
            lcout => OPEN,
            ltout => \ALU.d_RNIPFFDD1_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIBTSVI3_6_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__52709\,
            in1 => \_gnd_net_\,
            in2 => \N__52691\,
            in3 => \N__52493\,
            lcout => \ALU.N_863\,
            ltout => \ALU.N_863_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIGPBNB6_2_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__68935\,
            in1 => \_gnd_net_\,
            in2 => \N__52688\,
            in3 => \N__68174\,
            lcout => OPEN,
            ltout => \ALU.d_RNIGPBNB6Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIUDSOL9_2_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52683\,
            in2 => \N__52640\,
            in3 => \N__52499\,
            lcout => \ALU.a_15_m0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNINGV0T2_15_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__68934\,
            in1 => \N__69973\,
            in2 => \N__68556\,
            in3 => \N__52527\,
            lcout => \ALU.c_RNINGV0T2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIPFFDD1_6_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__66073\,
            in1 => \N__59640\,
            in2 => \N__62588\,
            in3 => \N__66765\,
            lcout => \ALU.d_RNIPFFDD1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_16_0_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60358\,
            in2 => \_gnd_net_\,
            in3 => \N__60319\,
            lcout => OPEN,
            ltout => \ALU.status_14_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_8_0_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__60280\,
            in1 => \N__59929\,
            in2 => \N__53363\,
            in3 => \N__61753\,
            lcout => \ALU.status_14_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_10_0_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__62338\,
            in1 => \N__62047\,
            in2 => \_gnd_net_\,
            in3 => \N__61492\,
            lcout => OPEN,
            ltout => \ALU.status_14_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_4_0_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__53036\,
            in1 => \N__63699\,
            in2 => \N__53345\,
            in3 => \N__63512\,
            lcout => \ALU.status_14_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIHLMGP_14_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__61014\,
            in1 => \N__63774\,
            in2 => \_gnd_net_\,
            in3 => \N__66736\,
            lcout => \ALU.N_979\,
            ltout => \ALU.N_979_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIUMNP22_15_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__63639\,
            in1 => \N__66742\,
            in2 => \N__53309\,
            in3 => \N__66076\,
            lcout => \ALU.N_968\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_22_0_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__53762\,
            in1 => \N__63638\,
            in2 => \N__63274\,
            in3 => \N__53177\,
            lcout => \ALU.status_RNO_22Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_9_0_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__59665\,
            in1 => \N__59353\,
            in2 => \_gnd_net_\,
            in3 => \N__66856\,
            lcout => \ALU.status_14_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIVHVMK_13_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__63225\,
            in1 => \N__61018\,
            in2 => \N__56839\,
            in3 => \_gnd_net_\,
            lcout => \ALU.c_RNIVHVMKZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_17_I_21_c_RNO_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__56719\,
            in1 => \N__63778\,
            in2 => \N__63613\,
            in3 => \N__74570\,
            lcout => \ALU.status_17_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIDDGOI_14_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__63779\,
            in1 => \N__63240\,
            in2 => \_gnd_net_\,
            in3 => \N__56718\,
            lcout => \ALU.c_RNIDDGOIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_e_0_RNO_0_2_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__69519\,
            in1 => \N__53690\,
            in2 => \_gnd_net_\,
            in3 => \N__63516\,
            lcout => OPEN,
            ltout => \ALU.status_e_0_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_e_0_2_LC_22_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56543\,
            in2 => \N__53732\,
            in3 => \N__53726\,
            lcout => \aluStatus_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73208\,
            ce => \N__56603\,
            sr => \_gnd_net_\
        );

    \ALU.c_RNI0NMSH_15_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__63241\,
            in1 => \_gnd_net_\,
            in2 => \N__63614\,
            in3 => \N__74569\,
            lcout => \ALU.c_RNI0NMSHZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_e_0_RNO_2_2_LC_22_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010001000"
        )
    port map (
            in0 => \N__74571\,
            in1 => \N__74856\,
            in2 => \_gnd_net_\,
            in3 => \N__63582\,
            lcout => OPEN,
            ltout => \ALU.N_570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_e_0_RNO_1_2_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__63242\,
            in1 => \_gnd_net_\,
            in2 => \N__53729\,
            in3 => \N__74528\,
            lcout => \ALU.status_e_0_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.g3_0_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__53689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53669\,
            lcout => \CONTROL.g3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_RNI9NEO1_15_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__53611\,
            in1 => \N__53588\,
            in2 => \N__53517\,
            in3 => \N__53478\,
            lcout => OPEN,
            ltout => \ALU.operand2_6_ns_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIKIDM2_15_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__54186\,
            in1 => \N__54328\,
            in2 => \N__53438\,
            in3 => \N__53434\,
            lcout => \ALU.N_1260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIILK02_15_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000011"
        )
    port map (
            in0 => \N__54329\,
            in1 => \N__54317\,
            in2 => \N__54308\,
            in3 => \N__54187\,
            lcout => OPEN,
            ltout => \ALU.N_1148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI2SRO3_15_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54161\,
            in2 => \N__54146\,
            in3 => \N__54140\,
            lcout => \aluOut_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI8VV95_15_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53990\,
            in1 => \N__53984\,
            in2 => \_gnd_net_\,
            in3 => \N__53968\,
            lcout => OPEN,
            ltout => \ALU.c_RNI8VV95Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIJTKD7_15_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53783\,
            in2 => \N__53765\,
            in3 => \N__71463\,
            lcout => \ALU.c_RNIJTKD7Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m320_bm_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010001000"
        )
    port map (
            in0 => \N__78776\,
            in1 => \N__77993\,
            in2 => \N__75965\,
            in3 => \N__77304\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m320_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m320_ns_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54401\,
            in2 => \N__53744\,
            in3 => \N__76475\,
            lcout => \PROM.ROMDATA.m320_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m413_am_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000011"
        )
    port map (
            in0 => \N__78774\,
            in1 => \N__77989\,
            in2 => \N__75964\,
            in3 => \N__77302\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m413_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m414_ns_1_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__79874\,
            in1 => \N__53741\,
            in2 => \N__53735\,
            in3 => \N__76474\,
            lcout => \PROM.ROMDATA.m414_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_2_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__54821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONTROL.dout_reto_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.un1_busState97_i_i_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__54782\,
            in1 => \N__54770\,
            in2 => \N__54752\,
            in3 => \N__54685\,
            lcout => \CONTROL.N_45_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m139_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__78773\,
            in1 => \N__77988\,
            in2 => \_gnd_net_\,
            in3 => \N__77301\,
            lcout => \PROM.ROMDATA.m139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m320_am_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000110010"
        )
    port map (
            in0 => \N__77303\,
            in1 => \N__75839\,
            in2 => \N__78054\,
            in3 => \N__78775\,
            lcout => \PROM.ROMDATA.m320_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m154_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110100000000"
        )
    port map (
            in0 => \N__75831\,
            in1 => \N__54395\,
            in2 => \N__64286\,
            in3 => \N__74061\,
            lcout => \PROM.ROMDATA.N_558_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m323_bm_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__78736\,
            in1 => \N__75832\,
            in2 => \N__79048\,
            in3 => \N__77982\,
            lcout => \PROM.ROMDATA.m323_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m49_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010101111"
        )
    port map (
            in0 => \N__77165\,
            in1 => \_gnd_net_\,
            in2 => \N__78049\,
            in3 => \N__78735\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m228_bm_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55222\,
            in2 => \N__54374\,
            in3 => \N__75830\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m228_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m229_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000100100010"
        )
    port map (
            in0 => \N__79842\,
            in1 => \N__54371\,
            in2 => \N__54365\,
            in3 => \N__76473\,
            lcout => \PROM.ROMDATA.m229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m226_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000100010"
        )
    port map (
            in0 => \N__78734\,
            in1 => \N__77977\,
            in2 => \_gnd_net_\,
            in3 => \N__77164\,
            lcout => \PROM.ROMDATA.m226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m312_bm_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__77981\,
            in1 => \N__73905\,
            in2 => \N__75963\,
            in3 => \N__78737\,
            lcout => \PROM.ROMDATA.m312_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m437_ns_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011010001"
        )
    port map (
            in0 => \N__54836\,
            in1 => \N__76460\,
            in2 => \N__64442\,
            in3 => \N__77121\,
            lcout => \PROM.ROMDATA.m437_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m11_bm_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101111001"
        )
    port map (
            in0 => \N__77118\,
            in1 => \N__75645\,
            in2 => \N__77973\,
            in3 => \N__78330\,
            lcout => \PROM.ROMDATA.m11_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m118_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101100011110"
        )
    port map (
            in0 => \N__78329\,
            in1 => \N__77796\,
            in2 => \N__75887\,
            in3 => \N__77117\,
            lcout => \PROM.ROMDATA.m118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m312_ns_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__76461\,
            in1 => \N__54857\,
            in2 => \_gnd_net_\,
            in3 => \N__54851\,
            lcout => \PROM.ROMDATA.m312_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m437_ns_1_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001111101"
        )
    port map (
            in0 => \N__78332\,
            in1 => \N__77803\,
            in2 => \N__75888\,
            in3 => \N__77120\,
            lcout => \PROM.ROMDATA.m437_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m18_bm_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011100001"
        )
    port map (
            in0 => \N__77119\,
            in1 => \N__75646\,
            in2 => \N__77974\,
            in3 => \N__78331\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m18_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m19_ns_1_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100110011"
        )
    port map (
            in0 => \N__54830\,
            in1 => \N__79841\,
            in2 => \N__54824\,
            in3 => \N__76458\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m19_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m19_ns_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101001010"
        )
    port map (
            in0 => \N__76459\,
            in1 => \N__54956\,
            in2 => \N__54944\,
            in3 => \N__54941\,
            lcout => \PROM.ROMDATA.m19_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m111_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101011010"
        )
    port map (
            in0 => \N__76911\,
            in1 => \N__78323\,
            in2 => \N__77838\,
            in3 => \N__75423\,
            lcout => \PROM.ROMDATA.m111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m117_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001111001111"
        )
    port map (
            in0 => \N__78321\,
            in1 => \N__77575\,
            in2 => \N__75709\,
            in3 => \N__76909\,
            lcout => \PROM.ROMDATA.m117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m33_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110110"
        )
    port map (
            in0 => \N__76913\,
            in1 => \N__78324\,
            in2 => \N__77839\,
            in3 => \N__75424\,
            lcout => \PROM.ROMDATA.m33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m211_ns_N_2L1_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100100011000"
        )
    port map (
            in0 => \N__78322\,
            in1 => \N__76173\,
            in2 => \N__75710\,
            in3 => \N__76910\,
            lcout => \PROM.ROMDATA.m211_ns_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIJA5J_1_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55064\,
            in1 => \N__54902\,
            in2 => \_gnd_net_\,
            in3 => \N__54890\,
            lcout => \N_416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNIH68I_1_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__54889\,
            in1 => \N__73787\,
            in2 => \_gnd_net_\,
            in3 => \N__55139\,
            lcout => OPEN,
            ltout => \CONTROL.programCounter_ret_1_RNIH68IZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_fast_RNI1RBH1_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55055\,
            in2 => \N__54875\,
            in3 => \N__54872\,
            lcout => \progRomAddress_1\,
            ltout => \progRomAddress_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m114_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100111010101"
        )
    port map (
            in0 => \N__75422\,
            in1 => \N__77576\,
            in2 => \N__54866\,
            in3 => \N__76912\,
            lcout => \PROM.ROMDATA.m114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m492_am_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100000000"
        )
    port map (
            in0 => \N__73542\,
            in1 => \N__73811\,
            in2 => \N__73741\,
            in3 => \N__77700\,
            lcout => \PROM.ROMDATA.m492_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m55_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000010010"
        )
    port map (
            in0 => \N__77073\,
            in1 => \N__75817\,
            in2 => \N__77895\,
            in3 => \N__78339\,
            lcout => \PROM.ROMDATA.m55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_RNINC8I_4_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__55184\,
            in1 => \N__55169\,
            in2 => \_gnd_net_\,
            in3 => \N__55137\,
            lcout => OPEN,
            ltout => \CONTROL.programCounter_ret_1_RNINC8IZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_18_fast_RNID7CH1_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55058\,
            in2 => \N__55013\,
            in3 => \N__55010\,
            lcout => \progRomAddress_4\,
            ltout => \progRomAddress_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m147_bm_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54998\,
            in2 => \N__54992\,
            in3 => \N__54989\,
            lcout => \PROM.ROMDATA.m147_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m140_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111101001"
        )
    port map (
            in0 => \N__77072\,
            in1 => \N__75816\,
            in2 => \N__77894\,
            in3 => \N__78338\,
            lcout => \PROM.ROMDATA.m140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m156_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__78337\,
            in1 => \N__77693\,
            in2 => \_gnd_net_\,
            in3 => \N__77071\,
            lcout => \PROM.ROMDATA.m156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m92_bm_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__54980\,
            in1 => \N__65183\,
            in2 => \_gnd_net_\,
            in3 => \N__76286\,
            lcout => \PROM.ROMDATA.m92_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m183_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011010011100"
        )
    port map (
            in0 => \N__64642\,
            in1 => \N__76264\,
            in2 => \N__64531\,
            in3 => \N__64485\,
            lcout => \PROM.ROMDATA.m183\,
            ltout => \PROM.ROMDATA.m183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m185_bm_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55244\,
            in2 => \N__55256\,
            in3 => \N__64919\,
            lcout => \PROM.ROMDATA.m185_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m166_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__76930\,
            in1 => \N__78790\,
            in2 => \N__77841\,
            in3 => \N__75631\,
            lcout => \PROM.ROMDATA.N_525_mux\,
            ltout => \PROM.ROMDATA.N_525_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m427_bm_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__75635\,
            in1 => \N__64017\,
            in2 => \N__55247\,
            in3 => \N__76287\,
            lcout => \PROM.ROMDATA.m427_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m164_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000001"
        )
    port map (
            in0 => \N__76929\,
            in1 => \N__78789\,
            in2 => \N__77840\,
            in3 => \N__75630\,
            lcout => \PROM.ROMDATA.m164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m132_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000101111"
        )
    port map (
            in0 => \N__78791\,
            in1 => \N__77590\,
            in2 => \N__75885\,
            in3 => \N__76931\,
            lcout => \PROM.ROMDATA.m132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m492_bm_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110001"
        )
    port map (
            in0 => \N__73553\,
            in1 => \N__64862\,
            in2 => \N__73742\,
            in3 => \N__73810\,
            lcout => \PROM.ROMDATA.m492_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m133_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__78788\,
            in1 => \N__77583\,
            in2 => \_gnd_net_\,
            in3 => \N__76928\,
            lcout => \PROM.ROMDATA.m133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m182_LC_22_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000010"
        )
    port map (
            in0 => \N__77145\,
            in1 => \N__76291\,
            in2 => \N__77975\,
            in3 => \N__78795\,
            lcout => \PROM.ROMDATA.i4_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m338_bm_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__55238\,
            in1 => \N__75828\,
            in2 => \_gnd_net_\,
            in3 => \N__55226\,
            lcout => \PROM.ROMDATA.m338_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m92_am_1_LC_22_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011101110010"
        )
    port map (
            in0 => \N__77147\,
            in1 => \N__76292\,
            in2 => \N__77976\,
            in3 => \N__75688\,
            lcout => \PROM.ROMDATA.m92_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m158_LC_22_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__78797\,
            in1 => \N__77816\,
            in2 => \N__75902\,
            in3 => \N__77148\,
            lcout => \PROM.ROMDATA.m158\,
            ltout => \PROM.ROMDATA.m158_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m162_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__79838\,
            in1 => \N__76293\,
            in2 => \N__55484\,
            in3 => \N__64925\,
            lcout => \PROM.ROMDATA.m162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m135_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010010000"
        )
    port map (
            in0 => \N__78796\,
            in1 => \N__77812\,
            in2 => \N__75901\,
            in3 => \N__77146\,
            lcout => \PROM.ROMDATA.m135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m202_LC_22_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__74065\,
            in1 => \N__72731\,
            in2 => \N__64142\,
            in3 => \N__55481\,
            lcout => \PROM_ROMDATA_dintern_6ro\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m317_am_LC_22_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100101100010"
        )
    port map (
            in0 => \N__78798\,
            in1 => \N__75829\,
            in2 => \N__73891\,
            in3 => \N__78989\,
            lcout => \PROM.ROMDATA.m317_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_19_4_LC_22_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55333\,
            lcout => \CONTROL.dout_reto_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_0_c_inv_LC_23_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66772\,
            in2 => \N__55283\,
            in3 => \N__60579\,
            lcout => \ALU.aluOut_i_0\,
            ltout => OPEN,
            carryin => \bfn_23_7_0_\,
            carryout => \ALU.status_19_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_1_c_inv_LC_23_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66084\,
            in2 => \N__55274\,
            in3 => \N__65537\,
            lcout => \ALU.aluOut_i_1\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_0\,
            carryout => \ALU.status_19_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_2_c_inv_LC_23_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68945\,
            in2 => \N__55265\,
            in3 => \N__66320\,
            lcout => \ALU.aluOut_i_2\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_1\,
            carryout => \ALU.status_19_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_3_c_inv_LC_23_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68525\,
            in2 => \N__56426\,
            in3 => \N__60266\,
            lcout => \ALU.aluOut_i_3\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_2\,
            carryout => \ALU.status_19_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_4_c_inv_LC_23_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56417\,
            in2 => \N__56285\,
            in3 => \N__59883\,
            lcout => \ALU.aluOut_i_4\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_3\,
            carryout => \ALU.status_19_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_5_c_inv_LC_23_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56276\,
            in2 => \N__56150\,
            in3 => \N__59644\,
            lcout => \ALU.aluOut_i_5\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_4\,
            carryout => \ALU.status_19_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_6_c_inv_LC_23_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56131\,
            in2 => \N__56003\,
            in3 => \N__62550\,
            lcout => \ALU.aluOut_i_6\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_5\,
            carryout => \ALU.status_19_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_7_c_inv_LC_23_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55991\,
            in2 => \N__55835\,
            in3 => \N__62298\,
            lcout => \ALU.aluOut_i_7\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_6\,
            carryout => \ALU.status_19_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_8_c_inv_LC_23_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55822\,
            in2 => \N__55697\,
            in3 => \N__62024\,
            lcout => \ALU.aluOut_i_8\,
            ltout => OPEN,
            carryin => \bfn_23_8_0_\,
            carryout => \ALU.status_19_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_9_c_inv_LC_23_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55687\,
            in2 => \N__55598\,
            in3 => \N__62889\,
            lcout => \ALU.aluOut_i_9\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_8\,
            carryout => \ALU.status_19_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_10_c_inv_LC_23_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55589\,
            in2 => \N__55517\,
            in3 => \N__61701\,
            lcout => \ALU.aluOut_i_10\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_9\,
            carryout => \ALU.status_19_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_11_c_inv_LC_23_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__61475\,
            in1 => \N__57053\,
            in2 => \N__56942\,
            in3 => \_gnd_net_\,
            lcout => \ALU.aluOut_i_11\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_10\,
            carryout => \ALU.status_19_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_12_c_inv_LC_23_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56933\,
            in2 => \N__56852\,
            in3 => \N__61226\,
            lcout => \ALU.aluOut_i_12\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_11\,
            carryout => \ALU.status_19_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_13_c_inv_LC_23_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56759\,
            in2 => \N__56843\,
            in3 => \N__61011\,
            lcout => \ALU.aluOut_i_13\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_12\,
            carryout => \ALU.status_19_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_14_c_inv_LC_23_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56749\,
            in2 => \N__56678\,
            in3 => \N__63852\,
            lcout => \ALU.aluOut_i_14\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_13\,
            carryout => \ALU.status_19_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_19_cry_15_c_inv_LC_23_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__63640\,
            in1 => \N__74603\,
            in2 => \N__56669\,
            in3 => \_gnd_net_\,
            lcout => \ALU.aluOut_i_15\,
            ltout => OPEN,
            carryin => \ALU.status_19_cry_14\,
            carryout => \ALU.status_19Z0Z_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_5_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__69513\,
            in1 => \N__56622\,
            in2 => \N__56647\,
            in3 => \N__56660\,
            lcout => \aluStatus_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_1_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__56621\,
            in1 => \N__63414\,
            in2 => \N__56542\,
            in3 => \N__63389\,
            lcout => \aluStatus_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI12L8C5_2_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__56492\,
            in1 => \N__68524\,
            in2 => \N__56472\,
            in3 => \N__68944\,
            lcout => \ALU.d_RNI12L8C5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_18_0_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011101000"
        )
    port map (
            in0 => \N__63113\,
            in1 => \N__60265\,
            in2 => \N__74902\,
            in3 => \N__68523\,
            lcout => \ALU.log_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_12_c_RNIP50IR3_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111110111"
        )
    port map (
            in0 => \N__57242\,
            in1 => \N__68565\,
            in2 => \N__67243\,
            in3 => \N__60835\,
            lcout => OPEN,
            ltout => \ALU.a_15_d_ns_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_558_c_RNIB75F9G_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100101110"
        )
    port map (
            in0 => \N__57185\,
            in1 => \N__57121\,
            in2 => \N__57176\,
            in3 => \N__67183\,
            lcout => \ALU.mult_558_c_RNIB75F9GZ0\,
            ltout => \ALU.mult_558_c_RNIB75F9GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_13_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__67493\,
            in1 => \_gnd_net_\,
            in2 => \N__57173\,
            in3 => \N__67450\,
            lcout => \ALU.aZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73165\,
            ce => \N__71214\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_d_s_10_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__59136\,
            in1 => \N__67179\,
            in2 => \_gnd_net_\,
            in3 => \N__69908\,
            lcout => \ALU.a_15_d_sZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJ7J1M5_0_2_LC_23_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__59159\,
            in1 => \N__57109\,
            in2 => \N__57122\,
            in3 => \N__57073\,
            lcout => \ALU.d_RNIJ7J1M5_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_m3_d_s_8_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__69907\,
            lcout => \ALU.a_15_m3_d_sZ0Z_8\,
            ltout => \ALU.a_15_m3_d_sZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIJ7J1M5_2_LC_23_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100001011"
        )
    port map (
            in0 => \N__59158\,
            in1 => \N__57110\,
            in2 => \N__57077\,
            in3 => \N__57074\,
            lcout => \ALU.d_RNIJ7J1M5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.f_12_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67754\,
            in1 => \N__67672\,
            in2 => \_gnd_net_\,
            in3 => \N__67603\,
            lcout => f_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73176\,
            ce => \N__67864\,
            sr => \_gnd_net_\
        );

    \ALU.f_13_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67449\,
            in1 => \N__67504\,
            in2 => \_gnd_net_\,
            in3 => \N__67390\,
            lcout => f_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73176\,
            ce => \N__67864\,
            sr => \_gnd_net_\
        );

    \ALU.f_14_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__68058\,
            in1 => \N__68123\,
            in2 => \_gnd_net_\,
            in3 => \N__68000\,
            lcout => f_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73176\,
            ce => \N__67864\,
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_13_c_RNIBVHEA1_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100011"
        )
    port map (
            in0 => \N__63701\,
            in1 => \N__59287\,
            in2 => \N__67270\,
            in3 => \N__57523\,
            lcout => \ALU.addsub_cry_13_c_RNIBVHEAZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_13_c_RNIBVHEA1_0_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__59288\,
            in1 => \N__67248\,
            in2 => \N__57527\,
            in3 => \N__63700\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_13_c_RNIBVHEA1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_13_c_RNIJMTGA5_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57503\,
            in2 => \N__57488\,
            in3 => \N__57485\,
            lcout => OPEN,
            ltout => \ALU.addsub_cry_13_c_RNIJMTGAZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.mult_561_c_RNI1EB5TL_LC_23_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__59107\,
            in1 => \N__67251\,
            in2 => \N__57479\,
            in3 => \N__57476\,
            lcout => \ALU.a_15_ns_rn_0_14\,
            ltout => \ALU.a_15_ns_rn_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_14_LC_23_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68122\,
            in2 => \N__57461\,
            in3 => \N__68087\,
            lcout => \ALU.aZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73187\,
            ce => \N__71200\,
            sr => \_gnd_net_\
        );

    \ALU.a_15_s_3_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__59286\,
            in1 => \N__59102\,
            in2 => \_gnd_net_\,
            in3 => \N__67244\,
            lcout => \ALU.a_15_sZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.a_15_ns_sn_14_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__67249\,
            in1 => \N__59106\,
            in2 => \_gnd_net_\,
            in3 => \N__59339\,
            lcout => \ALU.a_15_ns_snZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_6_c_RNIJ7U2L_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111001101"
        )
    port map (
            in0 => \N__59289\,
            in1 => \N__67250\,
            in2 => \N__59138\,
            in3 => \N__62048\,
            lcout => \ALU.a_15_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.h_3_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58817\,
            in2 => \N__58756\,
            in3 => \N__58677\,
            lcout => h_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73193\,
            ce => \N__69451\,
            sr => \_gnd_net_\
        );

    \ALU.h_10_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58562\,
            in1 => \N__58372\,
            in2 => \_gnd_net_\,
            in3 => \N__58301\,
            lcout => h_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73193\,
            ce => \N__69451\,
            sr => \_gnd_net_\
        );

    \ALU.h_11_LC_23_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58195\,
            in2 => \N__58127\,
            in3 => \N__58056\,
            lcout => h_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73193\,
            ce => \N__69451\,
            sr => \_gnd_net_\
        );

    \ALU.h_12_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67755\,
            in1 => \N__67687\,
            in2 => \_gnd_net_\,
            in3 => \N__67617\,
            lcout => h_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73193\,
            ce => \N__69451\,
            sr => \_gnd_net_\
        );

    \ALU.h_13_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67460\,
            in1 => \N__67517\,
            in2 => \_gnd_net_\,
            in3 => \N__67399\,
            lcout => h_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73193\,
            ce => \N__69451\,
            sr => \_gnd_net_\
        );

    \ALU.h_14_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__68078\,
            in1 => \N__68139\,
            in2 => \_gnd_net_\,
            in3 => \N__68002\,
            lcout => h_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73193\,
            ce => \N__69451\,
            sr => \_gnd_net_\
        );

    \CONTROL.addrstackptr_RNI0D361_4_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__57801\,
            in1 => \_gnd_net_\,
            in2 => \N__60818\,
            in3 => \N__60736\,
            lcout => \CONTROL.g1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_0_c_THRU_CRY_0_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63276\,
            in2 => \N__63297\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_23_14_0_\,
            carryout => \ALU.addsub_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI4KF5H_0_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60625\,
            in2 => \N__60386\,
            in3 => \N__60347\,
            lcout => \ALU.addsub_0\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_0_c_THRU_CO\,
            carryout => \ALU.addsub_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_0_c_RNISBATS_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65536\,
            in2 => \N__60344\,
            in3 => \N__60308\,
            lcout => \ALU.addsub_1\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_0\,
            carryout => \ALU.addsub_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_1_c_RNIRBVRO_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66303\,
            in2 => \N__60305\,
            in3 => \N__60269\,
            lcout => \ALU.addsub_2\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_1\,
            carryout => \ALU.addsub_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_2_c_RNIDOASJ_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60236\,
            in2 => \N__59957\,
            in3 => \N__59915\,
            lcout => \ALU.addsub_3\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_2\,
            carryout => \ALU.addsub_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_3_c_RNI67KIM_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59882\,
            in2 => \N__59693\,
            in3 => \N__59648\,
            lcout => \ALU.addsub_4\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_3\,
            carryout => \ALU.addsub_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_4_c_RNIDE0RM_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59639\,
            in2 => \N__59384\,
            in3 => \N__59342\,
            lcout => \ALU.addsub_5\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_4\,
            carryout => \ALU.addsub_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_5_c_RNIR5MEM_LC_23_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62586\,
            in2 => \N__62366\,
            in3 => \N__62327\,
            lcout => \ALU.addsub_6\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_5\,
            carryout => \ALU.addsub_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_6_c_RNI112DK_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62219\,
            in2 => \N__62060\,
            in3 => \N__62030\,
            lcout => \ALU.addsub_7\,
            ltout => OPEN,
            carryin => \bfn_23_15_0_\,
            carryout => \ALU.addsub_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_7_c_RNI7LOOL_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62027\,
            in2 => \N__61781\,
            in3 => \N__61742\,
            lcout => \ALU.addsub_8\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_7\,
            carryout => \ALU.addsub_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_8_c_RNINRS3M_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62801\,
            in2 => \N__62672\,
            in3 => \N__61739\,
            lcout => \ALU.addsub_9\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_8\,
            carryout => \ALU.addsub_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_9_c_RNI8MSRO_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61736\,
            in2 => \N__61710\,
            in3 => \N__61478\,
            lcout => \ALU.addsub_10\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_9\,
            carryout => \ALU.addsub_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_10_c_RNIS0BKM_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61364\,
            in2 => \N__61298\,
            in3 => \N__61247\,
            lcout => \ALU.addsub_11\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_10\,
            carryout => \ALU.addsub_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_11_c_RNI0C50P_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61244\,
            in2 => \N__61224\,
            in3 => \N__61028\,
            lcout => \ALU.addsub_12\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_11\,
            carryout => \ALU.addsub_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_12_c_RNIEV1GP_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61025\,
            in2 => \N__61019\,
            in3 => \N__63863\,
            lcout => \ALU.addsub_13\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_12\,
            carryout => \ALU.addsub_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_13_c_RNI9HJ8N_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63860\,
            in2 => \N__63819\,
            in3 => \N__63683\,
            lcout => \ALU.addsub_14\,
            ltout => OPEN,
            carryin => \ALU.addsub_cry_13\,
            carryout => \ALU.addsub_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_14_c_RNIORHUL_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63680\,
            in2 => \N__63612\,
            in3 => \N__63488\,
            lcout => \ALU.addsub_15\,
            ltout => OPEN,
            carryin => \bfn_23_16_0_\,
            carryout => \ALU.addsub_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.status_RNO_0_1_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__63442\,
            in1 => \N__63239\,
            in2 => \N__69496\,
            in3 => \N__63392\,
            lcout => \ALU.N_545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIPBAG72_14_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__69988\,
            in1 => \N__63360\,
            in2 => \_gnd_net_\,
            in3 => \N__62627\,
            lcout => \ALU.c_RNIPBAG72Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI70I1I_9_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__63238\,
            in1 => \N__62927\,
            in2 => \_gnd_net_\,
            in3 => \N__62881\,
            lcout => \ALU.d_RNI70I1IZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNISS7FV1_14_LC_23_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__62663\,
            in1 => \N__68933\,
            in2 => \_gnd_net_\,
            in3 => \N__66075\,
            lcout => \ALU.N_1029\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m500_ns_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010011101100"
        )
    port map (
            in0 => \N__79497\,
            in1 => \N__62621\,
            in2 => \N__63935\,
            in3 => \N__63869\,
            lcout => \PROM.ROMDATA.m500_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m498_am_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100111"
        )
    port map (
            in0 => \N__75995\,
            in1 => \N__78997\,
            in2 => \N__73919\,
            in3 => \N__78744\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m498_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m498_ns_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63950\,
            in2 => \N__63938\,
            in3 => \N__76572\,
            lcout => \PROM.ROMDATA.m498_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m317_bm_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010101100"
        )
    port map (
            in0 => \N__75996\,
            in1 => \N__78745\,
            in2 => \N__73918\,
            in3 => \N__78041\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m317_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m317_ns_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__63926\,
            in1 => \_gnd_net_\,
            in2 => \N__63914\,
            in3 => \N__76573\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m317_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m325_ns_1_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__63911\,
            in1 => \N__79498\,
            in2 => \N__63899\,
            in3 => \N__79895\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m325_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m325_ns_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__79499\,
            in1 => \N__74912\,
            in2 => \N__63896\,
            in3 => \N__63893\,
            lcout => \PROM.ROMDATA.m325_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m329_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__74070\,
            in1 => \N__72770\,
            in2 => \N__63884\,
            in3 => \N__64124\,
            lcout => OPEN,
            ltout => \PROM_ROMDATA_dintern_14ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.results_1_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__70882\,
            in1 => \N__64084\,
            in2 => \N__63872\,
            in3 => \N__72299\,
            lcout => \aluResults_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.results_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m494_ns_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__73829\,
            in1 => \N__65192\,
            in2 => \N__73469\,
            in3 => \N__76575\,
            lcout => \PROM.ROMDATA.m494_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m414_ns_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100100110001"
        )
    port map (
            in0 => \N__76574\,
            in1 => \N__64187\,
            in2 => \N__64181\,
            in3 => \N__64346\,
            lcout => \PROM.ROMDATA.m414_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m308_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__74069\,
            in1 => \N__74258\,
            in2 => \N__64157\,
            in3 => \N__72771\,
            lcout => OPEN,
            ltout => \PROM_ROMDATA_dintern_13ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.results_0_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__69270\,
            in1 => \N__64083\,
            in2 => \N__64145\,
            in3 => \N__72298\,
            lcout => \aluResults_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.results_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m198_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010010001"
        )
    port map (
            in0 => \N__78404\,
            in1 => \N__77896\,
            in2 => \N__75954\,
            in3 => \N__77252\,
            lcout => \PROM.ROMDATA.m198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m344_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__72697\,
            in1 => \N__74067\,
            in2 => \N__79064\,
            in3 => \N__64123\,
            lcout => OPEN,
            ltout => \PROM_ROMDATA_dintern_15ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.results_2_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__70913\,
            in1 => \N__64085\,
            in2 => \N__64070\,
            in3 => \N__72304\,
            lcout => \aluResults_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.results_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m367_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__65013\,
            in1 => \N__74066\,
            in2 => \N__64067\,
            in3 => \N__75800\,
            lcout => \PROM.ROMDATA.N_564_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m298_bm_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001100101100"
        )
    port map (
            in0 => \N__78406\,
            in1 => \N__77898\,
            in2 => \N__75955\,
            in3 => \N__77255\,
            lcout => \PROM.ROMDATA.m298_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m386_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__74068\,
            in1 => \N__64261\,
            in2 => \N__64018\,
            in3 => \N__75804\,
            lcout => \PROM.ROMDATA.N_565_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m287_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__78405\,
            in1 => \N__77897\,
            in2 => \_gnd_net_\,
            in3 => \N__77253\,
            lcout => \PROM.ROMDATA.m287\,
            ltout => \PROM.ROMDATA.m287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m410_bm_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__77254\,
            in1 => \N__77940\,
            in2 => \N__64349\,
            in3 => \N__75799\,
            lcout => \PROM.ROMDATA.m410_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m66_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111010"
        )
    port map (
            in0 => \N__77250\,
            in1 => \N__75668\,
            in2 => \N__78021\,
            in3 => \N__78359\,
            lcout => \PROM.ROMDATA.m66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m490_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001010000"
        )
    port map (
            in0 => \N__75669\,
            in1 => \N__74963\,
            in2 => \N__64328\,
            in3 => \N__76404\,
            lcout => \PROM.ROMDATA.m490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m446_am_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000001"
        )
    port map (
            in0 => \N__77251\,
            in1 => \N__75672\,
            in2 => \N__78022\,
            in3 => \N__78361\,
            lcout => \PROM.ROMDATA.m446_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m149_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111101110"
        )
    port map (
            in0 => \N__78358\,
            in1 => \N__77899\,
            in2 => \_gnd_net_\,
            in3 => \N__77249\,
            lcout => \PROM.ROMDATA.m149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m120_bm_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__76403\,
            in1 => \N__64277\,
            in2 => \_gnd_net_\,
            in3 => \N__64271\,
            lcout => \PROM.ROMDATA.m120_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m456_ns_1_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__75670\,
            in1 => \N__64793\,
            in2 => \N__79891\,
            in3 => \N__64966\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m456_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m456_ns_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000001010"
        )
    port map (
            in0 => \N__76405\,
            in1 => \N__64250\,
            in2 => \N__64202\,
            in3 => \N__75671\,
            lcout => \PROM.ROMDATA.m456_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m166_e_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010001"
        )
    port map (
            in0 => \N__78360\,
            in1 => \N__64524\,
            in2 => \N__73740\,
            in3 => \N__64486\,
            lcout => \PROM.ROMDATA.m166_e\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m107_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100010111010"
        )
    port map (
            in0 => \N__78482\,
            in1 => \N__77966\,
            in2 => \N__75795\,
            in3 => \N__77244\,
            lcout => \PROM.ROMDATA.m107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m361_am_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111000"
        )
    port map (
            in0 => \N__77245\,
            in1 => \N__75500\,
            in2 => \N__78573\,
            in3 => \N__79033\,
            lcout => \PROM.ROMDATA.m361_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m104_ns_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__75499\,
            in1 => \N__78988\,
            in2 => \N__79043\,
            in3 => \N__64433\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m104_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m109_bm_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64424\,
            in2 => \N__64418\,
            in3 => \N__76272\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m109_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m121_ns_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011000"
        )
    port map (
            in0 => \N__64355\,
            in1 => \N__64415\,
            in2 => \N__64400\,
            in3 => \N__79322\,
            lcout => \PROM.ROMDATA.m121_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m357_bm_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100111100000"
        )
    port map (
            in0 => \N__77246\,
            in1 => \N__75501\,
            in2 => \N__78043\,
            in3 => \N__78483\,
            lcout => \PROM.ROMDATA.m357_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m120_am_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__76271\,
            in1 => \N__64376\,
            in2 => \_gnd_net_\,
            in3 => \N__64370\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m120_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m121_ns_1_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__79321\,
            in1 => \N__79834\,
            in2 => \N__64364\,
            in3 => \N__64361\,
            lcout => \PROM.ROMDATA.m121_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m138_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011110001"
        )
    port map (
            in0 => \N__78334\,
            in1 => \N__77692\,
            in2 => \N__75909\,
            in3 => \N__77067\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m147_am_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64769\,
            in2 => \N__64763\,
            in3 => \N__76350\,
            lcout => \PROM.ROMDATA.m147_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m80_bm_1_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100111"
        )
    port map (
            in0 => \N__78333\,
            in1 => \N__77690\,
            in2 => \N__76498\,
            in3 => \N__77065\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m80_bm_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m80_bm_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010100010"
        )
    port map (
            in0 => \N__77691\,
            in1 => \N__76349\,
            in2 => \N__64760\,
            in3 => \N__75711\,
            lcout => \PROM.ROMDATA.m80_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m4_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111001010"
        )
    port map (
            in0 => \N__64740\,
            in1 => \N__64710\,
            in2 => \N__64662\,
            in3 => \N__77066\,
            lcout => \PROM.ROMDATA.m4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m347_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__77069\,
            in1 => \N__78336\,
            in2 => \_gnd_net_\,
            in3 => \N__77744\,
            lcout => \PROM.ROMDATA.m347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m292_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__73552\,
            in1 => \N__73809\,
            in2 => \N__73730\,
            in3 => \N__77070\,
            lcout => \PROM.ROMDATA.m292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m112_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__77068\,
            in1 => \N__78335\,
            in2 => \_gnd_net_\,
            in3 => \N__77743\,
            lcout => \PROM.ROMDATA.m112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m137_bm_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__76263\,
            in1 => \N__64544\,
            in2 => \_gnd_net_\,
            in3 => \N__64538\,
            lcout => \PROM.ROMDATA.m137_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m83_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__78793\,
            in1 => \N__77888\,
            in2 => \_gnd_net_\,
            in3 => \N__77238\,
            lcout => \PROM.ROMDATA.m83\,
            ltout => \PROM.ROMDATA.m83_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m161_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__76261\,
            in1 => \N__75636\,
            in2 => \N__64976\,
            in3 => \N__64940\,
            lcout => \PROM.ROMDATA.m161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m15_LC_23_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000010001"
        )
    port map (
            in0 => \N__78792\,
            in1 => \N__77887\,
            in2 => \_gnd_net_\,
            in3 => \N__77237\,
            lcout => \PROM.ROMDATA.m15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m128_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010101101"
        )
    port map (
            in0 => \N__77239\,
            in1 => \N__75637\,
            in2 => \N__78020\,
            in3 => \N__78794\,
            lcout => \PROM.ROMDATA.m128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m171_ns_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__64778\,
            in1 => \_gnd_net_\,
            in2 => \N__79890\,
            in3 => \N__65102\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m171_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m172_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__79454\,
            in1 => \_gnd_net_\,
            in2 => \N__64913\,
            in3 => \N__64910\,
            lcout => \PROM.ROMDATA.m172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m171_bm_LC_23_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__75638\,
            in1 => \N__76262\,
            in2 => \N__64876\,
            in3 => \N__64789\,
            lcout => \PROM.ROMDATA.m171_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m383_LC_23_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__77886\,
            in1 => \N__77236\,
            in2 => \N__75900\,
            in3 => \N__78506\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m427_am_LC_23_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__76448\,
            in1 => \N__74406\,
            in2 => \N__64772\,
            in3 => \N__75684\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m427_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m427_ns_LC_23_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65249\,
            in2 => \N__65240\,
            in3 => \N__79857\,
            lcout => \PROM.ROMDATA.m427_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m494_ns_1_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__76447\,
            in1 => \N__65213\,
            in2 => \N__65201\,
            in3 => \N__75680\,
            lcout => \PROM.ROMDATA.m494_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m88_LC_23_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100111001"
        )
    port map (
            in0 => \N__77884\,
            in1 => \N__77234\,
            in2 => \N__75899\,
            in3 => \N__78505\,
            lcout => \PROM.ROMDATA.m88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m181_LC_23_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__77235\,
            in1 => \N__78542\,
            in2 => \_gnd_net_\,
            in3 => \N__77885\,
            lcout => \PROM.ROMDATA.m181\,
            ltout => \PROM.ROMDATA.m181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m514_ns_LC_23_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__74489\,
            in1 => \N__65171\,
            in2 => \N__65153\,
            in3 => \N__79487\,
            lcout => \PROM.ROMDATA.m514_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m171_am_LC_23_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__76446\,
            in1 => \N__65114\,
            in2 => \_gnd_net_\,
            in3 => \N__65108\,
            lcout => \PROM.ROMDATA.m171_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_12_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67756\,
            in1 => \N__67686\,
            in2 => \_gnd_net_\,
            in3 => \N__67621\,
            lcout => \ALU.dZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73177\,
            ce => \N__70239\,
            sr => \_gnd_net_\
        );

    \ALU.d_13_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67451\,
            in1 => \N__67508\,
            in2 => \_gnd_net_\,
            in3 => \N__67389\,
            lcout => \ALU.dZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73177\,
            ce => \N__70239\,
            sr => \_gnd_net_\
        );

    \ALU.d_14_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__68144\,
            in1 => \N__68077\,
            in2 => \_gnd_net_\,
            in3 => \N__68012\,
            lcout => \ALU.dZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73177\,
            ce => \N__70239\,
            sr => \_gnd_net_\
        );

    \ALU.c_12_LC_24_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__67753\,
            in1 => \N__67685\,
            in2 => \_gnd_net_\,
            in3 => \N__67610\,
            lcout => \ALU.cZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73188\,
            ce => \N__71553\,
            sr => \_gnd_net_\
        );

    \ALU.c_13_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__67516\,
            in1 => \N__67459\,
            in2 => \_gnd_net_\,
            in3 => \N__67391\,
            lcout => \ALU.cZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73188\,
            ce => \N__71553\,
            sr => \_gnd_net_\
        );

    \ALU.c_14_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__68136\,
            in1 => \N__68076\,
            in2 => \_gnd_net_\,
            in3 => \N__68003\,
            lcout => \ALU.cZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73188\,
            ce => \N__71553\,
            sr => \_gnd_net_\
        );

    \ALU.addsub_cry_8_c_RNI6UUIV5_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111010"
        )
    port map (
            in0 => \N__67164\,
            in1 => \N__68150\,
            in2 => \N__66897\,
            in3 => \N__66860\,
            lcout => \ALU.a_15_d_ns_sx_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMGKJC1_0_2_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__66315\,
            in1 => \N__66085\,
            in2 => \N__65585\,
            in3 => \N__66761\,
            lcout => \ALU.d_RNIMGKJC1_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNIMGKJC1_2_LC_24_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__66762\,
            in1 => \N__66316\,
            in2 => \N__66089\,
            in3 => \N__65584\,
            lcout => OPEN,
            ltout => \ALU.d_RNIMGKJC1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNI0TK6H3_2_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65285\,
            in2 => \N__65279\,
            in3 => \N__65272\,
            lcout => OPEN,
            ltout => \ALU.N_859_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.d_RNISGV438_2_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__69188\,
            in1 => \N__68521\,
            in2 => \N__69176\,
            in3 => \N__68897\,
            lcout => OPEN,
            ltout => \ALU.rshift_15_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI0UFMPC_15_LC_24_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__68522\,
            in1 => \N__68567\,
            in2 => \N__69173\,
            in3 => \N__68167\,
            lcout => OPEN,
            ltout => \ALU.rshift_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNI98D92D_15_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__69150\,
            in1 => \_gnd_net_\,
            in2 => \N__69077\,
            in3 => \N__69057\,
            lcout => \ALU.c_RNI98D92DZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNICBIG85_15_LC_24_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__68896\,
            in1 => \N__68566\,
            in2 => \N__68531\,
            in3 => \N__68166\,
            lcout => \ALU.c_RNICBIG85Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.b_14_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__68140\,
            in1 => \N__68079\,
            in2 => \_gnd_net_\,
            in3 => \N__68011\,
            lcout => \ALU.bZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73209\,
            ce => \N__67921\,
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_8_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__70268\,
            in1 => \N__70891\,
            in2 => \N__69338\,
            in3 => \N__69284\,
            lcout => \ALU.un1_a41_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_4_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__70889\,
            in1 => \N__69333\,
            in2 => \N__70942\,
            in3 => \N__70259\,
            lcout => \ALU.un1_a41_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_operation_10_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__67820\,
            in1 => \N__69966\,
            in2 => \N__67808\,
            in3 => \N__69799\,
            lcout => \ALU.un1_operation_10_0\,
            ltout => \ALU.un1_operation_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_7_2_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100010001"
        )
    port map (
            in0 => \N__70931\,
            in1 => \N__71515\,
            in2 => \N__67787\,
            in3 => \N__71469\,
            lcout => \ALU.un1_a41_7_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_operation_13_2_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__69967\,
            in1 => \N__69798\,
            in2 => \N__69716\,
            in3 => \N__70157\,
            lcout => \ALU.un1_operation_13Z0Z_2\,
            ltout => \ALU.un1_operation_13Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_4_2_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000001010"
        )
    port map (
            in0 => \N__69283\,
            in1 => \N__71491\,
            in2 => \N__70262\,
            in3 => \N__71468\,
            lcout => \ALU.un1_a41_4_0_2\,
            ltout => \ALU.un1_a41_4_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_6_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__69337\,
            in1 => \N__70935\,
            in2 => \N__70253\,
            in3 => \N__70890\,
            lcout => \ALU.un1_a41_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_operation_7_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__70158\,
            in1 => \N__69968\,
            in2 => \N__69803\,
            in3 => \N__69697\,
            lcout => \ALU.un1_operationZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_2_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__71007\,
            in1 => \N__69332\,
            in2 => \N__70844\,
            in3 => \N__69282\,
            lcout => \ALU.un1_a41_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m160_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__78842\,
            in1 => \N__78066\,
            in2 => \N__76003\,
            in3 => \N__77317\,
            lcout => \PROM.ROMDATA.m160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_3_1_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69331\,
            in2 => \_gnd_net_\,
            in3 => \N__69281\,
            lcout => \ALU.un1_a41_3_0_1\,
            ltout => \ALU.un1_a41_3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_5_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__70940\,
            in1 => \N__70883\,
            in2 => \N__69248\,
            in3 => \N__71008\,
            lcout => \ALU.un1_a41_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_7_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__71009\,
            in1 => \N__70941\,
            in2 => \N__70892\,
            in3 => \N__71019\,
            lcout => \ALU.un1_a41_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_operation_13_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__71519\,
            in1 => \N__71490\,
            in2 => \_gnd_net_\,
            in3 => \N__71470\,
            lcout => \ALU.un1_operation_13_0\,
            ltout => \ALU.un1_operation_13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_9_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__70887\,
            in1 => \N__70936\,
            in2 => \N__71219\,
            in3 => \N__71020\,
            lcout => \ALU.un1_a41_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_3_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__71021\,
            in1 => \N__70888\,
            in2 => \N__70943\,
            in3 => \N__71006\,
            lcout => \ALU.un1_a41_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.un1_a41_2_1_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__70914\,
            in2 => \_gnd_net_\,
            in3 => \N__70865\,
            lcout => \ALU.un1_a41_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.ramAddReg_6_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__70835\,
            in1 => \N__70799\,
            in2 => \N__70613\,
            in3 => \N__70556\,
            lcout => \A6_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVCONTROL.ramAddReg_6C_net\,
            ce => \N__70329\,
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m281_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__78714\,
            in1 => \N__77907\,
            in2 => \_gnd_net_\,
            in3 => \N__77257\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m480_bm_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76559\,
            in2 => \N__70271\,
            in3 => \N__75808\,
            lcout => \PROM.ROMDATA.m480_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m60_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__78713\,
            in1 => \N__77906\,
            in2 => \_gnd_net_\,
            in3 => \N__77256\,
            lcout => \PROM.ROMDATA.m60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.programCounter_ret_1_7_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__73355\,
            lcout => \CONTROL.programCounter_1_reto_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__73258\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m480_am_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100000001000"
        )
    port map (
            in0 => \N__75809\,
            in1 => \N__72827\,
            in2 => \N__76616\,
            in3 => \N__74488\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m480_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m480_ns_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__72815\,
            in2 => \N__72809\,
            in3 => \N__79898\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m480_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m485_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111000"
        )
    port map (
            in0 => \N__72806\,
            in1 => \N__72696\,
            in2 => \N__72383\,
            in3 => \N__79502\,
            lcout => \PROM_ROMDATA_dintern_25ro\,
            ltout => \PROM_ROMDATA_dintern_25ro_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONTROL.romAddReg_7_9_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__72352\,
            in1 => \N__72318\,
            in2 => \N__71879\,
            in3 => \N__71875\,
            lcout => \CONTROL_romAddReg_7_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m262_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000100"
        )
    port map (
            in0 => \N__77247\,
            in1 => \N__75891\,
            in2 => \N__78839\,
            in3 => \N__77908\,
            lcout => \PROM.ROMDATA.m262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m447_ns_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__71615\,
            in1 => \N__71603\,
            in2 => \N__71588\,
            in3 => \N__79866\,
            lcout => \PROM.ROMDATA.m447_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m488_ns_1_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010010"
        )
    port map (
            in0 => \N__75892\,
            in1 => \N__78718\,
            in2 => \N__76601\,
            in3 => \N__77248\,
            lcout => \PROM.ROMDATA.m488_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m503_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__78719\,
            in1 => \N__74071\,
            in2 => \N__75986\,
            in3 => \N__73505\,
            lcout => \PROM.ROMDATA.N_570_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m493_am_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__73728\,
            in1 => \N__73565\,
            in2 => \N__73911\,
            in3 => \N__73812\,
            lcout => \PROM.ROMDATA.m493_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m493_bm_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__73813\,
            in1 => \N__73729\,
            in2 => \N__73573\,
            in3 => \N__73504\,
            lcout => \PROM.ROMDATA.m493_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m361_ns_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__74192\,
            in1 => \N__73454\,
            in2 => \_gnd_net_\,
            in3 => \N__76522\,
            lcout => \PROM.ROMDATA.m361_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m211_ns_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011010110100"
        )
    port map (
            in0 => \N__78473\,
            in1 => \N__77961\,
            in2 => \N__73448\,
            in3 => \N__77241\,
            lcout => \PROM.ROMDATA.m211_ns\,
            ltout => \PROM.ROMDATA.m211_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m221cf0_1_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__79323\,
            in2 => \N__73436\,
            in3 => \N__79831\,
            lcout => \PROM.ROMDATA.m221cf0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m221cf1_1_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011111"
        )
    port map (
            in0 => \N__79832\,
            in1 => \_gnd_net_\,
            in2 => \N__79414\,
            in3 => \N__73418\,
            lcout => \PROM.ROMDATA.m221cf1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m369_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111100011"
        )
    port map (
            in0 => \N__77242\,
            in1 => \N__75810\,
            in2 => \N__78042\,
            in3 => \N__78474\,
            lcout => \PROM.ROMDATA.m369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m373_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001001000101"
        )
    port map (
            in0 => \N__78475\,
            in1 => \N__77965\,
            in2 => \N__75959\,
            in3 => \N__77243\,
            lcout => \PROM.ROMDATA.m373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m303_ns_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__74270\,
            in1 => \N__79327\,
            in2 => \N__74360\,
            in3 => \N__74093\,
            lcout => \PROM.ROMDATA.m303_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m424_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__79833\,
            in1 => \N__74239\,
            in2 => \_gnd_net_\,
            in3 => \N__74225\,
            lcout => \PROM.ROMDATA.m424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m361_bm_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010110111111"
        )
    port map (
            in0 => \N__77172\,
            in1 => \N__75718\,
            in2 => \N__78035\,
            in3 => \N__78858\,
            lcout => \PROM.ROMDATA.m361_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m137_am_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__74186\,
            in1 => \N__76372\,
            in2 => \_gnd_net_\,
            in3 => \N__74171\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m137_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m148_ns_1_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__79452\,
            in1 => \N__79858\,
            in2 => \N__74165\,
            in3 => \N__74162\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m148_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m148_ns_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__74156\,
            in1 => \N__74150\,
            in2 => \N__74141\,
            in3 => \N__79453\,
            lcout => \PROM.ROMDATA.m148_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m301_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__76374\,
            in1 => \N__74125\,
            in2 => \N__74108\,
            in3 => \N__75720\,
            lcout => \PROM.ROMDATA.m301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m349_am_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111101110101"
        )
    port map (
            in0 => \N__78857\,
            in1 => \N__77933\,
            in2 => \N__75910\,
            in3 => \N__77171\,
            lcout => \PROM.ROMDATA.m349_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m357_am_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111011011"
        )
    port map (
            in0 => \N__77173\,
            in1 => \N__75719\,
            in2 => \N__78036\,
            in3 => \N__78859\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m357_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m357_ns_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74501\,
            in2 => \N__74495\,
            in3 => \N__76373\,
            lcout => \PROM.ROMDATA.m357_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m290_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__76533\,
            in1 => \N__74490\,
            in2 => \N__74411\,
            in3 => \N__75725\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m303_ns_1_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__74378\,
            in1 => \N__79457\,
            in2 => \N__74363\,
            in3 => \N__79860\,
            lcout => \PROM.ROMDATA.m303_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m363_ns_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__79456\,
            in1 => \N__74348\,
            in2 => \N__74339\,
            in3 => \N__74291\,
            lcout => \PROM.ROMDATA.m363_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m353_am_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111011101"
        )
    port map (
            in0 => \N__78720\,
            in1 => \N__77892\,
            in2 => \N__75911\,
            in3 => \N__77240\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m353_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m353_ns_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__76532\,
            in1 => \_gnd_net_\,
            in2 => \N__74312\,
            in3 => \N__74309\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m353_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m363_ns_1_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__74936\,
            in1 => \N__79455\,
            in2 => \N__74294\,
            in3 => \N__79859\,
            lcout => \PROM.ROMDATA.m363_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m349_bm_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__74972\,
            in1 => \N__74962\,
            in2 => \_gnd_net_\,
            in3 => \N__75721\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m349_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m349_ns_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74945\,
            in2 => \N__74939\,
            in3 => \N__76531\,
            lcout => \PROM.ROMDATA.m349_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m331_bm_LC_26_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100001000"
        )
    port map (
            in0 => \N__78843\,
            in1 => \N__78011\,
            in2 => \N__76010\,
            in3 => \N__77309\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m331_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m331_ns_LC_26_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74507\,
            in2 => \N__74930\,
            in3 => \N__76617\,
            lcout => \PROM.ROMDATA.m331_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m323_am_LC_26_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000111000"
        )
    port map (
            in0 => \N__78841\,
            in1 => \N__78069\,
            in2 => \N__76016\,
            in3 => \N__77310\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m323_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m323_ns_LC_26_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__74927\,
            in2 => \N__74915\,
            in3 => \N__76618\,
            lcout => \PROM.ROMDATA.m323_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU.c_RNIFS1RP_15_LC_26_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110111011"
        )
    port map (
            in0 => \N__74855\,
            in1 => \N__74618\,
            in2 => \_gnd_net_\,
            in3 => \N__74596\,
            lcout => \ALU.N_586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m331_am_LC_26_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101000"
        )
    port map (
            in0 => \N__76011\,
            in1 => \N__78840\,
            in2 => \N__79049\,
            in3 => \N__78068\,
            lcout => \PROM.ROMDATA.m331_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m341_ns_1_LC_26_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100111110"
        )
    port map (
            in0 => \N__78637\,
            in1 => \N__78067\,
            in2 => \N__76008\,
            in3 => \N__77318\,
            lcout => \PROM.ROMDATA.m341_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m343_ns_1_LC_26_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__79907\,
            in1 => \N__79415\,
            in2 => \N__78872\,
            in3 => \N__79883\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m343_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m343_ns_LC_26_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__79416\,
            in1 => \N__74978\,
            in2 => \N__79067\,
            in3 => \N__76661\,
            lcout => \PROM.ROMDATA.m343_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m334_ns_1_LC_26_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__76569\,
            in1 => \N__79044\,
            in2 => \_gnd_net_\,
            in3 => \N__78998\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m334_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m334_ns_LC_26_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100000000"
        )
    port map (
            in0 => \N__78061\,
            in1 => \N__78887\,
            in2 => \N__78875\,
            in3 => \N__78778\,
            lcout => \PROM.ROMDATA.i3_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m338_am_LC_26_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011110001100"
        )
    port map (
            in0 => \N__78777\,
            in1 => \N__78062\,
            in2 => \N__76009\,
            in3 => \N__77311\,
            lcout => OPEN,
            ltout => \PROM.ROMDATA.m338_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m338_ns_LC_26_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__76679\,
            in2 => \N__76664\,
            in3 => \N__76571\,
            lcout => \PROM.ROMDATA.m338_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PROM.ROMDATA.dintern_31_0__m341_ns_LC_26_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011010001"
        )
    port map (
            in0 => \N__76655\,
            in1 => \N__76570\,
            in2 => \N__76028\,
            in3 => \N__75983\,
            lcout => \PROM.ROMDATA.m341_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
