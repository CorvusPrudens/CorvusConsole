// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Aug 18 2020 14:56:44

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    TX,
    GPIO11,
    CLK,
    RX,
    GPIO9,
    GPIO3);

    output TX;
    output GPIO11;
    input CLK;
    input RX;
    output GPIO9;
    output GPIO3;

    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49515;
    wire N__49514;
    wire N__49513;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49469;
    wire N__49468;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49460;
    wire N__49457;
    wire N__49454;
    wire N__49451;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49443;
    wire N__49442;
    wire N__49441;
    wire N__49438;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49426;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49410;
    wire N__49407;
    wire N__49402;
    wire N__49397;
    wire N__49388;
    wire N__49387;
    wire N__49384;
    wire N__49383;
    wire N__49382;
    wire N__49379;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49368;
    wire N__49365;
    wire N__49362;
    wire N__49361;
    wire N__49360;
    wire N__49355;
    wire N__49352;
    wire N__49349;
    wire N__49346;
    wire N__49343;
    wire N__49340;
    wire N__49337;
    wire N__49334;
    wire N__49331;
    wire N__49328;
    wire N__49319;
    wire N__49310;
    wire N__49307;
    wire N__49304;
    wire N__49303;
    wire N__49300;
    wire N__49297;
    wire N__49294;
    wire N__49289;
    wire N__49288;
    wire N__49287;
    wire N__49286;
    wire N__49285;
    wire N__49282;
    wire N__49281;
    wire N__49278;
    wire N__49275;
    wire N__49272;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49262;
    wire N__49259;
    wire N__49248;
    wire N__49245;
    wire N__49244;
    wire N__49241;
    wire N__49236;
    wire N__49233;
    wire N__49230;
    wire N__49225;
    wire N__49220;
    wire N__49219;
    wire N__49218;
    wire N__49217;
    wire N__49214;
    wire N__49213;
    wire N__49212;
    wire N__49211;
    wire N__49208;
    wire N__49205;
    wire N__49204;
    wire N__49201;
    wire N__49198;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49184;
    wire N__49181;
    wire N__49178;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49162;
    wire N__49151;
    wire N__49148;
    wire N__49145;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49124;
    wire N__49123;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49112;
    wire N__49105;
    wire N__49102;
    wire N__49101;
    wire N__49098;
    wire N__49095;
    wire N__49094;
    wire N__49091;
    wire N__49090;
    wire N__49089;
    wire N__49086;
    wire N__49083;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49071;
    wire N__49068;
    wire N__49063;
    wire N__49056;
    wire N__49049;
    wire N__49048;
    wire N__49047;
    wire N__49046;
    wire N__49045;
    wire N__49044;
    wire N__49043;
    wire N__49040;
    wire N__49037;
    wire N__49034;
    wire N__49031;
    wire N__49028;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49013;
    wire N__49010;
    wire N__49007;
    wire N__49004;
    wire N__48999;
    wire N__48996;
    wire N__48991;
    wire N__48986;
    wire N__48983;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48965;
    wire N__48964;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48950;
    wire N__48947;
    wire N__48944;
    wire N__48943;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48933;
    wire N__48932;
    wire N__48931;
    wire N__48924;
    wire N__48921;
    wire N__48918;
    wire N__48917;
    wire N__48916;
    wire N__48909;
    wire N__48906;
    wire N__48903;
    wire N__48896;
    wire N__48893;
    wire N__48892;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48881;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48868;
    wire N__48867;
    wire N__48864;
    wire N__48863;
    wire N__48860;
    wire N__48857;
    wire N__48856;
    wire N__48851;
    wire N__48848;
    wire N__48845;
    wire N__48842;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48824;
    wire N__48815;
    wire N__48812;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48799;
    wire N__48796;
    wire N__48791;
    wire N__48790;
    wire N__48789;
    wire N__48788;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48777;
    wire N__48774;
    wire N__48771;
    wire N__48770;
    wire N__48765;
    wire N__48762;
    wire N__48759;
    wire N__48756;
    wire N__48753;
    wire N__48750;
    wire N__48749;
    wire N__48742;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48726;
    wire N__48723;
    wire N__48716;
    wire N__48715;
    wire N__48714;
    wire N__48713;
    wire N__48710;
    wire N__48707;
    wire N__48704;
    wire N__48701;
    wire N__48700;
    wire N__48697;
    wire N__48696;
    wire N__48695;
    wire N__48688;
    wire N__48685;
    wire N__48684;
    wire N__48681;
    wire N__48678;
    wire N__48675;
    wire N__48670;
    wire N__48667;
    wire N__48656;
    wire N__48655;
    wire N__48650;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48640;
    wire N__48639;
    wire N__48638;
    wire N__48637;
    wire N__48636;
    wire N__48635;
    wire N__48634;
    wire N__48633;
    wire N__48632;
    wire N__48631;
    wire N__48630;
    wire N__48629;
    wire N__48628;
    wire N__48627;
    wire N__48626;
    wire N__48625;
    wire N__48624;
    wire N__48623;
    wire N__48622;
    wire N__48621;
    wire N__48620;
    wire N__48619;
    wire N__48618;
    wire N__48617;
    wire N__48616;
    wire N__48615;
    wire N__48606;
    wire N__48599;
    wire N__48598;
    wire N__48597;
    wire N__48596;
    wire N__48595;
    wire N__48594;
    wire N__48593;
    wire N__48592;
    wire N__48591;
    wire N__48590;
    wire N__48589;
    wire N__48588;
    wire N__48587;
    wire N__48586;
    wire N__48585;
    wire N__48584;
    wire N__48583;
    wire N__48582;
    wire N__48581;
    wire N__48580;
    wire N__48579;
    wire N__48578;
    wire N__48577;
    wire N__48576;
    wire N__48575;
    wire N__48574;
    wire N__48573;
    wire N__48572;
    wire N__48571;
    wire N__48570;
    wire N__48569;
    wire N__48568;
    wire N__48567;
    wire N__48566;
    wire N__48565;
    wire N__48564;
    wire N__48563;
    wire N__48562;
    wire N__48561;
    wire N__48560;
    wire N__48557;
    wire N__48556;
    wire N__48555;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48535;
    wire N__48526;
    wire N__48517;
    wire N__48510;
    wire N__48509;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48497;
    wire N__48496;
    wire N__48495;
    wire N__48494;
    wire N__48493;
    wire N__48492;
    wire N__48491;
    wire N__48490;
    wire N__48489;
    wire N__48488;
    wire N__48487;
    wire N__48486;
    wire N__48485;
    wire N__48484;
    wire N__48483;
    wire N__48472;
    wire N__48469;
    wire N__48464;
    wire N__48461;
    wire N__48454;
    wire N__48447;
    wire N__48444;
    wire N__48437;
    wire N__48436;
    wire N__48435;
    wire N__48434;
    wire N__48433;
    wire N__48432;
    wire N__48431;
    wire N__48430;
    wire N__48427;
    wire N__48426;
    wire N__48425;
    wire N__48424;
    wire N__48423;
    wire N__48422;
    wire N__48421;
    wire N__48420;
    wire N__48419;
    wire N__48416;
    wire N__48413;
    wire N__48412;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48406;
    wire N__48401;
    wire N__48396;
    wire N__48389;
    wire N__48384;
    wire N__48375;
    wire N__48366;
    wire N__48363;
    wire N__48354;
    wire N__48349;
    wire N__48348;
    wire N__48347;
    wire N__48346;
    wire N__48345;
    wire N__48344;
    wire N__48341;
    wire N__48340;
    wire N__48339;
    wire N__48334;
    wire N__48331;
    wire N__48330;
    wire N__48329;
    wire N__48328;
    wire N__48317;
    wire N__48310;
    wire N__48301;
    wire N__48294;
    wire N__48291;
    wire N__48284;
    wire N__48275;
    wire N__48274;
    wire N__48273;
    wire N__48272;
    wire N__48271;
    wire N__48270;
    wire N__48269;
    wire N__48268;
    wire N__48267;
    wire N__48266;
    wire N__48265;
    wire N__48262;
    wire N__48261;
    wire N__48258;
    wire N__48255;
    wire N__48252;
    wire N__48251;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48227;
    wire N__48222;
    wire N__48215;
    wire N__48208;
    wire N__48203;
    wire N__48186;
    wire N__48183;
    wire N__48174;
    wire N__48171;
    wire N__48166;
    wire N__48161;
    wire N__48156;
    wire N__48153;
    wire N__48146;
    wire N__48137;
    wire N__48132;
    wire N__48127;
    wire N__48122;
    wire N__48113;
    wire N__48110;
    wire N__48109;
    wire N__48106;
    wire N__48105;
    wire N__48100;
    wire N__48097;
    wire N__48096;
    wire N__48095;
    wire N__48094;
    wire N__48093;
    wire N__48092;
    wire N__48089;
    wire N__48078;
    wire N__48077;
    wire N__48076;
    wire N__48075;
    wire N__48074;
    wire N__48065;
    wire N__48060;
    wire N__48055;
    wire N__48054;
    wire N__48049;
    wire N__48034;
    wire N__48031;
    wire N__48030;
    wire N__48029;
    wire N__48026;
    wire N__48023;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48007;
    wire N__48002;
    wire N__47997;
    wire N__47990;
    wire N__47987;
    wire N__47984;
    wire N__47979;
    wire N__47976;
    wire N__47971;
    wire N__47968;
    wire N__47963;
    wire N__47958;
    wire N__47953;
    wire N__47950;
    wire N__47941;
    wire N__47934;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47918;
    wire N__47913;
    wire N__47908;
    wire N__47905;
    wire N__47894;
    wire N__47893;
    wire N__47892;
    wire N__47889;
    wire N__47888;
    wire N__47887;
    wire N__47886;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47871;
    wire N__47868;
    wire N__47865;
    wire N__47864;
    wire N__47861;
    wire N__47858;
    wire N__47853;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47836;
    wire N__47833;
    wire N__47828;
    wire N__47827;
    wire N__47818;
    wire N__47815;
    wire N__47810;
    wire N__47809;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47798;
    wire N__47795;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47785;
    wire N__47782;
    wire N__47779;
    wire N__47778;
    wire N__47777;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47720;
    wire N__47719;
    wire N__47716;
    wire N__47713;
    wire N__47710;
    wire N__47707;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47692;
    wire N__47691;
    wire N__47690;
    wire N__47689;
    wire N__47688;
    wire N__47687;
    wire N__47686;
    wire N__47685;
    wire N__47684;
    wire N__47683;
    wire N__47682;
    wire N__47681;
    wire N__47680;
    wire N__47679;
    wire N__47678;
    wire N__47677;
    wire N__47676;
    wire N__47675;
    wire N__47674;
    wire N__47673;
    wire N__47672;
    wire N__47671;
    wire N__47670;
    wire N__47669;
    wire N__47668;
    wire N__47667;
    wire N__47666;
    wire N__47665;
    wire N__47664;
    wire N__47663;
    wire N__47662;
    wire N__47661;
    wire N__47660;
    wire N__47659;
    wire N__47658;
    wire N__47657;
    wire N__47656;
    wire N__47655;
    wire N__47654;
    wire N__47653;
    wire N__47652;
    wire N__47651;
    wire N__47650;
    wire N__47649;
    wire N__47648;
    wire N__47647;
    wire N__47646;
    wire N__47645;
    wire N__47644;
    wire N__47643;
    wire N__47642;
    wire N__47641;
    wire N__47640;
    wire N__47639;
    wire N__47638;
    wire N__47637;
    wire N__47636;
    wire N__47635;
    wire N__47634;
    wire N__47633;
    wire N__47632;
    wire N__47631;
    wire N__47630;
    wire N__47629;
    wire N__47628;
    wire N__47627;
    wire N__47626;
    wire N__47625;
    wire N__47624;
    wire N__47623;
    wire N__47622;
    wire N__47621;
    wire N__47620;
    wire N__47619;
    wire N__47618;
    wire N__47617;
    wire N__47616;
    wire N__47615;
    wire N__47614;
    wire N__47613;
    wire N__47612;
    wire N__47611;
    wire N__47610;
    wire N__47609;
    wire N__47608;
    wire N__47607;
    wire N__47606;
    wire N__47605;
    wire N__47604;
    wire N__47603;
    wire N__47602;
    wire N__47601;
    wire N__47600;
    wire N__47599;
    wire N__47408;
    wire N__47405;
    wire N__47402;
    wire N__47401;
    wire N__47398;
    wire N__47397;
    wire N__47394;
    wire N__47393;
    wire N__47390;
    wire N__47387;
    wire N__47384;
    wire N__47381;
    wire N__47378;
    wire N__47375;
    wire N__47372;
    wire N__47369;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47348;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47324;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47315;
    wire N__47314;
    wire N__47311;
    wire N__47310;
    wire N__47309;
    wire N__47308;
    wire N__47305;
    wire N__47304;
    wire N__47303;
    wire N__47300;
    wire N__47297;
    wire N__47294;
    wire N__47293;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47279;
    wire N__47278;
    wire N__47277;
    wire N__47274;
    wire N__47269;
    wire N__47264;
    wire N__47261;
    wire N__47260;
    wire N__47259;
    wire N__47256;
    wire N__47253;
    wire N__47246;
    wire N__47243;
    wire N__47238;
    wire N__47235;
    wire N__47234;
    wire N__47233;
    wire N__47232;
    wire N__47231;
    wire N__47230;
    wire N__47229;
    wire N__47224;
    wire N__47221;
    wire N__47220;
    wire N__47217;
    wire N__47212;
    wire N__47211;
    wire N__47210;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47194;
    wire N__47185;
    wire N__47180;
    wire N__47179;
    wire N__47178;
    wire N__47173;
    wire N__47170;
    wire N__47165;
    wire N__47160;
    wire N__47157;
    wire N__47154;
    wire N__47151;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47125;
    wire N__47116;
    wire N__47105;
    wire N__47102;
    wire N__47101;
    wire N__47100;
    wire N__47099;
    wire N__47098;
    wire N__47097;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47089;
    wire N__47088;
    wire N__47087;
    wire N__47084;
    wire N__47077;
    wire N__47074;
    wire N__47071;
    wire N__47068;
    wire N__47067;
    wire N__47064;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47051;
    wire N__47050;
    wire N__47049;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47032;
    wire N__47025;
    wire N__47022;
    wire N__47017;
    wire N__47014;
    wire N__47005;
    wire N__47002;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46979;
    wire N__46976;
    wire N__46975;
    wire N__46974;
    wire N__46973;
    wire N__46970;
    wire N__46967;
    wire N__46966;
    wire N__46965;
    wire N__46964;
    wire N__46963;
    wire N__46962;
    wire N__46961;
    wire N__46960;
    wire N__46957;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46946;
    wire N__46945;
    wire N__46944;
    wire N__46943;
    wire N__46942;
    wire N__46937;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46925;
    wire N__46922;
    wire N__46919;
    wire N__46918;
    wire N__46913;
    wire N__46912;
    wire N__46911;
    wire N__46908;
    wire N__46907;
    wire N__46904;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46890;
    wire N__46887;
    wire N__46884;
    wire N__46877;
    wire N__46876;
    wire N__46873;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46847;
    wire N__46840;
    wire N__46839;
    wire N__46838;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46820;
    wire N__46817;
    wire N__46814;
    wire N__46813;
    wire N__46808;
    wire N__46799;
    wire N__46794;
    wire N__46791;
    wire N__46788;
    wire N__46783;
    wire N__46780;
    wire N__46773;
    wire N__46770;
    wire N__46763;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46739;
    wire N__46736;
    wire N__46735;
    wire N__46734;
    wire N__46733;
    wire N__46730;
    wire N__46729;
    wire N__46728;
    wire N__46727;
    wire N__46724;
    wire N__46721;
    wire N__46720;
    wire N__46717;
    wire N__46716;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46700;
    wire N__46697;
    wire N__46694;
    wire N__46693;
    wire N__46690;
    wire N__46687;
    wire N__46686;
    wire N__46683;
    wire N__46682;
    wire N__46681;
    wire N__46676;
    wire N__46673;
    wire N__46672;
    wire N__46671;
    wire N__46670;
    wire N__46669;
    wire N__46666;
    wire N__46659;
    wire N__46658;
    wire N__46657;
    wire N__46654;
    wire N__46649;
    wire N__46648;
    wire N__46645;
    wire N__46642;
    wire N__46639;
    wire N__46638;
    wire N__46635;
    wire N__46630;
    wire N__46627;
    wire N__46626;
    wire N__46623;
    wire N__46622;
    wire N__46617;
    wire N__46616;
    wire N__46615;
    wire N__46612;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46559;
    wire N__46556;
    wire N__46551;
    wire N__46546;
    wire N__46543;
    wire N__46538;
    wire N__46535;
    wire N__46530;
    wire N__46525;
    wire N__46522;
    wire N__46517;
    wire N__46512;
    wire N__46509;
    wire N__46504;
    wire N__46495;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46475;
    wire N__46474;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46463;
    wire N__46462;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46449;
    wire N__46448;
    wire N__46445;
    wire N__46444;
    wire N__46443;
    wire N__46438;
    wire N__46433;
    wire N__46430;
    wire N__46427;
    wire N__46424;
    wire N__46421;
    wire N__46418;
    wire N__46413;
    wire N__46400;
    wire N__46397;
    wire N__46394;
    wire N__46393;
    wire N__46392;
    wire N__46391;
    wire N__46388;
    wire N__46385;
    wire N__46384;
    wire N__46383;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46367;
    wire N__46364;
    wire N__46363;
    wire N__46362;
    wire N__46359;
    wire N__46354;
    wire N__46353;
    wire N__46352;
    wire N__46349;
    wire N__46346;
    wire N__46343;
    wire N__46340;
    wire N__46335;
    wire N__46332;
    wire N__46331;
    wire N__46330;
    wire N__46327;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46317;
    wire N__46312;
    wire N__46311;
    wire N__46310;
    wire N__46305;
    wire N__46302;
    wire N__46299;
    wire N__46296;
    wire N__46293;
    wire N__46290;
    wire N__46285;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46266;
    wire N__46259;
    wire N__46256;
    wire N__46253;
    wire N__46250;
    wire N__46245;
    wire N__46240;
    wire N__46229;
    wire N__46226;
    wire N__46223;
    wire N__46220;
    wire N__46217;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46201;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46193;
    wire N__46192;
    wire N__46191;
    wire N__46190;
    wire N__46189;
    wire N__46186;
    wire N__46181;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46165;
    wire N__46164;
    wire N__46163;
    wire N__46162;
    wire N__46161;
    wire N__46160;
    wire N__46159;
    wire N__46158;
    wire N__46157;
    wire N__46156;
    wire N__46155;
    wire N__46154;
    wire N__46153;
    wire N__46152;
    wire N__46151;
    wire N__46150;
    wire N__46149;
    wire N__46148;
    wire N__46147;
    wire N__46144;
    wire N__46141;
    wire N__46138;
    wire N__46123;
    wire N__46122;
    wire N__46119;
    wire N__46118;
    wire N__46117;
    wire N__46114;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46085;
    wire N__46084;
    wire N__46083;
    wire N__46082;
    wire N__46081;
    wire N__46080;
    wire N__46079;
    wire N__46078;
    wire N__46077;
    wire N__46076;
    wire N__46073;
    wire N__46070;
    wire N__46067;
    wire N__46064;
    wire N__46061;
    wire N__46060;
    wire N__46057;
    wire N__46050;
    wire N__46047;
    wire N__46046;
    wire N__46045;
    wire N__46042;
    wire N__46041;
    wire N__46040;
    wire N__46037;
    wire N__46034;
    wire N__46033;
    wire N__46024;
    wire N__46017;
    wire N__46008;
    wire N__46005;
    wire N__46004;
    wire N__46003;
    wire N__46002;
    wire N__46001;
    wire N__46000;
    wire N__45997;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45990;
    wire N__45989;
    wire N__45986;
    wire N__45983;
    wire N__45980;
    wire N__45977;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45967;
    wire N__45962;
    wire N__45953;
    wire N__45950;
    wire N__45947;
    wire N__45940;
    wire N__45937;
    wire N__45934;
    wire N__45931;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45923;
    wire N__45920;
    wire N__45913;
    wire N__45910;
    wire N__45907;
    wire N__45904;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45893;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45877;
    wire N__45874;
    wire N__45873;
    wire N__45866;
    wire N__45857;
    wire N__45854;
    wire N__45843;
    wire N__45842;
    wire N__45837;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45808;
    wire N__45805;
    wire N__45798;
    wire N__45795;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45769;
    wire N__45766;
    wire N__45763;
    wire N__45760;
    wire N__45751;
    wire N__45748;
    wire N__45741;
    wire N__45734;
    wire N__45731;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45713;
    wire N__45710;
    wire N__45705;
    wire N__45700;
    wire N__45699;
    wire N__45698;
    wire N__45697;
    wire N__45692;
    wire N__45685;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45656;
    wire N__45653;
    wire N__45638;
    wire N__45635;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45622;
    wire N__45619;
    wire N__45616;
    wire N__45613;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45601;
    wire N__45598;
    wire N__45595;
    wire N__45592;
    wire N__45587;
    wire N__45586;
    wire N__45583;
    wire N__45580;
    wire N__45575;
    wire N__45574;
    wire N__45573;
    wire N__45572;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45538;
    wire N__45535;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45525;
    wire N__45522;
    wire N__45517;
    wire N__45514;
    wire N__45511;
    wire N__45508;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45498;
    wire N__45495;
    wire N__45490;
    wire N__45489;
    wire N__45486;
    wire N__45483;
    wire N__45476;
    wire N__45473;
    wire N__45468;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45447;
    wire N__45444;
    wire N__45439;
    wire N__45436;
    wire N__45431;
    wire N__45428;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45410;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45392;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45374;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45364;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45350;
    wire N__45349;
    wire N__45346;
    wire N__45343;
    wire N__45338;
    wire N__45337;
    wire N__45336;
    wire N__45335;
    wire N__45334;
    wire N__45333;
    wire N__45330;
    wire N__45323;
    wire N__45322;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45314;
    wire N__45313;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45300;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45288;
    wire N__45285;
    wire N__45284;
    wire N__45283;
    wire N__45282;
    wire N__45281;
    wire N__45280;
    wire N__45279;
    wire N__45278;
    wire N__45277;
    wire N__45276;
    wire N__45275;
    wire N__45270;
    wire N__45265;
    wire N__45262;
    wire N__45255;
    wire N__45252;
    wire N__45247;
    wire N__45242;
    wire N__45231;
    wire N__45228;
    wire N__45223;
    wire N__45216;
    wire N__45203;
    wire N__45200;
    wire N__45197;
    wire N__45194;
    wire N__45191;
    wire N__45188;
    wire N__45185;
    wire N__45182;
    wire N__45179;
    wire N__45176;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45158;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45148;
    wire N__45145;
    wire N__45142;
    wire N__45137;
    wire N__45136;
    wire N__45135;
    wire N__45130;
    wire N__45129;
    wire N__45128;
    wire N__45127;
    wire N__45126;
    wire N__45123;
    wire N__45122;
    wire N__45121;
    wire N__45120;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45112;
    wire N__45109;
    wire N__45104;
    wire N__45103;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45081;
    wire N__45080;
    wire N__45079;
    wire N__45078;
    wire N__45077;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45064;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45030;
    wire N__45027;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45009;
    wire N__45004;
    wire N__44987;
    wire N__44984;
    wire N__44981;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44963;
    wire N__44960;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44942;
    wire N__44939;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44927;
    wire N__44924;
    wire N__44921;
    wire N__44918;
    wire N__44915;
    wire N__44912;
    wire N__44909;
    wire N__44908;
    wire N__44907;
    wire N__44904;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44888;
    wire N__44885;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44873;
    wire N__44872;
    wire N__44871;
    wire N__44870;
    wire N__44867;
    wire N__44864;
    wire N__44861;
    wire N__44858;
    wire N__44853;
    wire N__44850;
    wire N__44849;
    wire N__44846;
    wire N__44841;
    wire N__44838;
    wire N__44837;
    wire N__44834;
    wire N__44831;
    wire N__44828;
    wire N__44825;
    wire N__44822;
    wire N__44819;
    wire N__44816;
    wire N__44813;
    wire N__44810;
    wire N__44807;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44792;
    wire N__44789;
    wire N__44780;
    wire N__44777;
    wire N__44774;
    wire N__44771;
    wire N__44770;
    wire N__44769;
    wire N__44768;
    wire N__44763;
    wire N__44760;
    wire N__44759;
    wire N__44758;
    wire N__44757;
    wire N__44756;
    wire N__44755;
    wire N__44754;
    wire N__44753;
    wire N__44750;
    wire N__44749;
    wire N__44748;
    wire N__44745;
    wire N__44744;
    wire N__44741;
    wire N__44726;
    wire N__44723;
    wire N__44720;
    wire N__44719;
    wire N__44718;
    wire N__44717;
    wire N__44714;
    wire N__44711;
    wire N__44708;
    wire N__44701;
    wire N__44698;
    wire N__44693;
    wire N__44688;
    wire N__44675;
    wire N__44672;
    wire N__44669;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44659;
    wire N__44656;
    wire N__44653;
    wire N__44648;
    wire N__44645;
    wire N__44642;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44612;
    wire N__44609;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44540;
    wire N__44539;
    wire N__44538;
    wire N__44537;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44527;
    wire N__44526;
    wire N__44525;
    wire N__44524;
    wire N__44523;
    wire N__44522;
    wire N__44521;
    wire N__44520;
    wire N__44519;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44501;
    wire N__44500;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44492;
    wire N__44491;
    wire N__44488;
    wire N__44487;
    wire N__44484;
    wire N__44481;
    wire N__44480;
    wire N__44479;
    wire N__44476;
    wire N__44471;
    wire N__44466;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44449;
    wire N__44448;
    wire N__44445;
    wire N__44444;
    wire N__44443;
    wire N__44442;
    wire N__44439;
    wire N__44438;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44426;
    wire N__44423;
    wire N__44422;
    wire N__44421;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44409;
    wire N__44404;
    wire N__44403;
    wire N__44396;
    wire N__44395;
    wire N__44394;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44384;
    wire N__44381;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44363;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44334;
    wire N__44331;
    wire N__44326;
    wire N__44325;
    wire N__44324;
    wire N__44323;
    wire N__44318;
    wire N__44315;
    wire N__44306;
    wire N__44303;
    wire N__44292;
    wire N__44285;
    wire N__44280;
    wire N__44275;
    wire N__44270;
    wire N__44267;
    wire N__44260;
    wire N__44249;
    wire N__44240;
    wire N__44237;
    wire N__44234;
    wire N__44231;
    wire N__44228;
    wire N__44227;
    wire N__44226;
    wire N__44225;
    wire N__44224;
    wire N__44223;
    wire N__44220;
    wire N__44219;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44207;
    wire N__44206;
    wire N__44205;
    wire N__44204;
    wire N__44203;
    wire N__44202;
    wire N__44199;
    wire N__44198;
    wire N__44195;
    wire N__44192;
    wire N__44189;
    wire N__44188;
    wire N__44187;
    wire N__44182;
    wire N__44179;
    wire N__44174;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44159;
    wire N__44156;
    wire N__44153;
    wire N__44152;
    wire N__44151;
    wire N__44150;
    wire N__44149;
    wire N__44148;
    wire N__44143;
    wire N__44140;
    wire N__44139;
    wire N__44134;
    wire N__44133;
    wire N__44122;
    wire N__44121;
    wire N__44118;
    wire N__44113;
    wire N__44108;
    wire N__44105;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44090;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44080;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44061;
    wire N__44060;
    wire N__44055;
    wire N__44050;
    wire N__44047;
    wire N__44044;
    wire N__44039;
    wire N__44038;
    wire N__44037;
    wire N__44030;
    wire N__44029;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43987;
    wire N__43984;
    wire N__43967;
    wire N__43964;
    wire N__43963;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43939;
    wire N__43938;
    wire N__43937;
    wire N__43934;
    wire N__43933;
    wire N__43930;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43881;
    wire N__43876;
    wire N__43873;
    wire N__43870;
    wire N__43865;
    wire N__43862;
    wire N__43861;
    wire N__43860;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43833;
    wire N__43830;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43800;
    wire N__43795;
    wire N__43792;
    wire N__43781;
    wire N__43776;
    wire N__43769;
    wire N__43768;
    wire N__43767;
    wire N__43764;
    wire N__43763;
    wire N__43762;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43754;
    wire N__43751;
    wire N__43748;
    wire N__43747;
    wire N__43744;
    wire N__43741;
    wire N__43736;
    wire N__43733;
    wire N__43730;
    wire N__43729;
    wire N__43728;
    wire N__43727;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43719;
    wire N__43716;
    wire N__43715;
    wire N__43714;
    wire N__43713;
    wire N__43708;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43690;
    wire N__43689;
    wire N__43688;
    wire N__43685;
    wire N__43684;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43676;
    wire N__43675;
    wire N__43674;
    wire N__43673;
    wire N__43670;
    wire N__43669;
    wire N__43668;
    wire N__43667;
    wire N__43666;
    wire N__43665;
    wire N__43664;
    wire N__43661;
    wire N__43654;
    wire N__43653;
    wire N__43650;
    wire N__43647;
    wire N__43642;
    wire N__43639;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43622;
    wire N__43621;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43609;
    wire N__43604;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43588;
    wire N__43587;
    wire N__43586;
    wire N__43585;
    wire N__43584;
    wire N__43583;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43559;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43545;
    wire N__43542;
    wire N__43533;
    wire N__43528;
    wire N__43525;
    wire N__43522;
    wire N__43517;
    wire N__43512;
    wire N__43511;
    wire N__43510;
    wire N__43507;
    wire N__43502;
    wire N__43495;
    wire N__43492;
    wire N__43491;
    wire N__43486;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43460;
    wire N__43455;
    wire N__43448;
    wire N__43443;
    wire N__43438;
    wire N__43429;
    wire N__43426;
    wire N__43419;
    wire N__43400;
    wire N__43397;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43373;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43346;
    wire N__43345;
    wire N__43344;
    wire N__43341;
    wire N__43340;
    wire N__43337;
    wire N__43334;
    wire N__43331;
    wire N__43328;
    wire N__43325;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43301;
    wire N__43298;
    wire N__43295;
    wire N__43292;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43247;
    wire N__43244;
    wire N__43241;
    wire N__43238;
    wire N__43235;
    wire N__43232;
    wire N__43231;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43211;
    wire N__43208;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43189;
    wire N__43186;
    wire N__43185;
    wire N__43184;
    wire N__43181;
    wire N__43180;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43172;
    wire N__43169;
    wire N__43166;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43152;
    wire N__43151;
    wire N__43150;
    wire N__43149;
    wire N__43144;
    wire N__43141;
    wire N__43140;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43125;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43110;
    wire N__43109;
    wire N__43106;
    wire N__43101;
    wire N__43098;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43090;
    wire N__43087;
    wire N__43082;
    wire N__43077;
    wire N__43072;
    wire N__43067;
    wire N__43064;
    wire N__43061;
    wire N__43056;
    wire N__43053;
    wire N__43048;
    wire N__43043;
    wire N__43038;
    wire N__43025;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42997;
    wire N__42996;
    wire N__42995;
    wire N__42994;
    wire N__42993;
    wire N__42992;
    wire N__42991;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42980;
    wire N__42977;
    wire N__42974;
    wire N__42973;
    wire N__42972;
    wire N__42971;
    wire N__42970;
    wire N__42969;
    wire N__42966;
    wire N__42963;
    wire N__42960;
    wire N__42959;
    wire N__42958;
    wire N__42957;
    wire N__42954;
    wire N__42951;
    wire N__42948;
    wire N__42947;
    wire N__42946;
    wire N__42945;
    wire N__42942;
    wire N__42939;
    wire N__42934;
    wire N__42933;
    wire N__42928;
    wire N__42927;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42916;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42906;
    wire N__42905;
    wire N__42904;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42892;
    wire N__42891;
    wire N__42886;
    wire N__42879;
    wire N__42874;
    wire N__42871;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42849;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42823;
    wire N__42822;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42810;
    wire N__42807;
    wire N__42800;
    wire N__42797;
    wire N__42790;
    wire N__42789;
    wire N__42788;
    wire N__42787;
    wire N__42782;
    wire N__42777;
    wire N__42774;
    wire N__42769;
    wire N__42764;
    wire N__42761;
    wire N__42758;
    wire N__42753;
    wire N__42748;
    wire N__42743;
    wire N__42738;
    wire N__42735;
    wire N__42724;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42698;
    wire N__42697;
    wire N__42696;
    wire N__42693;
    wire N__42692;
    wire N__42691;
    wire N__42690;
    wire N__42689;
    wire N__42688;
    wire N__42687;
    wire N__42684;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42676;
    wire N__42675;
    wire N__42668;
    wire N__42667;
    wire N__42666;
    wire N__42663;
    wire N__42662;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42644;
    wire N__42639;
    wire N__42636;
    wire N__42631;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42619;
    wire N__42616;
    wire N__42611;
    wire N__42608;
    wire N__42603;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42587;
    wire N__42584;
    wire N__42577;
    wire N__42572;
    wire N__42563;
    wire N__42560;
    wire N__42557;
    wire N__42554;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42539;
    wire N__42536;
    wire N__42533;
    wire N__42530;
    wire N__42527;
    wire N__42526;
    wire N__42523;
    wire N__42522;
    wire N__42519;
    wire N__42518;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42508;
    wire N__42507;
    wire N__42506;
    wire N__42505;
    wire N__42504;
    wire N__42503;
    wire N__42502;
    wire N__42499;
    wire N__42496;
    wire N__42495;
    wire N__42490;
    wire N__42487;
    wire N__42482;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42464;
    wire N__42463;
    wire N__42460;
    wire N__42459;
    wire N__42458;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42430;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42410;
    wire N__42407;
    wire N__42404;
    wire N__42401;
    wire N__42398;
    wire N__42395;
    wire N__42392;
    wire N__42389;
    wire N__42386;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42359;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42349;
    wire N__42346;
    wire N__42343;
    wire N__42340;
    wire N__42337;
    wire N__42332;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42322;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42311;
    wire N__42308;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42298;
    wire N__42297;
    wire N__42296;
    wire N__42289;
    wire N__42286;
    wire N__42283;
    wire N__42280;
    wire N__42277;
    wire N__42266;
    wire N__42265;
    wire N__42264;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42254;
    wire N__42253;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42233;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42199;
    wire N__42194;
    wire N__42193;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42181;
    wire N__42178;
    wire N__42175;
    wire N__42172;
    wire N__42169;
    wire N__42164;
    wire N__42163;
    wire N__42162;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42151;
    wire N__42150;
    wire N__42147;
    wire N__42146;
    wire N__42139;
    wire N__42136;
    wire N__42133;
    wire N__42130;
    wire N__42127;
    wire N__42126;
    wire N__42119;
    wire N__42114;
    wire N__42111;
    wire N__42108;
    wire N__42103;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42093;
    wire N__42092;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42080;
    wire N__42079;
    wire N__42078;
    wire N__42073;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42045;
    wire N__42038;
    wire N__42035;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42023;
    wire N__42020;
    wire N__42017;
    wire N__42016;
    wire N__42015;
    wire N__42014;
    wire N__42013;
    wire N__42012;
    wire N__42011;
    wire N__42006;
    wire N__42005;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41995;
    wire N__41994;
    wire N__41993;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41979;
    wire N__41978;
    wire N__41977;
    wire N__41976;
    wire N__41975;
    wire N__41974;
    wire N__41973;
    wire N__41966;
    wire N__41963;
    wire N__41960;
    wire N__41959;
    wire N__41956;
    wire N__41955;
    wire N__41952;
    wire N__41947;
    wire N__41944;
    wire N__41943;
    wire N__41942;
    wire N__41941;
    wire N__41938;
    wire N__41931;
    wire N__41928;
    wire N__41927;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41919;
    wire N__41916;
    wire N__41911;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41892;
    wire N__41887;
    wire N__41884;
    wire N__41883;
    wire N__41882;
    wire N__41879;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41861;
    wire N__41860;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41843;
    wire N__41840;
    wire N__41833;
    wire N__41830;
    wire N__41825;
    wire N__41820;
    wire N__41813;
    wire N__41810;
    wire N__41809;
    wire N__41804;
    wire N__41799;
    wire N__41794;
    wire N__41787;
    wire N__41782;
    wire N__41779;
    wire N__41776;
    wire N__41769;
    wire N__41766;
    wire N__41747;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41737;
    wire N__41736;
    wire N__41735;
    wire N__41730;
    wire N__41727;
    wire N__41726;
    wire N__41723;
    wire N__41722;
    wire N__41721;
    wire N__41720;
    wire N__41719;
    wire N__41716;
    wire N__41713;
    wire N__41710;
    wire N__41707;
    wire N__41706;
    wire N__41705;
    wire N__41704;
    wire N__41701;
    wire N__41696;
    wire N__41695;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41671;
    wire N__41668;
    wire N__41667;
    wire N__41664;
    wire N__41659;
    wire N__41654;
    wire N__41649;
    wire N__41646;
    wire N__41641;
    wire N__41638;
    wire N__41635;
    wire N__41628;
    wire N__41625;
    wire N__41620;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41548;
    wire N__41545;
    wire N__41544;
    wire N__41539;
    wire N__41538;
    wire N__41535;
    wire N__41534;
    wire N__41531;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41510;
    wire N__41509;
    wire N__41508;
    wire N__41507;
    wire N__41506;
    wire N__41503;
    wire N__41502;
    wire N__41501;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41490;
    wire N__41489;
    wire N__41488;
    wire N__41487;
    wire N__41486;
    wire N__41479;
    wire N__41478;
    wire N__41477;
    wire N__41476;
    wire N__41475;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41467;
    wire N__41458;
    wire N__41455;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41431;
    wire N__41430;
    wire N__41429;
    wire N__41428;
    wire N__41427;
    wire N__41426;
    wire N__41425;
    wire N__41424;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41413;
    wire N__41410;
    wire N__41409;
    wire N__41400;
    wire N__41399;
    wire N__41396;
    wire N__41391;
    wire N__41382;
    wire N__41375;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41340;
    wire N__41339;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41324;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41306;
    wire N__41301;
    wire N__41294;
    wire N__41293;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41281;
    wire N__41278;
    wire N__41271;
    wire N__41266;
    wire N__41261;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41244;
    wire N__41231;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41220;
    wire N__41219;
    wire N__41218;
    wire N__41215;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41207;
    wire N__41206;
    wire N__41205;
    wire N__41204;
    wire N__41203;
    wire N__41202;
    wire N__41201;
    wire N__41200;
    wire N__41199;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41183;
    wire N__41178;
    wire N__41163;
    wire N__41160;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41128;
    wire N__41123;
    wire N__41114;
    wire N__41113;
    wire N__41112;
    wire N__41109;
    wire N__41108;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41063;
    wire N__41062;
    wire N__41061;
    wire N__41060;
    wire N__41059;
    wire N__41058;
    wire N__41057;
    wire N__41056;
    wire N__41055;
    wire N__41054;
    wire N__41053;
    wire N__41052;
    wire N__41027;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40999;
    wire N__40998;
    wire N__40995;
    wire N__40994;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40981;
    wire N__40980;
    wire N__40979;
    wire N__40976;
    wire N__40969;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40959;
    wire N__40956;
    wire N__40951;
    wire N__40946;
    wire N__40943;
    wire N__40940;
    wire N__40937;
    wire N__40932;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40898;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40886;
    wire N__40883;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40862;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40849;
    wire N__40848;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40826;
    wire N__40823;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40805;
    wire N__40802;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40768;
    wire N__40767;
    wire N__40766;
    wire N__40765;
    wire N__40764;
    wire N__40763;
    wire N__40760;
    wire N__40753;
    wire N__40752;
    wire N__40751;
    wire N__40748;
    wire N__40747;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40718;
    wire N__40715;
    wire N__40712;
    wire N__40711;
    wire N__40708;
    wire N__40701;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40685;
    wire N__40682;
    wire N__40679;
    wire N__40674;
    wire N__40671;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40628;
    wire N__40627;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40617;
    wire N__40616;
    wire N__40615;
    wire N__40614;
    wire N__40611;
    wire N__40606;
    wire N__40601;
    wire N__40600;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40579;
    wire N__40574;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40526;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40432;
    wire N__40431;
    wire N__40430;
    wire N__40429;
    wire N__40428;
    wire N__40427;
    wire N__40426;
    wire N__40425;
    wire N__40424;
    wire N__40423;
    wire N__40420;
    wire N__40419;
    wire N__40414;
    wire N__40411;
    wire N__40410;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40402;
    wire N__40401;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40391;
    wire N__40390;
    wire N__40389;
    wire N__40388;
    wire N__40385;
    wire N__40380;
    wire N__40377;
    wire N__40372;
    wire N__40369;
    wire N__40368;
    wire N__40367;
    wire N__40366;
    wire N__40363;
    wire N__40362;
    wire N__40357;
    wire N__40354;
    wire N__40351;
    wire N__40348;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40319;
    wire N__40316;
    wire N__40311;
    wire N__40306;
    wire N__40301;
    wire N__40298;
    wire N__40293;
    wire N__40292;
    wire N__40291;
    wire N__40288;
    wire N__40283;
    wire N__40278;
    wire N__40277;
    wire N__40276;
    wire N__40271;
    wire N__40266;
    wire N__40263;
    wire N__40258;
    wire N__40253;
    wire N__40246;
    wire N__40241;
    wire N__40236;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40120;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40112;
    wire N__40111;
    wire N__40108;
    wire N__40107;
    wire N__40104;
    wire N__40103;
    wire N__40102;
    wire N__40099;
    wire N__40098;
    wire N__40095;
    wire N__40094;
    wire N__40093;
    wire N__40090;
    wire N__40087;
    wire N__40086;
    wire N__40085;
    wire N__40084;
    wire N__40083;
    wire N__40082;
    wire N__40081;
    wire N__40080;
    wire N__40079;
    wire N__40076;
    wire N__40075;
    wire N__40072;
    wire N__40071;
    wire N__40070;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40046;
    wire N__40045;
    wire N__40044;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40032;
    wire N__40029;
    wire N__40022;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40001;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39979;
    wire N__39976;
    wire N__39971;
    wire N__39968;
    wire N__39963;
    wire N__39960;
    wire N__39953;
    wire N__39950;
    wire N__39943;
    wire N__39940;
    wire N__39933;
    wire N__39928;
    wire N__39923;
    wire N__39920;
    wire N__39913;
    wire N__39904;
    wire N__39899;
    wire N__39890;
    wire N__39887;
    wire N__39884;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39860;
    wire N__39859;
    wire N__39856;
    wire N__39855;
    wire N__39854;
    wire N__39853;
    wire N__39852;
    wire N__39851;
    wire N__39850;
    wire N__39849;
    wire N__39848;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39838;
    wire N__39837;
    wire N__39836;
    wire N__39833;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39825;
    wire N__39822;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39814;
    wire N__39809;
    wire N__39808;
    wire N__39807;
    wire N__39804;
    wire N__39799;
    wire N__39796;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39753;
    wire N__39752;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39740;
    wire N__39737;
    wire N__39734;
    wire N__39731;
    wire N__39728;
    wire N__39725;
    wire N__39722;
    wire N__39717;
    wire N__39712;
    wire N__39709;
    wire N__39704;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39681;
    wire N__39676;
    wire N__39665;
    wire N__39656;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39607;
    wire N__39606;
    wire N__39605;
    wire N__39602;
    wire N__39601;
    wire N__39600;
    wire N__39599;
    wire N__39596;
    wire N__39595;
    wire N__39594;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39586;
    wire N__39579;
    wire N__39572;
    wire N__39571;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39540;
    wire N__39537;
    wire N__39532;
    wire N__39531;
    wire N__39528;
    wire N__39525;
    wire N__39518;
    wire N__39515;
    wire N__39506;
    wire N__39503;
    wire N__39500;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39472;
    wire N__39471;
    wire N__39468;
    wire N__39467;
    wire N__39464;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39453;
    wire N__39452;
    wire N__39449;
    wire N__39448;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39440;
    wire N__39435;
    wire N__39430;
    wire N__39427;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39398;
    wire N__39397;
    wire N__39396;
    wire N__39395;
    wire N__39394;
    wire N__39391;
    wire N__39390;
    wire N__39389;
    wire N__39388;
    wire N__39387;
    wire N__39386;
    wire N__39385;
    wire N__39384;
    wire N__39383;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39359;
    wire N__39356;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39323;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39308;
    wire N__39301;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39286;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39260;
    wire N__39253;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39232;
    wire N__39229;
    wire N__39224;
    wire N__39219;
    wire N__39212;
    wire N__39209;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39181;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39157;
    wire N__39152;
    wire N__39151;
    wire N__39150;
    wire N__39149;
    wire N__39148;
    wire N__39147;
    wire N__39146;
    wire N__39145;
    wire N__39144;
    wire N__39143;
    wire N__39142;
    wire N__39141;
    wire N__39140;
    wire N__39139;
    wire N__39134;
    wire N__39129;
    wire N__39122;
    wire N__39117;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39088;
    wire N__39085;
    wire N__39084;
    wire N__39083;
    wire N__39082;
    wire N__39081;
    wire N__39080;
    wire N__39079;
    wire N__39078;
    wire N__39077;
    wire N__39076;
    wire N__39071;
    wire N__39070;
    wire N__39069;
    wire N__39062;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39054;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39046;
    wire N__39045;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39037;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39022;
    wire N__39019;
    wire N__39018;
    wire N__39017;
    wire N__39016;
    wire N__39015;
    wire N__39014;
    wire N__39013;
    wire N__39012;
    wire N__39011;
    wire N__39010;
    wire N__39007;
    wire N__39006;
    wire N__39005;
    wire N__39002;
    wire N__38995;
    wire N__38986;
    wire N__38975;
    wire N__38974;
    wire N__38973;
    wire N__38972;
    wire N__38971;
    wire N__38970;
    wire N__38969;
    wire N__38968;
    wire N__38967;
    wire N__38966;
    wire N__38965;
    wire N__38962;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38923;
    wire N__38922;
    wire N__38919;
    wire N__38912;
    wire N__38907;
    wire N__38902;
    wire N__38897;
    wire N__38892;
    wire N__38889;
    wire N__38888;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38868;
    wire N__38865;
    wire N__38860;
    wire N__38855;
    wire N__38850;
    wire N__38847;
    wire N__38840;
    wire N__38835;
    wire N__38822;
    wire N__38819;
    wire N__38814;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38794;
    wire N__38785;
    wire N__38782;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38744;
    wire N__38743;
    wire N__38740;
    wire N__38739;
    wire N__38736;
    wire N__38735;
    wire N__38734;
    wire N__38733;
    wire N__38732;
    wire N__38731;
    wire N__38730;
    wire N__38729;
    wire N__38728;
    wire N__38727;
    wire N__38726;
    wire N__38725;
    wire N__38724;
    wire N__38723;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38715;
    wire N__38714;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38697;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38689;
    wire N__38686;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38678;
    wire N__38677;
    wire N__38676;
    wire N__38673;
    wire N__38668;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38653;
    wire N__38652;
    wire N__38649;
    wire N__38648;
    wire N__38647;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38593;
    wire N__38592;
    wire N__38591;
    wire N__38584;
    wire N__38579;
    wire N__38576;
    wire N__38571;
    wire N__38566;
    wire N__38561;
    wire N__38560;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38548;
    wire N__38541;
    wire N__38540;
    wire N__38529;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38517;
    wire N__38514;
    wire N__38509;
    wire N__38504;
    wire N__38495;
    wire N__38490;
    wire N__38485;
    wire N__38480;
    wire N__38477;
    wire N__38474;
    wire N__38469;
    wire N__38444;
    wire N__38441;
    wire N__38438;
    wire N__38437;
    wire N__38436;
    wire N__38433;
    wire N__38432;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38417;
    wire N__38414;
    wire N__38405;
    wire N__38402;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38375;
    wire N__38372;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38350;
    wire N__38345;
    wire N__38342;
    wire N__38339;
    wire N__38338;
    wire N__38337;
    wire N__38336;
    wire N__38333;
    wire N__38332;
    wire N__38331;
    wire N__38330;
    wire N__38329;
    wire N__38326;
    wire N__38325;
    wire N__38324;
    wire N__38323;
    wire N__38322;
    wire N__38319;
    wire N__38318;
    wire N__38317;
    wire N__38316;
    wire N__38315;
    wire N__38312;
    wire N__38311;
    wire N__38310;
    wire N__38309;
    wire N__38308;
    wire N__38307;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38299;
    wire N__38292;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38275;
    wire N__38274;
    wire N__38273;
    wire N__38272;
    wire N__38269;
    wire N__38264;
    wire N__38257;
    wire N__38250;
    wire N__38249;
    wire N__38248;
    wire N__38247;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38226;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38214;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38192;
    wire N__38191;
    wire N__38190;
    wire N__38183;
    wire N__38180;
    wire N__38179;
    wire N__38178;
    wire N__38177;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38163;
    wire N__38158;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38131;
    wire N__38126;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38100;
    wire N__38095;
    wire N__38092;
    wire N__38085;
    wire N__38076;
    wire N__38051;
    wire N__38048;
    wire N__38047;
    wire N__38046;
    wire N__38045;
    wire N__38042;
    wire N__38041;
    wire N__38038;
    wire N__38037;
    wire N__38036;
    wire N__38035;
    wire N__38034;
    wire N__38033;
    wire N__38030;
    wire N__38029;
    wire N__38028;
    wire N__38027;
    wire N__38026;
    wire N__38025;
    wire N__38024;
    wire N__38023;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38006;
    wire N__38003;
    wire N__38002;
    wire N__38001;
    wire N__37998;
    wire N__37997;
    wire N__37996;
    wire N__37995;
    wire N__37994;
    wire N__37987;
    wire N__37986;
    wire N__37985;
    wire N__37982;
    wire N__37981;
    wire N__37976;
    wire N__37969;
    wire N__37968;
    wire N__37963;
    wire N__37962;
    wire N__37961;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37937;
    wire N__37936;
    wire N__37935;
    wire N__37934;
    wire N__37933;
    wire N__37926;
    wire N__37923;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37883;
    wire N__37876;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37856;
    wire N__37847;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37827;
    wire N__37824;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37773;
    wire N__37770;
    wire N__37769;
    wire N__37768;
    wire N__37767;
    wire N__37764;
    wire N__37763;
    wire N__37762;
    wire N__37761;
    wire N__37760;
    wire N__37759;
    wire N__37758;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37746;
    wire N__37743;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37733;
    wire N__37732;
    wire N__37731;
    wire N__37730;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37718;
    wire N__37717;
    wire N__37716;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37704;
    wire N__37703;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37693;
    wire N__37688;
    wire N__37683;
    wire N__37680;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37664;
    wire N__37661;
    wire N__37660;
    wire N__37659;
    wire N__37658;
    wire N__37657;
    wire N__37656;
    wire N__37655;
    wire N__37654;
    wire N__37653;
    wire N__37652;
    wire N__37651;
    wire N__37648;
    wire N__37647;
    wire N__37646;
    wire N__37641;
    wire N__37636;
    wire N__37633;
    wire N__37628;
    wire N__37627;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37603;
    wire N__37596;
    wire N__37593;
    wire N__37586;
    wire N__37583;
    wire N__37578;
    wire N__37575;
    wire N__37570;
    wire N__37567;
    wire N__37560;
    wire N__37555;
    wire N__37538;
    wire N__37533;
    wire N__37514;
    wire N__37513;
    wire N__37510;
    wire N__37507;
    wire N__37504;
    wire N__37503;
    wire N__37502;
    wire N__37501;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37490;
    wire N__37489;
    wire N__37488;
    wire N__37487;
    wire N__37486;
    wire N__37485;
    wire N__37484;
    wire N__37481;
    wire N__37480;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37468;
    wire N__37463;
    wire N__37456;
    wire N__37451;
    wire N__37448;
    wire N__37447;
    wire N__37444;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37429;
    wire N__37428;
    wire N__37427;
    wire N__37426;
    wire N__37425;
    wire N__37420;
    wire N__37419;
    wire N__37418;
    wire N__37417;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37392;
    wire N__37391;
    wire N__37388;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37376;
    wire N__37373;
    wire N__37372;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37349;
    wire N__37348;
    wire N__37347;
    wire N__37342;
    wire N__37339;
    wire N__37334;
    wire N__37329;
    wire N__37326;
    wire N__37319;
    wire N__37318;
    wire N__37313;
    wire N__37302;
    wire N__37295;
    wire N__37290;
    wire N__37287;
    wire N__37280;
    wire N__37277;
    wire N__37272;
    wire N__37259;
    wire N__37256;
    wire N__37255;
    wire N__37254;
    wire N__37251;
    wire N__37246;
    wire N__37245;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37237;
    wire N__37236;
    wire N__37235;
    wire N__37234;
    wire N__37233;
    wire N__37232;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37218;
    wire N__37215;
    wire N__37214;
    wire N__37211;
    wire N__37206;
    wire N__37205;
    wire N__37204;
    wire N__37203;
    wire N__37202;
    wire N__37201;
    wire N__37200;
    wire N__37199;
    wire N__37196;
    wire N__37195;
    wire N__37194;
    wire N__37191;
    wire N__37188;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37169;
    wire N__37164;
    wire N__37159;
    wire N__37158;
    wire N__37157;
    wire N__37156;
    wire N__37153;
    wire N__37146;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37118;
    wire N__37117;
    wire N__37116;
    wire N__37115;
    wire N__37114;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37098;
    wire N__37095;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37069;
    wire N__37064;
    wire N__37059;
    wire N__37052;
    wire N__37049;
    wire N__37044;
    wire N__37037;
    wire N__37030;
    wire N__37021;
    wire N__37004;
    wire N__37003;
    wire N__37002;
    wire N__37001;
    wire N__37000;
    wire N__36999;
    wire N__36998;
    wire N__36997;
    wire N__36996;
    wire N__36995;
    wire N__36994;
    wire N__36993;
    wire N__36990;
    wire N__36989;
    wire N__36986;
    wire N__36985;
    wire N__36984;
    wire N__36983;
    wire N__36982;
    wire N__36981;
    wire N__36980;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36967;
    wire N__36966;
    wire N__36965;
    wire N__36964;
    wire N__36963;
    wire N__36962;
    wire N__36959;
    wire N__36958;
    wire N__36957;
    wire N__36954;
    wire N__36953;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36945;
    wire N__36944;
    wire N__36941;
    wire N__36940;
    wire N__36939;
    wire N__36938;
    wire N__36937;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36925;
    wire N__36922;
    wire N__36915;
    wire N__36912;
    wire N__36905;
    wire N__36902;
    wire N__36897;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36879;
    wire N__36878;
    wire N__36875;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36852;
    wire N__36845;
    wire N__36844;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36828;
    wire N__36825;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36813;
    wire N__36804;
    wire N__36801;
    wire N__36796;
    wire N__36791;
    wire N__36784;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36765;
    wire N__36760;
    wire N__36757;
    wire N__36754;
    wire N__36751;
    wire N__36748;
    wire N__36741;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36709;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36622;
    wire N__36617;
    wire N__36614;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36592;
    wire N__36591;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36554;
    wire N__36553;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36518;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36466;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36433;
    wire N__36430;
    wire N__36427;
    wire N__36424;
    wire N__36419;
    wire N__36416;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36395;
    wire N__36392;
    wire N__36391;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36329;
    wire N__36326;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36268;
    wire N__36265;
    wire N__36264;
    wire N__36261;
    wire N__36260;
    wire N__36259;
    wire N__36258;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36231;
    wire N__36228;
    wire N__36223;
    wire N__36218;
    wire N__36209;
    wire N__36206;
    wire N__36205;
    wire N__36204;
    wire N__36203;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36147;
    wire N__36140;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36124;
    wire N__36123;
    wire N__36120;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36104;
    wire N__36101;
    wire N__36100;
    wire N__36097;
    wire N__36094;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36046;
    wire N__36043;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36020;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36005;
    wire N__36004;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35989;
    wire N__35986;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35966;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35923;
    wire N__35912;
    wire N__35911;
    wire N__35910;
    wire N__35907;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35894;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35876;
    wire N__35875;
    wire N__35872;
    wire N__35871;
    wire N__35870;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35853;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35841;
    wire N__35838;
    wire N__35833;
    wire N__35830;
    wire N__35823;
    wire N__35810;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35798;
    wire N__35795;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35762;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35754;
    wire N__35753;
    wire N__35752;
    wire N__35749;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35738;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35713;
    wire N__35710;
    wire N__35709;
    wire N__35708;
    wire N__35707;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35699;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35672;
    wire N__35671;
    wire N__35668;
    wire N__35663;
    wire N__35658;
    wire N__35653;
    wire N__35648;
    wire N__35645;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35615;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35599;
    wire N__35596;
    wire N__35591;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35583;
    wire N__35582;
    wire N__35581;
    wire N__35578;
    wire N__35577;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35532;
    wire N__35531;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35488;
    wire N__35483;
    wire N__35478;
    wire N__35475;
    wire N__35462;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35447;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35435;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35410;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35396;
    wire N__35395;
    wire N__35394;
    wire N__35391;
    wire N__35386;
    wire N__35385;
    wire N__35384;
    wire N__35379;
    wire N__35378;
    wire N__35377;
    wire N__35376;
    wire N__35375;
    wire N__35374;
    wire N__35371;
    wire N__35368;
    wire N__35367;
    wire N__35366;
    wire N__35365;
    wire N__35362;
    wire N__35357;
    wire N__35356;
    wire N__35353;
    wire N__35352;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35303;
    wire N__35300;
    wire N__35299;
    wire N__35298;
    wire N__35297;
    wire N__35294;
    wire N__35289;
    wire N__35280;
    wire N__35275;
    wire N__35272;
    wire N__35265;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35242;
    wire N__35241;
    wire N__35236;
    wire N__35233;
    wire N__35232;
    wire N__35231;
    wire N__35230;
    wire N__35229;
    wire N__35226;
    wire N__35225;
    wire N__35224;
    wire N__35223;
    wire N__35222;
    wire N__35221;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35202;
    wire N__35199;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35187;
    wire N__35184;
    wire N__35183;
    wire N__35180;
    wire N__35175;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35135;
    wire N__35134;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35102;
    wire N__35097;
    wire N__35094;
    wire N__35087;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35033;
    wire N__35032;
    wire N__35031;
    wire N__35030;
    wire N__35029;
    wire N__35028;
    wire N__35027;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34995;
    wire N__34994;
    wire N__34993;
    wire N__34988;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34947;
    wire N__34934;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34884;
    wire N__34883;
    wire N__34882;
    wire N__34877;
    wire N__34872;
    wire N__34869;
    wire N__34868;
    wire N__34867;
    wire N__34864;
    wire N__34863;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34855;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34827;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34787;
    wire N__34784;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34770;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34764;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34748;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34721;
    wire N__34720;
    wire N__34717;
    wire N__34716;
    wire N__34715;
    wire N__34714;
    wire N__34711;
    wire N__34710;
    wire N__34709;
    wire N__34708;
    wire N__34705;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34691;
    wire N__34688;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34682;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34657;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34617;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34605;
    wire N__34604;
    wire N__34601;
    wire N__34594;
    wire N__34589;
    wire N__34582;
    wire N__34579;
    wire N__34568;
    wire N__34567;
    wire N__34566;
    wire N__34563;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34509;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34497;
    wire N__34496;
    wire N__34495;
    wire N__34494;
    wire N__34489;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34475;
    wire N__34474;
    wire N__34473;
    wire N__34470;
    wire N__34469;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34454;
    wire N__34447;
    wire N__34444;
    wire N__34439;
    wire N__34434;
    wire N__34431;
    wire N__34424;
    wire N__34415;
    wire N__34412;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34404;
    wire N__34403;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34395;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34364;
    wire N__34361;
    wire N__34346;
    wire N__34345;
    wire N__34344;
    wire N__34343;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34326;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34310;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34288;
    wire N__34283;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34269;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34250;
    wire N__34249;
    wire N__34248;
    wire N__34247;
    wire N__34246;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34215;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34190;
    wire N__34181;
    wire N__34180;
    wire N__34179;
    wire N__34176;
    wire N__34175;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34128;
    wire N__34125;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34094;
    wire N__34091;
    wire N__34090;
    wire N__34089;
    wire N__34088;
    wire N__34087;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34031;
    wire N__34030;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34022;
    wire N__34021;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33962;
    wire N__33959;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33940;
    wire N__33939;
    wire N__33936;
    wire N__33935;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33921;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33906;
    wire N__33903;
    wire N__33900;
    wire N__33895;
    wire N__33890;
    wire N__33881;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33873;
    wire N__33872;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33864;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33853;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33834;
    wire N__33831;
    wire N__33818;
    wire N__33817;
    wire N__33816;
    wire N__33815;
    wire N__33814;
    wire N__33813;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33758;
    wire N__33757;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33749;
    wire N__33748;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33713;
    wire N__33708;
    wire N__33705;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33662;
    wire N__33661;
    wire N__33660;
    wire N__33659;
    wire N__33656;
    wire N__33655;
    wire N__33654;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33623;
    wire N__33620;
    wire N__33615;
    wire N__33612;
    wire N__33605;
    wire N__33604;
    wire N__33603;
    wire N__33602;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33591;
    wire N__33590;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33557;
    wire N__33552;
    wire N__33539;
    wire N__33536;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33476;
    wire N__33473;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33442;
    wire N__33439;
    wire N__33438;
    wire N__33435;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33385;
    wire N__33384;
    wire N__33381;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33362;
    wire N__33359;
    wire N__33358;
    wire N__33357;
    wire N__33356;
    wire N__33355;
    wire N__33354;
    wire N__33351;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33335;
    wire N__33332;
    wire N__33331;
    wire N__33330;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33318;
    wire N__33317;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33303;
    wire N__33302;
    wire N__33301;
    wire N__33300;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33287;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33275;
    wire N__33272;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33264;
    wire N__33263;
    wire N__33262;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33246;
    wire N__33245;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33227;
    wire N__33220;
    wire N__33213;
    wire N__33210;
    wire N__33205;
    wire N__33200;
    wire N__33197;
    wire N__33192;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33149;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33089;
    wire N__33086;
    wire N__33085;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33065;
    wire N__33064;
    wire N__33063;
    wire N__33062;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__32996;
    wire N__32995;
    wire N__32994;
    wire N__32993;
    wire N__32992;
    wire N__32991;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32983;
    wire N__32980;
    wire N__32975;
    wire N__32972;
    wire N__32971;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32963;
    wire N__32960;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32885;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32840;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32798;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32767;
    wire N__32764;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32716;
    wire N__32715;
    wire N__32712;
    wire N__32707;
    wire N__32704;
    wire N__32701;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32670;
    wire N__32667;
    wire N__32666;
    wire N__32665;
    wire N__32662;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32627;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32608;
    wire N__32605;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32585;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32471;
    wire N__32468;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32444;
    wire N__32439;
    wire N__32436;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32363;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32327;
    wire N__32326;
    wire N__32323;
    wire N__32322;
    wire N__32321;
    wire N__32320;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32308;
    wire N__32303;
    wire N__32294;
    wire N__32293;
    wire N__32292;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32228;
    wire N__32225;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32215;
    wire N__32214;
    wire N__32213;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32193;
    wire N__32188;
    wire N__32185;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32080;
    wire N__32079;
    wire N__32074;
    wire N__32073;
    wire N__32070;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32066;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32049;
    wire N__32044;
    wire N__32041;
    wire N__32040;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32028;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32011;
    wire N__32006;
    wire N__31999;
    wire N__31992;
    wire N__31987;
    wire N__31984;
    wire N__31979;
    wire N__31964;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31922;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31901;
    wire N__31898;
    wire N__31895;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31883;
    wire N__31880;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31862;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31772;
    wire N__31771;
    wire N__31768;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31751;
    wire N__31748;
    wire N__31745;
    wire N__31742;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31597;
    wire N__31594;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31502;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31442;
    wire N__31441;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31423;
    wire N__31420;
    wire N__31417;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31396;
    wire N__31393;
    wire N__31390;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31264;
    wire N__31263;
    wire N__31262;
    wire N__31261;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31250;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31198;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31180;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31157;
    wire N__31154;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31046;
    wire N__31045;
    wire N__31044;
    wire N__31043;
    wire N__31042;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31015;
    wire N__31014;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__30999;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30983;
    wire N__30974;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30941;
    wire N__30938;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30809;
    wire N__30808;
    wire N__30807;
    wire N__30806;
    wire N__30805;
    wire N__30802;
    wire N__30797;
    wire N__30794;
    wire N__30789;
    wire N__30784;
    wire N__30783;
    wire N__30782;
    wire N__30781;
    wire N__30780;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30750;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30635;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30623;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30610;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30557;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30539;
    wire N__30536;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30479;
    wire N__30478;
    wire N__30477;
    wire N__30472;
    wire N__30471;
    wire N__30470;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30455;
    wire N__30452;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30418;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30386;
    wire N__30385;
    wire N__30384;
    wire N__30381;
    wire N__30380;
    wire N__30379;
    wire N__30378;
    wire N__30377;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30359;
    wire N__30356;
    wire N__30349;
    wire N__30346;
    wire N__30341;
    wire N__30338;
    wire N__30337;
    wire N__30336;
    wire N__30333;
    wire N__30328;
    wire N__30323;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30315;
    wire N__30314;
    wire N__30311;
    wire N__30306;
    wire N__30303;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30292;
    wire N__30291;
    wire N__30290;
    wire N__30289;
    wire N__30286;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30269;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30253;
    wire N__30250;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30223;
    wire N__30218;
    wire N__30217;
    wire N__30216;
    wire N__30215;
    wire N__30212;
    wire N__30211;
    wire N__30208;
    wire N__30207;
    wire N__30206;
    wire N__30205;
    wire N__30202;
    wire N__30201;
    wire N__30200;
    wire N__30197;
    wire N__30196;
    wire N__30195;
    wire N__30194;
    wire N__30193;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30181;
    wire N__30176;
    wire N__30173;
    wire N__30172;
    wire N__30171;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30153;
    wire N__30148;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30136;
    wire N__30135;
    wire N__30132;
    wire N__30131;
    wire N__30130;
    wire N__30129;
    wire N__30122;
    wire N__30117;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30098;
    wire N__30093;
    wire N__30090;
    wire N__30083;
    wire N__30074;
    wire N__30059;
    wire N__30058;
    wire N__30057;
    wire N__30056;
    wire N__30055;
    wire N__30054;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30046;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30032;
    wire N__30031;
    wire N__30030;
    wire N__30027;
    wire N__30026;
    wire N__30025;
    wire N__30024;
    wire N__30023;
    wire N__30022;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30014;
    wire N__30013;
    wire N__30012;
    wire N__30007;
    wire N__30002;
    wire N__29995;
    wire N__29994;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29956;
    wire N__29955;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29926;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29898;
    wire N__29891;
    wire N__29888;
    wire N__29883;
    wire N__29880;
    wire N__29875;
    wire N__29870;
    wire N__29865;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29837;
    wire N__29836;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29818;
    wire N__29815;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29788;
    wire N__29785;
    wire N__29780;
    wire N__29773;
    wire N__29756;
    wire N__29755;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29746;
    wire N__29745;
    wire N__29742;
    wire N__29741;
    wire N__29740;
    wire N__29739;
    wire N__29736;
    wire N__29735;
    wire N__29730;
    wire N__29729;
    wire N__29728;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29703;
    wire N__29702;
    wire N__29701;
    wire N__29698;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29688;
    wire N__29683;
    wire N__29682;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29678;
    wire N__29673;
    wire N__29668;
    wire N__29659;
    wire N__29654;
    wire N__29649;
    wire N__29644;
    wire N__29639;
    wire N__29632;
    wire N__29623;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29587;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29521;
    wire N__29520;
    wire N__29519;
    wire N__29518;
    wire N__29517;
    wire N__29514;
    wire N__29507;
    wire N__29502;
    wire N__29495;
    wire N__29494;
    wire N__29493;
    wire N__29492;
    wire N__29491;
    wire N__29490;
    wire N__29483;
    wire N__29480;
    wire N__29475;
    wire N__29468;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29437;
    wire N__29436;
    wire N__29435;
    wire N__29434;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29413;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29405;
    wire N__29404;
    wire N__29403;
    wire N__29402;
    wire N__29399;
    wire N__29394;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29380;
    wire N__29379;
    wire N__29378;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29367;
    wire N__29362;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29342;
    wire N__29339;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29316;
    wire N__29311;
    wire N__29310;
    wire N__29309;
    wire N__29306;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29292;
    wire N__29289;
    wire N__29284;
    wire N__29279;
    wire N__29276;
    wire N__29267;
    wire N__29266;
    wire N__29263;
    wire N__29262;
    wire N__29261;
    wire N__29258;
    wire N__29251;
    wire N__29250;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29238;
    wire N__29235;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29219;
    wire N__29216;
    wire N__29215;
    wire N__29210;
    wire N__29207;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29195;
    wire N__29194;
    wire N__29193;
    wire N__29190;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29171;
    wire N__29168;
    wire N__29167;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29072;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29051;
    wire N__29048;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29015;
    wire N__29012;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28979;
    wire N__28976;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28952;
    wire N__28949;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28909;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28781;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28759;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28703;
    wire N__28700;
    wire N__28697;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28636;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28601;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28565;
    wire N__28562;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28496;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28426;
    wire N__28423;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28394;
    wire N__28391;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28159;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28141;
    wire N__28138;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28126;
    wire N__28125;
    wire N__28122;
    wire N__28117;
    wire N__28114;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28090;
    wire N__28089;
    wire N__28088;
    wire N__28087;
    wire N__28086;
    wire N__28085;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28071;
    wire N__28070;
    wire N__28069;
    wire N__28068;
    wire N__28065;
    wire N__28060;
    wire N__28057;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28036;
    wire N__28035;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28027;
    wire N__28026;
    wire N__28025;
    wire N__28020;
    wire N__28015;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__27999;
    wire N__27996;
    wire N__27991;
    wire N__27988;
    wire N__27983;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27898;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27883;
    wire N__27880;
    wire N__27875;
    wire N__27874;
    wire N__27871;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27802;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27728;
    wire N__27727;
    wire N__27724;
    wire N__27723;
    wire N__27720;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27607;
    wire N__27604;
    wire N__27603;
    wire N__27602;
    wire N__27601;
    wire N__27600;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27596;
    wire N__27595;
    wire N__27594;
    wire N__27593;
    wire N__27590;
    wire N__27589;
    wire N__27588;
    wire N__27587;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27570;
    wire N__27567;
    wire N__27566;
    wire N__27559;
    wire N__27558;
    wire N__27555;
    wire N__27554;
    wire N__27551;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27536;
    wire N__27535;
    wire N__27534;
    wire N__27531;
    wire N__27526;
    wire N__27521;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27511;
    wire N__27508;
    wire N__27503;
    wire N__27500;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27446;
    wire N__27443;
    wire N__27436;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27414;
    wire N__27405;
    wire N__27400;
    wire N__27395;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27349;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27338;
    wire N__27337;
    wire N__27336;
    wire N__27331;
    wire N__27326;
    wire N__27325;
    wire N__27322;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27304;
    wire N__27299;
    wire N__27296;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27196;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27185;
    wire N__27182;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27155;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27134;
    wire N__27133;
    wire N__27132;
    wire N__27131;
    wire N__27130;
    wire N__27129;
    wire N__27128;
    wire N__27127;
    wire N__27126;
    wire N__27125;
    wire N__27124;
    wire N__27121;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27109;
    wire N__27108;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27062;
    wire N__27059;
    wire N__27054;
    wire N__27041;
    wire N__27040;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27029;
    wire N__27028;
    wire N__27027;
    wire N__27026;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26997;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26945;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26881;
    wire N__26880;
    wire N__26879;
    wire N__26874;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26828;
    wire N__26827;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26750;
    wire N__26747;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26729;
    wire N__26728;
    wire N__26727;
    wire N__26722;
    wire N__26717;
    wire N__26716;
    wire N__26715;
    wire N__26712;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26690;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26678;
    wire N__26673;
    wire N__26668;
    wire N__26665;
    wire N__26660;
    wire N__26651;
    wire N__26650;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26627;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26605;
    wire N__26604;
    wire N__26603;
    wire N__26602;
    wire N__26601;
    wire N__26600;
    wire N__26599;
    wire N__26598;
    wire N__26597;
    wire N__26596;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26588;
    wire N__26583;
    wire N__26578;
    wire N__26577;
    wire N__26576;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26568;
    wire N__26565;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26554;
    wire N__26553;
    wire N__26550;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26535;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26523;
    wire N__26518;
    wire N__26515;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26503;
    wire N__26500;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26496;
    wire N__26495;
    wire N__26494;
    wire N__26487;
    wire N__26484;
    wire N__26477;
    wire N__26468;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26428;
    wire N__26425;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26380;
    wire N__26379;
    wire N__26376;
    wire N__26375;
    wire N__26370;
    wire N__26363;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26346;
    wire N__26341;
    wire N__26334;
    wire N__26329;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26303;
    wire N__26298;
    wire N__26285;
    wire N__26284;
    wire N__26283;
    wire N__26282;
    wire N__26281;
    wire N__26280;
    wire N__26279;
    wire N__26278;
    wire N__26277;
    wire N__26276;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26259;
    wire N__26254;
    wire N__26253;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26237;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26201;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26059;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25631;
    wire N__25628;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25538;
    wire N__25535;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25506;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25462;
    wire N__25461;
    wire N__25454;
    wire N__25453;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25442;
    wire N__25439;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25423;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25378;
    wire N__25377;
    wire N__25374;
    wire N__25373;
    wire N__25372;
    wire N__25371;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25356;
    wire N__25355;
    wire N__25354;
    wire N__25353;
    wire N__25352;
    wire N__25349;
    wire N__25348;
    wire N__25345;
    wire N__25344;
    wire N__25343;
    wire N__25342;
    wire N__25341;
    wire N__25340;
    wire N__25335;
    wire N__25330;
    wire N__25327;
    wire N__25326;
    wire N__25323;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25290;
    wire N__25289;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25274;
    wire N__25269;
    wire N__25264;
    wire N__25259;
    wire N__25252;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25225;
    wire N__25222;
    wire N__25221;
    wire N__25220;
    wire N__25217;
    wire N__25216;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25206;
    wire N__25205;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25170;
    wire N__25169;
    wire N__25166;
    wire N__25165;
    wire N__25164;
    wire N__25159;
    wire N__25156;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25140;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25123;
    wire N__25122;
    wire N__25119;
    wire N__25118;
    wire N__25111;
    wire N__25108;
    wire N__25103;
    wire N__25100;
    wire N__25091;
    wire N__25084;
    wire N__25079;
    wire N__25076;
    wire N__25061;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25053;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25039;
    wire N__25036;
    wire N__25031;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25013;
    wire N__25010;
    wire N__25009;
    wire N__25008;
    wire N__25003;
    wire N__25000;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24985;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24973;
    wire N__24970;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24906;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24872;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24853;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24772;
    wire N__24769;
    wire N__24768;
    wire N__24767;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24753;
    wire N__24746;
    wire N__24743;
    wire N__24742;
    wire N__24741;
    wire N__24740;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24723;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24711;
    wire N__24708;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24688;
    wire N__24683;
    wire N__24682;
    wire N__24681;
    wire N__24680;
    wire N__24677;
    wire N__24670;
    wire N__24667;
    wire N__24662;
    wire N__24661;
    wire N__24660;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24645;
    wire N__24636;
    wire N__24633;
    wire N__24632;
    wire N__24631;
    wire N__24628;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24612;
    wire N__24609;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24595;
    wire N__24594;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24580;
    wire N__24579;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24563;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24515;
    wire N__24512;
    wire N__24511;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24427;
    wire N__24424;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24376;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24341;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24329;
    wire N__24326;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24318;
    wire N__24317;
    wire N__24316;
    wire N__24315;
    wire N__24314;
    wire N__24313;
    wire N__24312;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24298;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24253;
    wire N__24250;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24235;
    wire N__24234;
    wire N__24233;
    wire N__24232;
    wire N__24231;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24209;
    wire N__24202;
    wire N__24197;
    wire N__24194;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24161;
    wire N__24154;
    wire N__24153;
    wire N__24150;
    wire N__24149;
    wire N__24148;
    wire N__24145;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24094;
    wire N__24091;
    wire N__24082;
    wire N__24065;
    wire N__24064;
    wire N__24061;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24043;
    wire N__24042;
    wire N__24039;
    wire N__24034;
    wire N__24031;
    wire N__24030;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24015;
    wire N__24014;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23991;
    wire N__23988;
    wire N__23983;
    wire N__23980;
    wire N__23975;
    wire N__23974;
    wire N__23973;
    wire N__23972;
    wire N__23969;
    wire N__23964;
    wire N__23961;
    wire N__23954;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23940;
    wire N__23939;
    wire N__23938;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23922;
    wire N__23921;
    wire N__23920;
    wire N__23919;
    wire N__23918;
    wire N__23917;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23868;
    wire N__23863;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23779;
    wire N__23776;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23750;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23707;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23617;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23569;
    wire N__23568;
    wire N__23567;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23559;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23544;
    wire N__23539;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23524;
    wire N__23523;
    wire N__23520;
    wire N__23513;
    wire N__23508;
    wire N__23501;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23493;
    wire N__23490;
    wire N__23489;
    wire N__23488;
    wire N__23487;
    wire N__23486;
    wire N__23485;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23469;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23457;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23409;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23338;
    wire N__23337;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23316;
    wire N__23313;
    wire N__23308;
    wire N__23305;
    wire N__23300;
    wire N__23299;
    wire N__23294;
    wire N__23291;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23279;
    wire N__23278;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23192;
    wire N__23189;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23144;
    wire N__23143;
    wire N__23142;
    wire N__23141;
    wire N__23138;
    wire N__23137;
    wire N__23134;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23118;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23093;
    wire N__23090;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23053;
    wire N__23052;
    wire N__23049;
    wire N__23044;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22898;
    wire N__22895;
    wire N__22894;
    wire N__22893;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22840;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22729;
    wire N__22726;
    wire N__22725;
    wire N__22724;
    wire N__22723;
    wire N__22722;
    wire N__22721;
    wire N__22720;
    wire N__22719;
    wire N__22716;
    wire N__22715;
    wire N__22712;
    wire N__22707;
    wire N__22700;
    wire N__22699;
    wire N__22698;
    wire N__22697;
    wire N__22696;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22688;
    wire N__22687;
    wire N__22686;
    wire N__22685;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22677;
    wire N__22676;
    wire N__22675;
    wire N__22674;
    wire N__22669;
    wire N__22666;
    wire N__22657;
    wire N__22654;
    wire N__22645;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22623;
    wire N__22618;
    wire N__22601;
    wire N__22600;
    wire N__22599;
    wire N__22598;
    wire N__22597;
    wire N__22596;
    wire N__22595;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22584;
    wire N__22583;
    wire N__22582;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22574;
    wire N__22573;
    wire N__22570;
    wire N__22569;
    wire N__22566;
    wire N__22559;
    wire N__22556;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22537;
    wire N__22530;
    wire N__22527;
    wire N__22526;
    wire N__22525;
    wire N__22520;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22494;
    wire N__22493;
    wire N__22492;
    wire N__22489;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22468;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22442;
    wire N__22441;
    wire N__22440;
    wire N__22439;
    wire N__22438;
    wire N__22437;
    wire N__22436;
    wire N__22433;
    wire N__22432;
    wire N__22431;
    wire N__22430;
    wire N__22423;
    wire N__22420;
    wire N__22419;
    wire N__22410;
    wire N__22409;
    wire N__22408;
    wire N__22407;
    wire N__22406;
    wire N__22405;
    wire N__22404;
    wire N__22403;
    wire N__22402;
    wire N__22397;
    wire N__22392;
    wire N__22389;
    wire N__22388;
    wire N__22387;
    wire N__22386;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22366;
    wire N__22361;
    wire N__22354;
    wire N__22345;
    wire N__22342;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22322;
    wire N__22321;
    wire N__22320;
    wire N__22319;
    wire N__22316;
    wire N__22307;
    wire N__22300;
    wire N__22299;
    wire N__22298;
    wire N__22297;
    wire N__22296;
    wire N__22295;
    wire N__22294;
    wire N__22293;
    wire N__22292;
    wire N__22291;
    wire N__22286;
    wire N__22285;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22277;
    wire N__22276;
    wire N__22275;
    wire N__22274;
    wire N__22267;
    wire N__22258;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22241;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22204;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22138;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22107;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22072;
    wire N__22069;
    wire N__22068;
    wire N__22067;
    wire N__22066;
    wire N__22065;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22057;
    wire N__22054;
    wire N__22049;
    wire N__22048;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22022;
    wire N__22019;
    wire N__22014;
    wire N__22007;
    wire N__22004;
    wire N__22003;
    wire N__22002;
    wire N__21997;
    wire N__21992;
    wire N__21987;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21888;
    wire N__21887;
    wire N__21884;
    wire N__21883;
    wire N__21880;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21860;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21787;
    wire N__21786;
    wire N__21785;
    wire N__21784;
    wire N__21781;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21766;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21754;
    wire N__21749;
    wire N__21746;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21728;
    wire N__21725;
    wire N__21724;
    wire N__21723;
    wire N__21722;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21700;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21688;
    wire N__21683;
    wire N__21674;
    wire N__21671;
    wire N__21670;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21564;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21546;
    wire N__21539;
    wire N__21536;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21487;
    wire N__21486;
    wire N__21485;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21471;
    wire N__21470;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21431;
    wire N__21428;
    wire N__21421;
    wire N__21416;
    wire N__21413;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21313;
    wire N__21312;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21277;
    wire N__21274;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21235;
    wire N__21234;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21095;
    wire N__21094;
    wire N__21093;
    wire N__21090;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21057;
    wire N__21054;
    wire N__21049;
    wire N__21044;
    wire N__21041;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20971;
    wire N__20970;
    wire N__20967;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20950;
    wire N__20945;
    wire N__20944;
    wire N__20941;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20926;
    wire N__20921;
    wire N__20918;
    wire N__20917;
    wire N__20916;
    wire N__20915;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20895;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20873;
    wire N__20870;
    wire N__20869;
    wire N__20868;
    wire N__20867;
    wire N__20866;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20833;
    wire N__20830;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20767;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20701;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20668;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20587;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20572;
    wire N__20567;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20555;
    wire N__20554;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20542;
    wire N__20541;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20483;
    wire N__20480;
    wire N__20479;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20462;
    wire N__20459;
    wire N__20458;
    wire N__20457;
    wire N__20456;
    wire N__20455;
    wire N__20454;
    wire N__20453;
    wire N__20450;
    wire N__20445;
    wire N__20436;
    wire N__20435;
    wire N__20428;
    wire N__20425;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20365;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20329;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20302;
    wire N__20301;
    wire N__20294;
    wire N__20291;
    wire N__20290;
    wire N__20289;
    wire N__20286;
    wire N__20281;
    wire N__20278;
    wire N__20277;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20089;
    wire N__20088;
    wire N__20087;
    wire N__20084;
    wire N__20083;
    wire N__20082;
    wire N__20069;
    wire N__20066;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20041;
    wire N__20040;
    wire N__20037;
    wire N__20032;
    wire N__20027;
    wire N__20024;
    wire N__20023;
    wire N__20022;
    wire N__20015;
    wire N__20014;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19981;
    wire N__19980;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19930;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19853;
    wire N__19850;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19842;
    wire N__19839;
    wire N__19838;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19820;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19789;
    wire N__19788;
    wire N__19785;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19767;
    wire N__19764;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19733;
    wire N__19732;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19696;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19677;
    wire N__19672;
    wire N__19669;
    wire N__19664;
    wire N__19661;
    wire N__19660;
    wire N__19655;
    wire N__19652;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19640;
    wire N__19639;
    wire N__19634;
    wire N__19631;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19585;
    wire N__19580;
    wire N__19577;
    wire N__19576;
    wire N__19575;
    wire N__19572;
    wire N__19567;
    wire N__19562;
    wire N__19559;
    wire N__19558;
    wire N__19557;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19540;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19522;
    wire N__19519;
    wire N__19514;
    wire N__19511;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19405;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19270;
    wire N__19269;
    wire N__19266;
    wire N__19261;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19225;
    wire N__19220;
    wire N__19217;
    wire N__19216;
    wire N__19215;
    wire N__19212;
    wire N__19207;
    wire N__19204;
    wire N__19199;
    wire N__19198;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19172;
    wire N__19171;
    wire N__19170;
    wire N__19169;
    wire N__19164;
    wire N__19159;
    wire N__19156;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19144;
    wire N__19141;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19102;
    wire N__19099;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19091;
    wire N__19090;
    wire N__19089;
    wire N__19086;
    wire N__19085;
    wire N__19082;
    wire N__19081;
    wire N__19080;
    wire N__19077;
    wire N__19074;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19055;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19003;
    wire N__19002;
    wire N__18997;
    wire N__18994;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18972;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18952;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18940;
    wire N__18939;
    wire N__18936;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18835;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18794;
    wire N__18791;
    wire N__18790;
    wire N__18785;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18775;
    wire N__18772;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18739;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18731;
    wire N__18730;
    wire N__18729;
    wire N__18728;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18717;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18703;
    wire N__18698;
    wire N__18695;
    wire N__18690;
    wire N__18685;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18669;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18648;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18632;
    wire N__18629;
    wire N__18628;
    wire N__18627;
    wire N__18624;
    wire N__18619;
    wire N__18618;
    wire N__18615;
    wire N__18614;
    wire N__18609;
    wire N__18600;
    wire N__18597;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18550;
    wire N__18549;
    wire N__18546;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18530;
    wire N__18527;
    wire N__18526;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18502;
    wire N__18497;
    wire N__18494;
    wire N__18489;
    wire N__18482;
    wire N__18481;
    wire N__18476;
    wire N__18475;
    wire N__18474;
    wire N__18471;
    wire N__18466;
    wire N__18463;
    wire N__18458;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18419;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18347;
    wire N__18344;
    wire N__18343;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18316;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18245;
    wire N__18242;
    wire N__18241;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18151;
    wire N__18146;
    wire N__18143;
    wire N__18142;
    wire N__18141;
    wire N__18140;
    wire N__18139;
    wire N__18138;
    wire N__18127;
    wire N__18124;
    wire N__18123;
    wire N__18122;
    wire N__18121;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18105;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18091;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18079;
    wire N__18074;
    wire N__18065;
    wire N__18062;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18054;
    wire N__18053;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18039;
    wire N__18034;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18022;
    wire N__18019;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17938;
    wire N__17937;
    wire N__17930;
    wire N__17927;
    wire N__17926;
    wire N__17925;
    wire N__17924;
    wire N__17923;
    wire N__17922;
    wire N__17921;
    wire N__17918;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17897;
    wire N__17888;
    wire N__17885;
    wire N__17884;
    wire N__17883;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17862;
    wire N__17855;
    wire N__17854;
    wire N__17853;
    wire N__17852;
    wire N__17849;
    wire N__17848;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17840;
    wire N__17839;
    wire N__17836;
    wire N__17823;
    wire N__17820;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17808;
    wire N__17803;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17764;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17746;
    wire N__17745;
    wire N__17744;
    wire N__17743;
    wire N__17740;
    wire N__17731;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17716;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17647;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17590;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17575;
    wire N__17570;
    wire N__17567;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17555;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17533;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17492;
    wire N__17491;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17461;
    wire N__17456;
    wire N__17455;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17354;
    wire N__17353;
    wire N__17348;
    wire N__17345;
    wire N__17344;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17299;
    wire N__17296;
    wire N__17295;
    wire N__17294;
    wire N__17291;
    wire N__17284;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17251;
    wire N__17250;
    wire N__17247;
    wire N__17244;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17228;
    wire N__17225;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17214;
    wire N__17213;
    wire N__17212;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17198;
    wire N__17195;
    wire N__17186;
    wire N__17185;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17170;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17137;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17125;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17098;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17027;
    wire N__17024;
    wire N__17023;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16996;
    wire N__16993;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16981;
    wire N__16980;
    wire N__16977;
    wire N__16972;
    wire N__16967;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16952;
    wire N__16949;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16931;
    wire N__16928;
    wire N__16927;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16864;
    wire N__16863;
    wire N__16860;
    wire N__16855;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16843;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16768;
    wire N__16763;
    wire N__16760;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16742;
    wire N__16741;
    wire N__16736;
    wire N__16733;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16725;
    wire N__16722;
    wire N__16717;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16687;
    wire N__16686;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16674;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16618;
    wire N__16617;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16603;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16591;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16574;
    wire N__16573;
    wire N__16572;
    wire N__16567;
    wire N__16564;
    wire N__16559;
    wire N__16556;
    wire N__16555;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16499;
    wire N__16496;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16450;
    wire N__16449;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16430;
    wire N__16427;
    wire N__16426;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16399;
    wire N__16394;
    wire N__16393;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16369;
    wire N__16368;
    wire N__16365;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16349;
    wire N__16346;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16313;
    wire N__16312;
    wire N__16309;
    wire N__16308;
    wire N__16307;
    wire N__16304;
    wire N__16301;
    wire N__16296;
    wire N__16293;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16279;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16240;
    wire N__16235;
    wire N__16232;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16189;
    wire N__16186;
    wire N__16185;
    wire N__16182;
    wire N__16181;
    wire N__16178;
    wire N__16171;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16157;
    wire N__16156;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16121;
    wire N__16120;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16102;
    wire N__16101;
    wire N__16098;
    wire N__16093;
    wire N__16090;
    wire N__16085;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16052;
    wire N__16051;
    wire N__16050;
    wire N__16049;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16031;
    wire N__16028;
    wire N__16027;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15988;
    wire N__15985;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15925;
    wire N__15922;
    wire N__15921;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15902;
    wire N__15901;
    wire N__15898;
    wire N__15897;
    wire N__15896;
    wire N__15893;
    wire N__15892;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15870;
    wire N__15863;
    wire N__15862;
    wire N__15861;
    wire N__15858;
    wire N__15857;
    wire N__15854;
    wire N__15851;
    wire N__15850;
    wire N__15847;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15818;
    wire N__15815;
    wire N__15814;
    wire N__15813;
    wire N__15812;
    wire N__15811;
    wire N__15806;
    wire N__15803;
    wire N__15798;
    wire N__15795;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15766;
    wire N__15763;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15575;
    wire N__15572;
    wire N__15571;
    wire N__15570;
    wire N__15567;
    wire N__15562;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15478;
    wire N__15477;
    wire N__15476;
    wire N__15473;
    wire N__15468;
    wire N__15463;
    wire N__15460;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15445;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15361;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15280;
    wire N__15277;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15250;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15226;
    wire N__15225;
    wire N__15224;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15205;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15184;
    wire N__15181;
    wire N__15176;
    wire N__15173;
    wire GNDG0;
    wire VCCG0;
    wire \INVFTDI.RXbuffer_3C_net ;
    wire \INVFTDI.RXbuffer_0C_net ;
    wire ctrlOut_8;
    wire \ALU.m289_nsZ0Z_1_cascade_ ;
    wire ctrlOut_5;
    wire \ALU.N_223_0_cascade_ ;
    wire \ALU.a9_b_3_cascade_ ;
    wire \ALU.a7_b_5 ;
    wire \ALU.a9_b_3 ;
    wire \ALU.g0_0_a3_2_0_cascade_ ;
    wire \ALU.madd_315_0_cascade_ ;
    wire \ALU.a12_b_1 ;
    wire \ALU.madd_315_0 ;
    wire \ALU.a12_b_1_cascade_ ;
    wire \ALU.madd_264 ;
    wire \ALU.madd_141_0_cascade_ ;
    wire \ALU.N_1545_0 ;
    wire \ALU.madd_166_0 ;
    wire \ALU.madd_254_0_tz_cascade_ ;
    wire \ALU.madd_141 ;
    wire \ALU.madd_254_cascade_ ;
    wire \ALU.madd_254_0_tz ;
    wire \ALU.m292_nsZ0Z_1 ;
    wire \ALU.N_90_0_cascade_ ;
    wire ctrlOut_6;
    wire \ALU.N_217_0_cascade_ ;
    wire \ALU.un9_addsub_axb_10_cascade_ ;
    wire \ALU.a3_b_0_10_cascade_ ;
    wire \ALU.g0_2_cascade_ ;
    wire \ALU.N_1555_0 ;
    wire \ALU.N_1527_0 ;
    wire \ALU.madd_171_cascade_ ;
    wire \ALU.madd_161_0_cascade_ ;
    wire \ALU.madd_161 ;
    wire \ALU.madd_166 ;
    wire \ALU.madd_171 ;
    wire \ALU.madd_161_cascade_ ;
    wire \ALU.a8_b_3_cascade_ ;
    wire \ALU.a8_b_3 ;
    wire \ALU.g0_0_2 ;
    wire \ALU.g0_0_cascade_ ;
    wire \ALU.N_1527_1_0 ;
    wire \ALU.g2_0_1 ;
    wire \ALU.g1 ;
    wire \ALU.g0_1_0 ;
    wire \ALU.madd_124_0_cascade_ ;
    wire \ALU.madd_124_cascade_ ;
    wire \ALU.madd_144_cascade_ ;
    wire \ALU.madd_324_cascade_ ;
    wire \ALU.madd_N_9_cascade_ ;
    wire \ALU.madd_191_0 ;
    wire \ALU.madd_186 ;
    wire \ALU.madd_191_0_cascade_ ;
    wire \ALU.madd_324 ;
    wire \ALU.madd_326_cascade_ ;
    wire \ALU.madd_325 ;
    wire clkdivZ0Z_0;
    wire bfn_1_16_0_;
    wire clkdivZ0Z_1;
    wire clkdiv_cry_0;
    wire clkdivZ0Z_2;
    wire clkdiv_cry_1;
    wire clkdivZ0Z_3;
    wire clkdiv_cry_2;
    wire clkdivZ0Z_4;
    wire clkdiv_cry_3;
    wire clkdivZ0Z_5;
    wire clkdiv_cry_4;
    wire clkdivZ0Z_6;
    wire clkdiv_cry_5;
    wire clkdivZ0Z_7;
    wire clkdiv_cry_6;
    wire clkdiv_cry_7;
    wire clkdivZ0Z_8;
    wire bfn_1_17_0_;
    wire clkdivZ0Z_9;
    wire clkdiv_cry_8;
    wire clkdivZ0Z_10;
    wire clkdiv_cry_9;
    wire clkdivZ0Z_11;
    wire clkdiv_cry_10;
    wire clkdivZ0Z_12;
    wire clkdiv_cry_11;
    wire clkdivZ0Z_13;
    wire clkdiv_cry_12;
    wire clkdivZ0Z_14;
    wire clkdiv_cry_13;
    wire clkdivZ0Z_15;
    wire clkdiv_cry_14;
    wire clkdiv_cry_15;
    wire clkdivZ0Z_16;
    wire bfn_1_18_0_;
    wire clkdivZ0Z_17;
    wire clkdiv_cry_16;
    wire clkdivZ0Z_18;
    wire clkdiv_cry_17;
    wire clkdivZ0Z_19;
    wire clkdiv_cry_18;
    wire clkdivZ0Z_20;
    wire clkdiv_cry_19;
    wire clkdivZ0Z_21;
    wire clkdiv_cry_20;
    wire clkdivZ0Z_22;
    wire clkdiv_cry_21;
    wire clkdiv_cry_22;
    wire GPIO3_c;
    wire testWordZ0Z_13;
    wire \ALU.m304_nsZ0Z_1_cascade_ ;
    wire \ALU.i73_mux_1_cascade_ ;
    wire RXbuffer_0;
    wire RXbuffer_7;
    wire RXbuffer_1;
    wire RXbuffer_3;
    wire N_661_0_cascade_;
    wire \ALU.un2_addsub_axb_8_cascade_ ;
    wire \ALU.N_275_0_cascade_ ;
    wire \ALU.g0_0_0_N_3L3 ;
    wire \ALU.g0_0_0_N_4L5_cascade_ ;
    wire \ALU.g0_0_0_N_3L3_0 ;
    wire \ALU.a5_b_9_cascade_ ;
    wire \ALU.operand2_8_cascade_ ;
    wire \ALU.a1_b_8 ;
    wire \ALU.a1_b_8_cascade_ ;
    wire \ALU.a4_b_8_cascade_ ;
    wire \ALU.madd_269 ;
    wire \ALU.madd_i1_mux_cascade_ ;
    wire \ALU.g0_14 ;
    wire \ALU.madd_i3_mux_cascade_ ;
    wire \ALU.madd_331_cascade_ ;
    wire \ALU.madd_328 ;
    wire \ALU.madd_340_0 ;
    wire \ALU.g0_1_cascade_ ;
    wire \ALU.g2 ;
    wire \ALU.N_1545_1 ;
    wire \ALU.g0_3_cascade_ ;
    wire \ALU.madd_350_0 ;
    wire \ALU.madd_350_0_cascade_ ;
    wire \ALU.madd_335 ;
    wire \ALU.madd_i1_mux_2 ;
    wire \ALU.madd_289 ;
    wire \ALU.madd_227 ;
    wire \ALU.madd_227_cascade_ ;
    wire \ALU.madd_165_0_0_cascade_ ;
    wire \ALU.madd_170_0_tz_cascade_ ;
    wire \ALU.madd_90 ;
    wire \ALU.madd_223_0_cascade_ ;
    wire \ALU.N_1533_0 ;
    wire \ALU.N_1559_0 ;
    wire \ALU.madd_165_0_tz ;
    wire \ALU.madd_165_0 ;
    wire \ALU.a5_b_5 ;
    wire \ALU.a5_b_5_cascade_ ;
    wire \ALU.a4_b_6 ;
    wire \ALU.madd_175_cascade_ ;
    wire \ALU.madd_232 ;
    wire \ALU.madd_175 ;
    wire \ALU.madd_213_0 ;
    wire \ALU.a7_b_4_cascade_ ;
    wire \ALU.madd_208 ;
    wire \ALU.N_225_0_cascade_ ;
    wire \ALU.madd_290_0_cascade_ ;
    wire \ALU.madd_299_cascade_ ;
    wire \ALU.g0_11 ;
    wire \ALU.madd_299 ;
    wire \ALU.madd_223_0 ;
    wire \ALU.madd_228 ;
    wire \ALU.madd_170 ;
    wire \ALU.madd_265_0_cascade_ ;
    wire \ALU.madd_280 ;
    wire \ALU.madd_280_cascade_ ;
    wire \ALU.madd_285 ;
    wire \ALU.madd_326 ;
    wire \ALU.a4_b_7 ;
    wire \ALU.a4_b_7_cascade_ ;
    wire \ALU.madd_233_cascade_ ;
    wire \ALU.madd_237 ;
    wire \ALU.madd_242 ;
    wire \ALU.madd_247_cascade_ ;
    wire \ALU.madd_295_0 ;
    wire \ALU.madd_N_10 ;
    wire \ALU.madd_247 ;
    wire \ALU.madd_N_10_cascade_ ;
    wire \ALU.madd_N_5_0 ;
    wire \ALU.madd_190 ;
    wire \ALU.madd_238_0 ;
    wire \ALU.madd_233 ;
    wire \ALU.madd_327 ;
    wire \ALU.un2_addsub_axb_7_cascade_ ;
    wire \ALU.a0_b_8_cascade_ ;
    wire \ALU.madd_103 ;
    wire \ALU.madd_124 ;
    wire \ALU.madd_148 ;
    wire \ALU.madd_148_cascade_ ;
    wire \ALU.madd_247_0_tz_0 ;
    wire \ALU.madd_143 ;
    wire \ALU.madd_181 ;
    wire \ALU.madd_129 ;
    wire \ALU.a5_b_4 ;
    wire \ALU.a5_b_4_cascade_ ;
    wire \ALU.madd_133_cascade_ ;
    wire \ALU.madd_237_0_tz_0 ;
    wire \ALU.madd_133 ;
    wire \ALU.madd_138 ;
    wire \ALU.madd_128_0_0_0_cascade_ ;
    wire \ALU.madd_70 ;
    wire \ALU.madd_237_0_tz_0_1_cascade_ ;
    wire \ALU.g0_0_0 ;
    wire \ALU.N_1537_0_0_1 ;
    wire \ALU.i6_mux_cascade_ ;
    wire N_51_0_cascade_;
    wire testWordZ0Z_15;
    wire N_662_0_cascade_;
    wire N_665_0;
    wire N_301_0_cascade_;
    wire N_668_0_cascade_;
    wire \ALU.m300_nsZ0Z_1 ;
    wire N_662_0;
    wire N_670_0_cascade_;
    wire \CONTROL.results_cnvZ0Z_0 ;
    wire \ALU.un2_addsub_axb_14 ;
    wire \ALU.un2_addsub_axb_9_cascade_ ;
    wire \ALU.a13_b_1_cascade_ ;
    wire \ALU.a11_b_3 ;
    wire \ALU.a11_b_3_cascade_ ;
    wire ctrlOut_14;
    wire RXbuffer_6;
    wire testWordZ0Z_14;
    wire \ALU.a7_b_6_cascade_ ;
    wire \ALU.a6_b_7 ;
    wire \ALU.a7_b_6 ;
    wire \ALU.madd_324_0 ;
    wire \ALU.madd_324_0_cascade_ ;
    wire \ALU.madd_372 ;
    wire \ALU.madd_396 ;
    wire \ALU.madd_484_21 ;
    wire \ALU.madd_411_cascade_ ;
    wire \ALU.madd_484_24 ;
    wire \ALU.a8_b_6 ;
    wire \ALU.a9_b_5 ;
    wire \ALU.madd_377 ;
    wire \ALU.madd_372_0 ;
    wire \ALU.madd_382 ;
    wire \ALU.madd_377_cascade_ ;
    wire \ALU.a13_b_1 ;
    wire \ALU.madd_397 ;
    wire \ALU.madd_392 ;
    wire \ALU.madd_397_cascade_ ;
    wire \ALU.madd_339 ;
    wire \ALU.madd_406 ;
    wire \ALU.a5_b_8_cascade_ ;
    wire \ALU.madd_387 ;
    wire \ALU.madd_329_0 ;
    wire \ALU.madd_387_cascade_ ;
    wire \ALU.madd_402 ;
    wire \ALU.madd_402_cascade_ ;
    wire \ALU.madd_354 ;
    wire \ALU.madd_412_cascade_ ;
    wire \ALU.madd_329 ;
    wire \ALU.madd_407 ;
    wire \ALU.madd_412 ;
    wire \ALU.madd_i3_mux_1 ;
    wire \ALU.madd_330 ;
    wire \ALU.madd_141_1 ;
    wire \ALU.madd_270_0 ;
    wire \ALU.madd_250_0 ;
    wire \ALU.madd_250_0_cascade_ ;
    wire \ALU.madd_250 ;
    wire \ALU.a3_b_9 ;
    wire \ALU.madd_250_cascade_ ;
    wire \ALU.madd_207 ;
    wire \ALU.madd_274 ;
    wire \ALU.madd_320 ;
    wire \ALU.madd_325_0 ;
    wire \ALU.madd_274_cascade_ ;
    wire \ALU.madd_254 ;
    wire \ALU.madd_344 ;
    wire \ALU.madd_29_cascade_ ;
    wire \ALU.madd_47_cascade_ ;
    wire \ALU.madd_265_0 ;
    wire \ALU.madd_260 ;
    wire \ALU.a2_b_6 ;
    wire \ALU.a0_b_8 ;
    wire \ALU.a2_b_6_cascade_ ;
    wire \ALU.a5_b_6_cascade_ ;
    wire \ALU.operand2_5_cascade_ ;
    wire \ALU.madd_176_0 ;
    wire \ALU.madd_218_0 ;
    wire \ALU.a7_b_4 ;
    wire \ALU.a6_b_5 ;
    wire \ALU.a5_b_6 ;
    wire \ALU.madd_275_0 ;
    wire \ALU.madd_42_cascade_ ;
    wire \ALU.madd_42_0 ;
    wire \ALU.e_RNIM09HZ0Z_7_cascade_ ;
    wire \ALU.operand2_7_ns_1_7_cascade_ ;
    wire \ALU.g1_2_cascade_ ;
    wire \ALU.a4_b_0_7 ;
    wire \ALU.g2_0_0_0 ;
    wire \ALU.un2_addsub_axb_5_cascade_ ;
    wire \ALU.a6_b_0_7 ;
    wire \ALU.a6_b_0_cascade_ ;
    wire \ALU.madd_41_cascade_ ;
    wire \ALU.madd_46_cascade_ ;
    wire \ALU.madd_39_cascade_ ;
    wire \ALU.a6_b_3 ;
    wire \ALU.madd_78_0_tz_cascade_ ;
    wire \ALU.madd_78_0 ;
    wire \ALU.madd_39 ;
    wire \ALU.madd_78_0_cascade_ ;
    wire \ALU.madd_114_cascade_ ;
    wire testClock_0_cascade_;
    wire \ALU.a_cnv_0Z0Z_0_cascade_ ;
    wire \ALU.N_53_0 ;
    wire aluResults_0;
    wire testClock_0;
    wire testClockZ0;
    wire \ALU.a_cnv_0Z0Z_0 ;
    wire aluResults_1;
    wire \ALU.b_cnv_0Z0Z_0 ;
    wire aluResults_2;
    wire \ALU.N_169_0 ;
    wire \ALU.c_RNIEP354Z0Z_14_cascade_ ;
    wire \ALU.c_RNIJENJ8_0Z0Z_15 ;
    wire \ALU.rshift_3_ns_1_6_cascade_ ;
    wire \ALU.N_474_cascade_ ;
    wire \ALU.rshift_15_ns_1_6 ;
    wire \ALU.rshift_6_cascade_ ;
    wire \ALU.N_291_0 ;
    wire \ALU.dout_6_ns_1_14_cascade_ ;
    wire \ALU.aluOut_15_cascade_ ;
    wire \ALU.N_761 ;
    wire \ALU.N_713 ;
    wire \ALU.a_15_m2_ns_1Z0Z_14_cascade_ ;
    wire \ALU.lshift_15_ns_1_14_cascade_ ;
    wire \ALU.lshift_14_cascade_ ;
    wire \ALU.a_15_m2_14 ;
    wire \ALU.a_15_m4_14_cascade_ ;
    wire \ALU.a_15_m3_14 ;
    wire \ALU.dout_3_ns_1_12_cascade_ ;
    wire \ALU.dout_6_ns_1_12_cascade_ ;
    wire \ALU.N_711 ;
    wire \ALU.N_759_cascade_ ;
    wire \ALU.aluOut_12_cascade_ ;
    wire \ALU.a12_b_2 ;
    wire \ALU.N_90_0 ;
    wire ctrlOut_3;
    wire \ALU.N_235_0_cascade_ ;
    wire \ALU.a12_b_3_cascade_ ;
    wire ctrlOut_4;
    wire \ALU.a9_b_4 ;
    wire \ALU.a10_b_3_cascade_ ;
    wire \ALU.madd_319 ;
    wire \ALU.madd_366 ;
    wire \ALU.madd_484_11 ;
    wire \ALU.madd_376 ;
    wire \ALU.madd_484_17_cascade_ ;
    wire \ALU.madd_484_15 ;
    wire \ALU.madd_484_20 ;
    wire \ALU.madd_309 ;
    wire \ALU.madd_362 ;
    wire \ALU.madd_391 ;
    wire \ALU.a5_b_9 ;
    wire \ALU.a6_b_8 ;
    wire \ALU.a7_b_7_cascade_ ;
    wire \ALU.madd_381 ;
    wire \ALU.madd_484_16 ;
    wire \ALU.un9_addsub_axb_12_cascade_ ;
    wire \ALU.d_RNIV96U8Z0Z_13_cascade_ ;
    wire \ALU.madd_314 ;
    wire \ALU.madd_310_0_cascade_ ;
    wire \ALU.madd_334 ;
    wire \ALU.a1_b_12 ;
    wire \ALU.a2_b_9_cascade_ ;
    wire \ALU.operand2_8 ;
    wire \ALU.N_199_0 ;
    wire \ALU.a3_b_8 ;
    wire \ALU.madd_275 ;
    wire \ALU.madd_217 ;
    wire \ALU.madd_222 ;
    wire \ALU.madd_212 ;
    wire \ALU.madd_284 ;
    wire \ALU.madd_279_cascade_ ;
    wire \ALU.madd_349 ;
    wire \ALU.d_RNIV96U8Z0Z_13 ;
    wire \ALU.madd_310_0 ;
    wire \ALU.madd_330_0 ;
    wire \ALU.c_RNIF549Z0Z_10_cascade_ ;
    wire \ALU.a_RNIBLBOZ0Z_10 ;
    wire \ALU.operand2_7_ns_1_10_cascade_ ;
    wire \ALU.operand2_10_cascade_ ;
    wire \ALU.a4_b_10 ;
    wire \ALU.a3_b_10 ;
    wire \ALU.a3_b_10_cascade_ ;
    wire \ALU.madd_305 ;
    wire \ALU.madd_5_cascade_ ;
    wire \ALU.madd_19 ;
    wire \ALU.madd_17 ;
    wire \ALU.madd_19_cascade_ ;
    wire \ALU.madd_47 ;
    wire \ALU.g0_0_a3_0 ;
    wire \ALU.a8_b_0_cascade_ ;
    wire \ALU.madd_10_cascade_ ;
    wire \ALU.madd_24 ;
    wire \ALU.madd_29 ;
    wire \ALU.madd_24_cascade_ ;
    wire \ALU.madd_i1_mux_1 ;
    wire \ALU.madd_i3_mux_0 ;
    wire \ALU.a4_b_2 ;
    wire \ALU.a6_b_0 ;
    wire \ALU.madd_12_cascade_ ;
    wire \ALU.madd_34 ;
    wire \ALU.madd_42 ;
    wire \ALU.madd_34_cascade_ ;
    wire \ALU.madd_37 ;
    wire \ALU.madd_56_cascade_ ;
    wire \ALU.madd_52_0 ;
    wire \ALU.madd_25 ;
    wire \ALU.madd_12 ;
    wire \ALU.un2_addsub_axb_6_cascade_ ;
    wire \ALU.madd_64_0 ;
    wire \ALU.madd_74_0_cascade_ ;
    wire \ALU.madd_83 ;
    wire \ALU.madd_46 ;
    wire \ALU.madd_69 ;
    wire \ALU.madd_74_0 ;
    wire \ALU.madd_79_0 ;
    wire \ALU.madd_51 ;
    wire \ALU.madd_58 ;
    wire \ALU.madd_79_0_cascade_ ;
    wire \ALU.madd_56 ;
    wire \ALU.madd_88_cascade_ ;
    wire \ALU.madd_114 ;
    wire \ALU.madd_41 ;
    wire \ALU.madd_73_cascade_ ;
    wire \ALU.operand2_7 ;
    wire \ALU.a0_b_7 ;
    wire \ALU.madd_144 ;
    wire \ALU.madd_113 ;
    wire \ALU.madd_154_cascade_ ;
    wire \ALU.madd_99 ;
    wire \ALU.madd_73 ;
    wire \ALU.madd_109 ;
    wire \ALU.madd_154 ;
    wire \ALU.madd_118 ;
    wire \ALU.m641_nsZ0Z_1 ;
    wire \ALU.m645_nsZ0Z_1 ;
    wire \ALU.N_283_0_cascade_ ;
    wire \ALU.m55_bmZ0 ;
    wire \ALU.m55_amZ0 ;
    wire \ALU.m650_nsZ0Z_1_cascade_ ;
    wire \ALU.N_15_0 ;
    wire N_727;
    wire \ALU.N_577_cascade_ ;
    wire \ALU.N_528_cascade_ ;
    wire \ALU.N_633 ;
    wire \ALU.d_RNI8DL9U1Z0Z_3_cascade_ ;
    wire \ALU.N_221_cascade_ ;
    wire \ALU.N_588_cascade_ ;
    wire \ALU.N_575 ;
    wire \ALU.N_575_cascade_ ;
    wire \ALU.rshift_3_ns_1_8 ;
    wire \ALU.lshift_3_ns_1_15 ;
    wire \ALU.dout_3_ns_1_14 ;
    wire \ALU.lshift_3_ns_1_14_cascade_ ;
    wire \ALU.N_256 ;
    wire \ALU.N_224_cascade_ ;
    wire \ALU.N_220_cascade_ ;
    wire \ALU.N_222 ;
    wire \ALU.madd_484_4 ;
    wire \ALU.N_241_0 ;
    wire \ALU.N_240_0_i_cascade_ ;
    wire \ALU.N_9_0 ;
    wire \ALU.N_10_0 ;
    wire \ALU.N_253_0 ;
    wire \ALU.d_RNIUV3H4Z0Z_0 ;
    wire \ALU.N_635_0 ;
    wire \ALU.N_724 ;
    wire \ALU.N_283_0 ;
    wire ctrlOut_7;
    wire \ALU.N_211_0 ;
    wire ctrlOut_9;
    wire \ALU.madd_367 ;
    wire \ALU.d_RNIRV558Z0Z_13 ;
    wire \ALU.d_RNIRV558Z0Z_13_cascade_ ;
    wire \ALU.madd_371 ;
    wire \ALU.a2_b_12 ;
    wire \ALU.madd_259 ;
    wire \ALU.N_186_0_cascade_ ;
    wire \ALU.a1_b_11 ;
    wire \ALU.a0_b_12 ;
    wire \ALU.a1_b_11_cascade_ ;
    wire \ALU.madd_255 ;
    wire \ALU.dout_6_ns_1_8_cascade_ ;
    wire \ALU.dout_3_ns_1_8 ;
    wire \ALU.N_707_cascade_ ;
    wire \ALU.N_755 ;
    wire \ALU.m272_nsZ0Z_1_cascade_ ;
    wire \ALU.N_191_0_0 ;
    wire ctrlOut_10;
    wire \ALU.N_191_0 ;
    wire \ALU.N_191_0_cascade_ ;
    wire \ALU.operand2_10 ;
    wire \ALU.a1_b_10 ;
    wire \ALU.a1_b_10_cascade_ ;
    wire \ALU.madd_203 ;
    wire \ALU.a9_b_2 ;
    wire \ALU.dout_3_ns_1_9_cascade_ ;
    wire \ALU.N_708_cascade_ ;
    wire \ALU.dout_6_ns_1_9_cascade_ ;
    wire \ALU.N_756 ;
    wire \ALU.N_751_cascade_ ;
    wire \ALU.N_703 ;
    wire \ALU.rshift_3_ns_1_4_cascade_ ;
    wire \ALU.N_472 ;
    wire \ALU.N_472_cascade_ ;
    wire \ALU.N_476 ;
    wire \ALU.N_706_cascade_ ;
    wire \ALU.N_754 ;
    wire \ALU.aluOut_7_cascade_ ;
    wire \ALU.a7_b_0_6 ;
    wire \ALU.m271_nsZ0Z_1 ;
    wire \ALU.madd_20_0_cascade_ ;
    wire \ALU.madd_20 ;
    wire ctrlOut_2;
    wire \ALU.N_5_0_cascade_ ;
    wire \ALU.N_240_0_cascade_ ;
    wire \ALU.madd_24_0_tz ;
    wire \ALU.madd_8_0 ;
    wire \ALU.madd_5 ;
    wire \ALU.madd_8_0_cascade_ ;
    wire \ALU.a7_b_0_cascade_ ;
    wire \ALU.madd_59 ;
    wire \ALU.madd_484_5 ;
    wire \ALU.madd_128_0_tz_0 ;
    wire \ALU.madd_104 ;
    wire \ALU.madd_149 ;
    wire \ALU.madd_128_0_tz ;
    wire \ALU.madd_128_0 ;
    wire \ALU.madd_N_1_i ;
    wire \ALU.madd_33 ;
    wire \ALU.madd_68_0_tz ;
    wire \ALU.madd_68 ;
    wire \ALU.madd_89_0 ;
    wire \ALU.madd_68_cascade_ ;
    wire \ALU.a7_b_1 ;
    wire \ALU.madd_108 ;
    wire \ALU.madd_108_cascade_ ;
    wire \ALU.madd_134 ;
    wire \ALU.madd_153 ;
    wire \FTDI.N_201_2 ;
    wire \INVFTDI.RXreadyC_net ;
    wire aluOperation_3;
    wire \ALU.m681Z0Z_1_cascade_ ;
    wire \ALU.N_730_mux ;
    wire \FTDI.N_28 ;
    wire \ALU.a_15_m1_0 ;
    wire \ALU.a_15_m4_ns_1_0_cascade_ ;
    wire \ALU.a_15_m4_0_cascade_ ;
    wire \ALU.a_15_m3_0 ;
    wire \ALU.a_15_m4_bm_1Z0Z_8 ;
    wire \ALU.a_15_m0_0 ;
    wire i53_mux_0;
    wire \ALU.N_273_0 ;
    wire \ALU.N_461 ;
    wire \ALU.N_474 ;
    wire \ALU.N_530_cascade_ ;
    wire \ALU.N_635 ;
    wire \ALU.d_RNIP8ITN1Z0Z_5_cascade_ ;
    wire \ALU.d_RNILBFG4Z0Z_2 ;
    wire \ALU.a_15_m3_2_cascade_ ;
    wire \ALU.d_RNIE937BZ0Z_0_cascade_ ;
    wire \ALU.a_15_m4_2 ;
    wire \ALU.N_257 ;
    wire \ALU.N_249_cascade_ ;
    wire \ALU.N_253 ;
    wire \ALU.c_RNIUGCLVZ0Z_11_cascade_ ;
    wire \ALU.N_415 ;
    wire \ALU.N_310 ;
    wire \ALU.lshift_3_ns_1_4_cascade_ ;
    wire \ALU.N_220 ;
    wire \ALU.N_250 ;
    wire \ALU.N_250_cascade_ ;
    wire \ALU.N_254 ;
    wire \ALU.N_218 ;
    wire \ALU.N_218_cascade_ ;
    wire \ALU.N_361_cascade_ ;
    wire \ALU.N_252 ;
    wire \ALU.m270_nsZ0Z_1_cascade_ ;
    wire ctrlOut_12;
    wire ctrlOut_15;
    wire \ALU.N_7_0_cascade_ ;
    wire \ALU.N_179_0 ;
    wire \ALU.a_15_m2_ns_1Z0Z_13_cascade_ ;
    wire \ALU.operand2_9 ;
    wire \ALU.N_205_0 ;
    wire \ALU.operand2_9_cascade_ ;
    wire \ALU.a_15_m2_ns_1Z0Z_9_cascade_ ;
    wire \ALU.d_RNIO7LUZ0Z_13_cascade_ ;
    wire \ALU.operand2_13_cascade_ ;
    wire \ALU.N_177_0_cascade_ ;
    wire \ALU.madd_484_3 ;
    wire \ALU.madd_484_1 ;
    wire \ALU.madd_484_2_cascade_ ;
    wire \ALU.madd_484_0 ;
    wire \ALU.madd_484_12 ;
    wire \ALU.a0_b_11 ;
    wire bfn_6_9_0_;
    wire \ALU.un2_addsub_cry_0 ;
    wire \ALU.d_RNIEDJEAZ0Z_2 ;
    wire \ALU.N_240_0_i ;
    wire \ALU.un2_addsub_cry_1 ;
    wire \ALU.un2_addsub_cry_2 ;
    wire \ALU.un2_addsub_cry_3 ;
    wire \ALU.d_RNIVR3QAZ0Z_5 ;
    wire \ALU.un2_addsub_cry_4 ;
    wire \ALU.d_RNIGLK5BZ0Z_6 ;
    wire \ALU.un2_addsub_cry_5 ;
    wire \ALU.d_RNITAM9DZ0Z_7 ;
    wire \ALU.un2_addsub_cry_6 ;
    wire \ALU.un2_addsub_cry_7 ;
    wire \ALU.N_201_0 ;
    wire \ALU.d_RNIQ74VBZ0Z_8 ;
    wire bfn_6_10_0_;
    wire \ALU.d_RNI6B7KDZ0Z_9 ;
    wire \ALU.un2_addsub_cry_8 ;
    wire \ALU.N_192_0_i ;
    wire \ALU.un2_addsub_cry_9 ;
    wire \ALU.un2_addsub_cry_10 ;
    wire \ALU.N_180_0_i ;
    wire \ALU.un2_addsub_cry_11 ;
    wire \ALU.un2_addsub_cry_12 ;
    wire \ALU.N_171_0 ;
    wire \ALU.d_RNI1M3JEZ0Z_14 ;
    wire \ALU.un2_addsub_cry_13 ;
    wire \ALU.un2_addsub_cry_14 ;
    wire \ALU.g0_7_a3_0Z0Z_0 ;
    wire \ALU.N_8_1_cascade_ ;
    wire \ALU.g0_2Z0Z_1 ;
    wire \ALU.g0_7_m4_0_1_cascade_ ;
    wire \ALU.N_9_2 ;
    wire \ALU.dout_3_ns_1_0_cascade_ ;
    wire \ALU.dout_6_ns_1_0_cascade_ ;
    wire \ALU.N_747_cascade_ ;
    wire \ALU.aluOut_0_cascade_ ;
    wire \ALU.g0_0_0_N_2L1 ;
    wire \ALU.dout_3_ns_1_7 ;
    wire \ALU.a_15_m5_0 ;
    wire \ALU.d_RNI9BO713Z0Z_0_cascade_ ;
    wire \ALU.operand2_7_ns_1_0_cascade_ ;
    wire ctrlOut_0;
    wire \ALU.operand2_0_cascade_ ;
    wire \ALU.hZ0Z_0 ;
    wire \ALU.d_RNIE4R7Z0Z_0 ;
    wire \ALU.g_RNIT0COZ0Z_1_cascade_ ;
    wire \ALU.operand2_7_ns_1_1_cascade_ ;
    wire \ALU.e_RNIPKVJZ0Z_1 ;
    wire \ALU.madd_4 ;
    wire \ALU.madd_12_0_tz ;
    wire \ALU.dout_6_ns_1_15_cascade_ ;
    wire \ALU.N_752_cascade_ ;
    wire \ALU.dout_3_ns_1_5_cascade_ ;
    wire \ALU.N_704 ;
    wire \ALU.un2_addsub_axb_4_cascade_ ;
    wire \ALU.d_RNI312TBZ0Z_4 ;
    wire \ALU.N_223_0 ;
    wire \ALU.operand2_5 ;
    wire \ALU.a3_b_5_cascade_ ;
    wire \ALU.madd_94 ;
    wire \ALU.a4_b_4 ;
    wire \ALU.a3_b_5 ;
    wire \ALU.a4_b_4_cascade_ ;
    wire \ALU.madd_98 ;
    wire \ALU.N_207_0 ;
    wire \ALU.madd_98_cascade_ ;
    wire \ALU.madd_93 ;
    wire \ALU.madd_139 ;
    wire RX_c;
    wire RXready;
    wire ctrlOut_1;
    wire \ALU.N_41_0_0_cascade_ ;
    wire \ALU.rshift_3_ns_1_5 ;
    wire \ALU.N_473_cascade_ ;
    wire \ALU.m42_nsZ0Z_1 ;
    wire testWordZ0Z_1;
    wire testWordZ0Z_4;
    wire testWordZ0Z_2;
    wire testWordZ0Z_3;
    wire \ALU.N_469_cascade_ ;
    wire \ALU.N_473 ;
    wire \ALU.rshift_15_ns_1_1_cascade_ ;
    wire N_305_0;
    wire \CONTROL.aluParams_cnvZ0Z_0 ;
    wire \ALU.rshift_3_ns_1_9_cascade_ ;
    wire \ALU.rshift_3_ns_1_1 ;
    wire \ALU.d_RNINEO9E_0Z0Z_1 ;
    wire \ALU.N_217 ;
    wire \ALU.lshift_7_ns_1_9 ;
    wire \ALU.N_311_cascade_ ;
    wire \ALU.lshift_9_cascade_ ;
    wire \ALU.a_15_m2_9 ;
    wire \ALU.N_292_0 ;
    wire \ALU.rshift_1 ;
    wire \ALU.d_RNIA28GU1Z0Z_1_cascade_ ;
    wire \ALU.d_RNIJ1PCQZ0Z_1 ;
    wire \ALU.N_225 ;
    wire \ALU.N_223 ;
    wire \ALU.N_221 ;
    wire \ALU.lshift_7_ns_1_13_cascade_ ;
    wire \ALU.N_219 ;
    wire \ALU.N_315_cascade_ ;
    wire \ALU.lshift_13_cascade_ ;
    wire \ALU.a_15_m2_13 ;
    wire \ALU.a_15_m4_13_cascade_ ;
    wire \ALU.N_247 ;
    wire \ALU.lshift_15_ns_1_15 ;
    wire \ALU.N_416 ;
    wire \ALU.N_377 ;
    wire \ALU.N_377_cascade_ ;
    wire \ALU.N_216 ;
    wire \ALU.N_404 ;
    wire \ALU.N_246 ;
    wire \ALU.N_376_cascade_ ;
    wire \ALU.d_RNIEBMRAZ0Z_0_cascade_ ;
    wire \ALU.d_RNI1GH4VZ0Z_7 ;
    wire \ALU.N_468 ;
    wire \ALU.a1_b_3 ;
    wire \ALU.a0_b_4 ;
    wire \ALU.a1_b_3_cascade_ ;
    wire \ALU.madd_0 ;
    wire \ALU.a0_b_3 ;
    wire \ALU.N_375 ;
    wire \ALU.rshift_3_ns_1_0 ;
    wire \ALU.N_249 ;
    wire \ALU.N_245 ;
    wire \ALU.lshift_10 ;
    wire \ALU.a_15_m3_10 ;
    wire \ALU.a_15_m4_10_cascade_ ;
    wire \ALU.a_15_m2_10 ;
    wire \ALU.a_15_m2_ns_1Z0Z_10 ;
    wire \ALU.un2_addsub_cry_9_c_RNIVCOFAZ0 ;
    wire un9_addsub_cry_9_c_RNI8H83V_cascade_;
    wire c_RNI5V90O2_10;
    wire aluOperation_RNINNN4N3_0_cascade_;
    wire \ALU.dout_6_ns_1_11_cascade_ ;
    wire \ALU.dout_3_ns_1_11_cascade_ ;
    wire \ALU.N_758 ;
    wire \ALU.N_710_cascade_ ;
    wire \ALU.aluOut_11_cascade_ ;
    wire \ALU.madd_484_6 ;
    wire \ALU.un2_addsub_axb_1_cascade_ ;
    wire \ALU.d_RNIC4AT9Z0Z_1 ;
    wire \ALU.dout_7_ns_1_1_cascade_ ;
    wire \ALU.N_247_0 ;
    wire \ALU.operand2_1 ;
    wire \ALU.N_249_0 ;
    wire \ALU.N_249_0_cascade_ ;
    wire \ALU.d_RNI61SHAZ0Z_1_cascade_ ;
    wire \ALU.d_RNIJM067Z0Z_1 ;
    wire \ALU.a_15_m2_1 ;
    wire \ALU.g_RNIK6LLZ0Z_4_cascade_ ;
    wire \ALU.e_RNIGQ8HZ0Z_4 ;
    wire \ALU.a1_b_4 ;
    wire \ALU.a2_b_4 ;
    wire \ALU.operand2_7_ns_1_4 ;
    wire \ALU.operand2_4 ;
    wire \ALU.N_229_0 ;
    wire \ALU.operand2_4_cascade_ ;
    wire \ALU.N_231_0_cascade_ ;
    wire \ALU.madd_93_0 ;
    wire \ALU.aZ0Z_10 ;
    wire \ALU.dout_3_ns_1_10_cascade_ ;
    wire \ALU.dout_6_ns_1_10_cascade_ ;
    wire \ALU.N_757_cascade_ ;
    wire \ALU.N_709 ;
    wire \ALU.dout_6_ns_1_5 ;
    wire \ALU.N_865_cascade_ ;
    wire \ALU.operand2_3_ns_1_6_cascade_ ;
    wire \ALU.N_817 ;
    wire \ALU.a6_b_6 ;
    wire \ALU.a3_b_6 ;
    wire \ALU.operand2_6_ns_1_6 ;
    wire \ALU.N_750_cascade_ ;
    wire \ALU.operand2_3_cascade_ ;
    wire \ALU.a3_b_3 ;
    wire aluReadBus_rep1;
    wire \ALU.a2_b_3 ;
    wire \ALU.operand2_3 ;
    wire \ALU.N_235_0 ;
    wire \ALU.un2_addsub_axb_3 ;
    wire \ALU.d_RNIDK21BZ0Z_3 ;
    wire \ALU.dout_3_ns_1_3_cascade_ ;
    wire \ALU.N_702 ;
    wire \ALU.g_RNII4LLZ0Z_3 ;
    wire \ALU.e_RNITOVJZ0Z_3_cascade_ ;
    wire \ALU.operand2_7_ns_1_3 ;
    wire \ALU.un2_addsub_cry_6_c_RNIL4LMIZ0 ;
    wire \ALU.a7_b_0 ;
    wire \ALU.a5_b_2 ;
    wire \ALU.madd_63 ;
    wire \ALU.a2_b_1 ;
    wire \ALU.a3_b_0 ;
    wire \ALU.a1_b_2 ;
    wire \ALU.d_RNI2B0LZ0Z_9 ;
    wire \ALU.hZ0Z_10 ;
    wire \ALU.d_RNII1LUZ0Z_10 ;
    wire \ALU.d_RNIO00LZ0Z_4 ;
    wire \FTDI.RXstateZ0Z_2 ;
    wire \FTDI.N_23_cascade_ ;
    wire \FTDI.RXstateZ0Z_1 ;
    wire \FTDI.m13_ns_1 ;
    wire \FTDI.RXstateZ0Z_0 ;
    wire \FTDI.RXstateZ0Z_3 ;
    wire \INVFTDI.gap_0C_net ;
    wire \ALU.a_15_sm0_cascade_ ;
    wire \ALU.a_15_m2_ns_1Z0Z_12_cascade_ ;
    wire \ALU.log_2_sqmuxa ;
    wire \ALU.a_15_m4_bm_1Z0Z_2_cascade_ ;
    wire \ALU.d_RNIII58AZ0Z_2 ;
    wire \ALU.rshift_3_ns_1_2_cascade_ ;
    wire \ALU.N_470 ;
    wire \ALU.N_376 ;
    wire \ALU.N_589_cascade_ ;
    wire \ALU.rshift_1_13_cascade_ ;
    wire \ALU.a_15_m3_13 ;
    wire \ALU.N_576_cascade_ ;
    wire \ALU.N_636_cascade_ ;
    wire \ALU.N_272_0 ;
    wire \ALU.N_264_0 ;
    wire \ALU.aluOut_12 ;
    wire \ALU.N_462 ;
    wire \ALU.N_270_0 ;
    wire aluReadBus_fast;
    wire \ALU.N_175_0 ;
    wire \ALU.N_175_0_cascade_ ;
    wire \ALU.operand2_13 ;
    wire \ALU.un2_addsub_axb_13_cascade_ ;
    wire \ALU.N_177_0 ;
    wire \ALU.d_RNI9FOTEZ0Z_13 ;
    wire ctrlOut_11;
    wire \ALU.N_186_0_i ;
    wire \ALU.N_186_0_i_cascade_ ;
    wire \ALU.c_RNIA7OEEZ0Z_11 ;
    wire RXbuffer_5;
    wire \ALU.hZ0Z_12 ;
    wire \ALU.c_RNIJ949Z0Z_12_cascade_ ;
    wire \ALU.a_RNIFPBOZ0Z_12 ;
    wire \ALU.d_RNIM5LUZ0Z_12 ;
    wire \ALU.operand2_7_ns_1_12_cascade_ ;
    wire \ALU.operand2_12 ;
    wire \ALU.d_RNICJE9BZ0Z_8 ;
    wire \ALU.d_RNIEUKR11Z0Z_0 ;
    wire \ALU.a_15_m3_8 ;
    wire \ALU.a_15_m4_8_cascade_ ;
    wire \ALU.a_15_m5_8 ;
    wire \ALU.fZ0Z_8 ;
    wire \ALU.dZ0Z_8 ;
    wire \ALU.operand2_6_ns_1_8_cascade_ ;
    wire \ALU.N_867 ;
    wire \ALU.hZ0Z_8 ;
    wire \ALU.fZ0Z_15 ;
    wire \ALU.madd_cry_0_ma ;
    wire bfn_9_9_0_;
    wire \ALU.madd_cry_1_ma ;
    wire \ALU.madd_cry_0 ;
    wire \ALU.madd_axb_2_l_fx ;
    wire \ALU.madd_6 ;
    wire \ALU.madd_cry_1 ;
    wire \ALU.madd_13 ;
    wire \ALU.madd_18 ;
    wire \ALU.madd_cry_2 ;
    wire \ALU.madd_axb_4_l_fx ;
    wire \ALU.madd_30 ;
    wire \ALU.madd_cry_3 ;
    wire \ALU.madd_52 ;
    wire \ALU.madd_axb_5_l_fx ;
    wire \ALU.madd_cry_4 ;
    wire \ALU.madd_cry_5 ;
    wire \ALU.madd_axb_7 ;
    wire \ALU.madd_cry_6_THRU_CO ;
    wire \ALU.madd_cry_6 ;
    wire \ALU.madd_cry_7 ;
    wire \ALU.madd_axb_8_l_fx ;
    wire \ALU.madd_159 ;
    wire bfn_9_10_0_;
    wire \ALU.madd_cry_9_ma ;
    wire \ALU.madd_axb_9_l_ofx ;
    wire \ALU.madd_cry_8 ;
    wire \ALU.madd_cry_10_ma ;
    wire \ALU.madd_axb_10_l_ofx ;
    wire \ALU.madd_cry_9 ;
    wire \ALU.madd_axb_11 ;
    wire \ALU.madd_cry_10 ;
    wire \ALU.madd_axb_12_l_fx ;
    wire \ALU.madd_360 ;
    wire \ALU.madd_cry_11 ;
    wire \ALU.madd_cry_13_ma ;
    wire \ALU.madd_axb_13_l_ofx ;
    wire \ALU.madd_cry_12 ;
    wire \ALU.madd_axb_14 ;
    wire \ALU.madd_cry_13 ;
    wire \ALU.operand2_6 ;
    wire aluReadBus;
    wire \ALU.N_217_0 ;
    wire \ALU.dout_3_ns_1_15_cascade_ ;
    wire \ALU.dout_6_ns_1_2_cascade_ ;
    wire \ALU.N_749_cascade_ ;
    wire \ALU.N_701 ;
    wire \ALU.dout_3_ns_1_2 ;
    wire \ALU.dout_6_ns_1_7 ;
    wire \ALU.f_RNIQQJ01Z0Z_7 ;
    wire testWordZ0Z_8;
    wire \ALU.fZ0Z_10 ;
    wire \ALU.b_RNIEHSD1Z0Z_10 ;
    wire \ALU.dout_3_ns_1_4 ;
    wire \ALU.eZ0Z_4 ;
    wire \ALU.e_RNIS97JZ0Z_1 ;
    wire \ALU.eZ0Z_1 ;
    wire \ALU.g_RNI0MJNZ0Z_1 ;
    wire \ALU.dout_6_ns_1_3 ;
    wire aluOperand1_2_rep1;
    wire \ALU.dout_6_ns_1_4 ;
    wire \ALU.N_747 ;
    wire \ALU.N_699 ;
    wire \ALU.N_404_1 ;
    wire \ALU.dout_6_ns_1_6 ;
    wire \ALU.N_753_cascade_ ;
    wire testWordZ0Z_9;
    wire aluOperand1_fast_1;
    wire aluOperand1_fast_2;
    wire \ALU.dout_3_ns_1_6_cascade_ ;
    wire \ALU.N_705 ;
    wire testWordZ0Z_7;
    wire \CONTROL.operand1_cnvZ0Z_0 ;
    wire \ALU.c_RNI72MICZ0Z_15_cascade_ ;
    wire \ALU.d_RNI4HG101Z0Z_7 ;
    wire \INVFTDI.baudAcc_0C_net ;
    wire \ALU.aluOut_10 ;
    wire \ALU.N_475_cascade_ ;
    wire \ALU.rshift_7 ;
    wire \ALU.rshift_15_ns_1_7 ;
    wire \ALU.rshift_3_ns_1_3_cascade_ ;
    wire \ALU.N_471_cascade_ ;
    wire \ALU.N_475 ;
    wire \ALU.rshift_3_ns_1_7 ;
    wire \ALU.N_576 ;
    wire \ALU.a_15_m5_5_cascade_ ;
    wire \ALU.mult_5 ;
    wire \ALU.d_RNIPFIBI1Z0Z_9 ;
    wire \ALU.a_15_m2_ns_1Z0Z_5_cascade_ ;
    wire \ALU.N_225_0 ;
    wire \ALU.a_15_m2_5_cascade_ ;
    wire \ALU.N_420 ;
    wire \ALU.a_15_m4_5 ;
    wire a_4;
    wire a_6;
    wire a_7;
    wire \ALU.a_15_m2_12 ;
    wire \ALU.a_15_m4_12_cascade_ ;
    wire \ALU.un2_addsub_cry_11_c_RNII7OFZ0Z9 ;
    wire un2_addsub_cry_11_c_RNIQ9LMU_cascade_;
    wire c_RNIC8RDN2_12;
    wire aluOperation_RNIGPL5M3_0_cascade_;
    wire \ALU.aZ0Z_12 ;
    wire \ALU.N_271_0 ;
    wire \ALU.a_15_m3_12 ;
    wire \ALU.N_314 ;
    wire \ALU.lshift_12 ;
    wire \ALU.fZ0Z_9 ;
    wire \ALU.bZ0Z_9 ;
    wire \ALU.f_RNIUUJ01Z0Z_9 ;
    wire \ALU.bZ0Z_12 ;
    wire \ALU.fZ0Z_12 ;
    wire \ALU.b_RNIILSD1Z0Z_12 ;
    wire \ALU.fZ0Z_14 ;
    wire \ALU.bZ0Z_14 ;
    wire \ALU.g0_3_1_cascade_ ;
    wire \ALU.N_703_0_0 ;
    wire \ALU.N_4 ;
    wire \ALU.N_5 ;
    wire \ALU.fZ0Z_11 ;
    wire \ALU.bZ0Z_11 ;
    wire \ALU.b_RNIKNSD1Z0Z_13 ;
    wire \ALU.dZ0Z_10 ;
    wire \ALU.dZ0Z_12 ;
    wire \ALU.eZ0Z_10 ;
    wire \ALU.eZ0Z_12 ;
    wire \ALU.d_RNIPER7Z0Z_5 ;
    wire \ALU.bZ0Z_10 ;
    wire \ALU.bZ0Z_15 ;
    wire \ALU.un2_addsub_cry_12_c_RNIUL1GKZ0 ;
    wire un2_addsub_cry_12_c_RNIG3PMU_cascade_;
    wire c_RNI88B4N2_13;
    wire aluOperation_RNI2J9SL3_0_cascade_;
    wire \ALU.mult_2 ;
    wire \ALU.a_15_m5_2 ;
    wire \ALU.d_RNIIFMN04Z0Z_2_cascade_ ;
    wire \ALU.eZ0Z_3 ;
    wire \ALU.eZ0Z_6 ;
    wire \ALU.eZ0Z_7 ;
    wire \ALU.eZ0Z_2 ;
    wire a_2;
    wire \ALU.g_RNIV2COZ0Z_2_cascade_ ;
    wire \ALU.e_RNIRMVJZ0Z_2 ;
    wire \ALU.operand2_7_ns_1_2_cascade_ ;
    wire \ALU.operand2_2 ;
    wire \ALU.eZ0Z_0 ;
    wire a_0;
    wire \ALU.e_RNINIVJZ0Z_0 ;
    wire \ALU.g_RNIM8LLZ0Z_5 ;
    wire \ALU.e_RNI1TVJZ0Z_5_cascade_ ;
    wire \ALU.operand2_7_ns_1_5 ;
    wire \ALU.eZ0Z_5 ;
    wire \ALU.g_RNIRUBOZ0Z_0 ;
    wire \ALU.d_RNIG6R7Z0Z_1 ;
    wire \ALU.d_RNI45J9Z0Z_1 ;
    wire \ALU.d_RNII8R7Z0Z_2 ;
    wire \ALU.cZ0Z_0 ;
    wire \ALU.cZ0Z_1 ;
    wire \ALU.cZ0Z_2 ;
    wire \ALU.cZ0Z_3 ;
    wire \ALU.cZ0Z_4 ;
    wire \ALU.cZ0Z_5 ;
    wire \ALU.cZ0Z_6 ;
    wire \ALU.dZ0Z_4 ;
    wire \ALU.gZ0Z_6 ;
    wire \FTDI.gapZ0Z_2 ;
    wire \FTDI.gapZ0Z_0 ;
    wire \FTDI.gap8 ;
    wire \FTDI.gapZ0Z_1 ;
    wire \INVFTDI.gap_2C_net ;
    wire \FTDI.TXstate_e_1_0 ;
    wire \FTDI.N_169_0_cascade_ ;
    wire \FTDI.N_169_0 ;
    wire \FTDI.TXstate_cnst_0_0_2_cascade_ ;
    wire \INVFTDI.TXstate_0C_net ;
    wire \FTDI.N_217_0_cascade_ ;
    wire \FTDI.N_216_0 ;
    wire \FTDI.TXready_cascade_ ;
    wire \FTDI.baudAccZ0Z_0 ;
    wire \FTDI.baudAccZ0Z_1 ;
    wire \ALU.N_290_0 ;
    wire \ALU.rshift_5 ;
    wire \ALU.a_15_m3_5 ;
    wire \FTDI.TXstateZ1Z_0 ;
    wire \FTDI.TXstateZ1Z_1 ;
    wire \FTDI.N_170_0 ;
    wire \FTDI.TXstate_e_1_3_cascade_ ;
    wire \INVFTDI.baudAcc_1C_net ;
    wire \ALU.N_11_0 ;
    wire \ALU.N_5_0 ;
    wire \ALU.c_RNI1OCN4Z0Z_15_cascade_ ;
    wire \ALU.N_762 ;
    wire \ALU.N_714 ;
    wire \ALU.N_621_1_cascade_ ;
    wire \ALU.N_589 ;
    wire \ALU.N_621_1 ;
    wire \ALU.c_RNI4JFV4_0Z0Z_15 ;
    wire \ALU.N_274_0 ;
    wire \ALU.d_RNI36KJ21Z0Z_9 ;
    wire \FTDI.TXready ;
    wire \FTDI.baudAccZ0Z_2 ;
    wire TXstartZ0;
    wire testStateZ0Z_0;
    wire ctrlOut_13;
    wire busState_2;
    wire aluReadBus_rep2;
    wire busState_0;
    wire \ALU.N_9_1 ;
    wire testStateZ0Z_2;
    wire testState_i_2;
    wire \ALU.eZ0Z_14 ;
    wire \ALU.un2_addsub_cry_13_c_RNINVE5KZ0 ;
    wire un2_addsub_cry_13_c_RNI2LH1U_cascade_;
    wire c_RNIFCGVL2_14;
    wire aluOperation_RNIR872K3_0_cascade_;
    wire \ALU.a_RNIJTBOZ0Z_14 ;
    wire \ALU.operand2_7_ns_1_14_cascade_ ;
    wire \ALU.b_RNIMPSD1Z0Z_14 ;
    wire \ALU.operand2_14 ;
    wire \ALU.hZ0Z_14 ;
    wire \ALU.dZ0Z_14 ;
    wire \ALU.d_RNIQ9LUZ0Z_14 ;
    wire \ALU.un2_addsub_cry_7_c_RNIL8JHGZ0 ;
    wire \ALU.aZ0Z_8 ;
    wire aluOperand2_fast_1;
    wire \ALU.eZ0Z_8 ;
    wire \ALU.gZ0Z_8 ;
    wire \ALU.cZ0Z_8 ;
    wire \ALU.operand2_3_ns_1_8_cascade_ ;
    wire \ALU.N_819 ;
    wire \ALU.addsub_0_sqmuxa_cascade_ ;
    wire \ALU.un2_addsub_cry_8_c_RNIKR81JZ0 ;
    wire \ALU.un9_addsub_cry_8_c_RNIKTS9SZ0_cascade_ ;
    wire \ALU.a_15_m5_9 ;
    wire \ALU.a_15_ns_1_9_cascade_ ;
    wire \ALU.eZ0Z_11 ;
    wire aluOperand2_0_rep1;
    wire \ALU.a_RNICNBOZ0Z_11_cascade_ ;
    wire \ALU.operand2_7_ns_1_11_cascade_ ;
    wire \ALU.b_RNIGJSD1Z0Z_11 ;
    wire \ALU.operand2_11 ;
    wire \ALU.dZ0Z_11 ;
    wire \ALU.d_RNIK3LUZ0Z_11 ;
    wire \ALU.hZ0Z_11 ;
    wire \ALU.c_RNIG749Z0Z_11 ;
    wire \ALU.a_RNIHRBOZ0Z_13_cascade_ ;
    wire \ALU.c_RNILB49Z0Z_13 ;
    wire \ALU.operand2_7_ns_1_13 ;
    wire \ALU.eZ0Z_15 ;
    wire \ALU.a_RNILVBOZ0Z_15_cascade_ ;
    wire \ALU.c_RNIPF49Z0Z_15 ;
    wire \ALU.operand2_7_ns_1_15_cascade_ ;
    wire \ALU.b_RNIORSD1Z0Z_15 ;
    wire \ALU.operand2_15 ;
    wire \ALU.cZ0Z_11 ;
    wire \ALU.cZ0Z_12 ;
    wire \ALU.cZ0Z_14 ;
    wire \ALU.c_RNIND49Z0Z_14 ;
    wire \ALU.cZ0Z_15 ;
    wire \ALU.c_cnvZ0Z_0 ;
    wire \ALU.hZ0Z_1 ;
    wire \ALU.hZ0Z_2 ;
    wire \ALU.hZ0Z_5 ;
    wire \ALU.aZ0Z_14 ;
    wire \ALU.aZ0Z_15 ;
    wire \ALU.f_RNI0P6LZ0Z_1 ;
    wire \ALU.f_RNICQEJZ0Z_1 ;
    wire \ALU.cZ0Z_7 ;
    wire \ALU.g_RNIQCLLZ0Z_7 ;
    wire \ALU.f_RNIL2FJZ0Z_5 ;
    wire \ALU.m286_bmZ0 ;
    wire \ALU.m286_amZ0 ;
    wire \ALU.f_RNIAOEJZ0Z_0 ;
    wire aluOperand2_fast_0;
    wire aluOperand2_2_rep1;
    wire \ALU.bZ0Z_2 ;
    wire \ALU.f_RNIESEJZ0Z_2 ;
    wire \ALU.gZ0Z_0 ;
    wire \ALU.gZ0Z_1 ;
    wire \ALU.gZ0Z_2 ;
    wire \ALU.gZ0Z_3 ;
    wire \ALU.gZ0Z_4 ;
    wire \ALU.gZ0Z_5 ;
    wire \ALU.gZ0Z_7 ;
    wire \ALU.N_578 ;
    wire \ALU.N_477 ;
    wire \ALU.N_634 ;
    wire CONSTANT_ONE_NET;
    wire \FTDI.un3_TX_0 ;
    wire RXbuffer_4;
    wire testWordZ0Z_12;
    wire TXbufferZ0Z_0;
    wire TXbufferZ0Z_3;
    wire \FTDI.TXshiftZ0Z_5 ;
    wire TXbufferZ0Z_4;
    wire \FTDI.TXshiftZ0Z_4 ;
    wire \FTDI.TXshiftZ0Z_3 ;
    wire TXbufferZ0Z_2;
    wire TXbufferZ0Z_6;
    wire \FTDI.TXshiftZ0Z_6 ;
    wire TXbufferZ0Z_7;
    wire \FTDI.TXshiftZ0Z_7 ;
    wire \INVFTDI.TXshift_0C_net ;
    wire \ALU.un2_addsub_cry_10_c_RNIUS1OJZ0 ;
    wire \ALU.a_15_m2_ns_1Z0Z_11_cascade_ ;
    wire \ALU.a_15_m2_11_cascade_ ;
    wire \ALU.lshift_11 ;
    wire \ALU.a_15_m4_11_cascade_ ;
    wire \ALU.a_15_m3_11 ;
    wire c_RNID7K8N2_11_cascade_;
    wire un2_addsub_cry_10_c_RNIEBKOT;
    wire aluOperation_RNI5QD2L3_0_cascade_;
    wire \ALU.aZ0Z_11 ;
    wire \ALU.e_cnvZ0Z_0 ;
    wire \ALU.g_RNIVGLLZ0Z_9_cascade_ ;
    wire \ALU.operand2_7_ns_1_9 ;
    wire \ALU.hZ0Z_9 ;
    wire \ALU.dZ0Z_9 ;
    wire \ALU.g0_0_0_m2_1 ;
    wire \ALU.N_11_cascade_ ;
    wire \ALU.N_13 ;
    wire \ALU.cZ0Z_9 ;
    wire \ALU.g0_0_0_m2_0_1 ;
    wire \ALU.N_12 ;
    wire \ALU.aluOut_15 ;
    wire \ALU.a_15_m2_ns_1Z0Z_15_cascade_ ;
    wire \ALU.N_7_0 ;
    wire \ALU.a_15_m2_15_cascade_ ;
    wire \ALU.lshift_15 ;
    wire \ALU.a_15_m4_15_cascade_ ;
    wire \ALU.a_15_m3_15 ;
    wire \ALU.c_RNIR4QHM2Z0Z_15_cascade_ ;
    wire \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93_cascade_ ;
    wire \ALU.hZ0Z_15 ;
    wire \ALU.dZ0Z_15 ;
    wire \ALU.d_RNISBLUZ0Z_15 ;
    wire \CONTROL.aluOperation_cnvZ0Z_0 ;
    wire N_723;
    wire testWordZ0Z_5;
    wire aluOperation_5;
    wire \ALU.a2_b_0 ;
    wire \ALU.madd_axb_1_l_ofx ;
    wire aluOperand2_0_rep2;
    wire aluOperand2_0;
    wire aluOperand2_1_rep1;
    wire \ALU.cZ0Z_10 ;
    wire aluOperand2_fast_2;
    wire \ALU.g0_7_m4_1 ;
    wire N_287_0;
    wire G_566;
    wire testWordZ0Z_11;
    wire aluOperand2_1;
    wire \ALU.mult_10 ;
    wire aluOperation_RNINNN4N3_0;
    wire \ALU.gZ0Z_10 ;
    wire aluOperation_RNI5QD2L3_0;
    wire \ALU.mult_11 ;
    wire \ALU.gZ0Z_11 ;
    wire aluOperation_RNIGPL5M3_0;
    wire \ALU.mult_12 ;
    wire \ALU.gZ0Z_12 ;
    wire aluOperation_RNI2J9SL3_0;
    wire \ALU.mult_13 ;
    wire aluOperation_RNIR872K3_0;
    wire \ALU.mult_14 ;
    wire \ALU.gZ0Z_14 ;
    wire \ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93 ;
    wire \ALU.mult_15 ;
    wire \ALU.gZ0Z_15 ;
    wire \ALU.a_15_ns_1_9 ;
    wire \ALU.mult_9 ;
    wire \ALU.gZ0Z_9 ;
    wire \ALU.g_cnvZ0Z_0 ;
    wire \ALU.eZ0Z_13 ;
    wire \ALU.aZ0Z_13 ;
    wire aluOperand1_2_rep2;
    wire aluOperand1_1_rep1;
    wire \ALU.cZ0Z_13 ;
    wire \ALU.dout_3_ns_1_13_cascade_ ;
    wire \ALU.gZ0Z_13 ;
    wire \ALU.bZ0Z_13 ;
    wire aluOperand1_1_rep2;
    wire \ALU.fZ0Z_13 ;
    wire aluOperand1_2;
    wire \ALU.hZ0Z_13 ;
    wire \ALU.dZ0Z_13 ;
    wire \ALU.dout_6_ns_1_13_cascade_ ;
    wire aluOperand1_1;
    wire \ALU.N_712 ;
    wire \ALU.N_760_cascade_ ;
    wire aluOperand1_0;
    wire \ALU.aluOut_13_cascade_ ;
    wire \ALU.a13_b_0 ;
    wire \ALU.fZ0Z_0 ;
    wire \ALU.fZ0Z_1 ;
    wire \ALU.fZ0Z_2 ;
    wire \ALU.fZ0Z_5 ;
    wire \ALU.fZ0Z_6 ;
    wire \ALU.fZ0Z_7 ;
    wire \ALU.f_cnvZ0Z_0 ;
    wire \ALU.N_1700_i ;
    wire \ALU.d_RNIO75MAZ0Z_0_cascade_ ;
    wire \ALU.bZ0Z_0 ;
    wire \ALU.madd_axb_0_l_ofx ;
    wire \ALU.mult_1_cascade_ ;
    wire \ALU.a_15_m5_1 ;
    wire \ALU.d_RNIEICQ63Z0Z_1_cascade_ ;
    wire \ALU.bZ0Z_1 ;
    wire \ALU.d_RNIEICQ63Z0Z_1 ;
    wire \ALU.dZ0Z_1 ;
    wire \ALU.hZ0Z_4 ;
    wire \FTDI.un3_TX_0_i ;
    wire bfn_13_2_0_;
    wire \FTDI.un3_TX_axb_3 ;
    wire \FTDI.un3_TX_cry_2 ;
    wire \FTDI.TXshiftZ0Z_0 ;
    wire \FTDI.un3_TX_cry_3 ;
    wire FTDI_TX_0_i;
    wire \ALU.N_361 ;
    wire \ALU.N_244 ;
    wire aluParams_1;
    wire \ALU.N_588 ;
    wire aluParams_2;
    wire \ALU.N_590 ;
    wire \ALU.eZ0Z_9 ;
    wire \ALU.aZ0Z_9 ;
    wire \ALU.e_RNIR49HZ0Z_9 ;
    wire \ALU.N_252_0 ;
    wire \ALU.aluOut_0 ;
    wire \ALU.a0_b_2 ;
    wire bfn_13_7_0_;
    wire \ALU.N_249_0_i ;
    wire \ALU.aluOut_1 ;
    wire \ALU.un9_addsub_cry_0 ;
    wire \ALU.N_240_0 ;
    wire \ALU.aluOut_2 ;
    wire \ALU.un9_addsub_cry_1 ;
    wire \ALU.N_237_0_i ;
    wire \ALU.un9_addsub_cry_2 ;
    wire \ALU.N_231_0_i ;
    wire \ALU.un9_addsub_cry_3 ;
    wire \ALU.aluOut_5 ;
    wire \ALU.N_225_0_i ;
    wire \ALU.un9_addsub_cry_4 ;
    wire \ALU.N_219_0_i ;
    wire \ALU.un9_addsub_cry_5 ;
    wire \ALU.N_213_0_i ;
    wire \ALU.un9_addsub_cry_6_c_RNI2EFHZ0Z8 ;
    wire \ALU.un9_addsub_cry_6 ;
    wire \ALU.un9_addsub_cry_7 ;
    wire \ALU.aluOut_8 ;
    wire \ALU.N_201_0_i ;
    wire \ALU.un9_addsub_cry_7_c_RNIU7FZ0Z18 ;
    wire bfn_13_8_0_;
    wire \ALU.aluOut_9 ;
    wire \ALU.N_207_0_i ;
    wire \ALU.un9_addsub_cry_8_c_RNIPV1SZ0Z8 ;
    wire \ALU.un9_addsub_cry_8 ;
    wire \ALU.N_192_0 ;
    wire \ALU.a_RNIV2S0FZ0Z_10 ;
    wire \ALU.un9_addsub_cry_9_c_RNI22U6KZ0 ;
    wire \ALU.un9_addsub_cry_9 ;
    wire \ALU.N_186_0 ;
    wire \ALU.aluOut_11 ;
    wire \ALU.un9_addsub_cry_10_c_RNI9C0KZ0Z9 ;
    wire \ALU.un9_addsub_cry_10 ;
    wire \ALU.N_180_0 ;
    wire \ALU.d_RNIFKNTEZ0Z_12 ;
    wire \ALU.un9_addsub_cry_11_c_RNI10BQKZ0 ;
    wire \ALU.un9_addsub_cry_11 ;
    wire \ALU.aluOut_13 ;
    wire \ALU.N_177_0_i ;
    wire \ALU.un9_addsub_cry_12_c_RNIBB5QZ0Z9 ;
    wire \ALU.un9_addsub_cry_12 ;
    wire \ALU.aluOut_14 ;
    wire \ALU.N_171_0_i ;
    wire \ALU.un9_addsub_cry_13_c_RNI4JGFZ0Z9 ;
    wire \ALU.un9_addsub_cry_13 ;
    wire \ALU.un9_addsub_axb_15 ;
    wire \ALU.un2_addsub_cry_14_c_RNINOKZ0Z69 ;
    wire \ALU.un9_addsub_cry_14 ;
    wire \ALU.un9_addsub_cry_14_c_RNIS374JZ0 ;
    wire \ALU.c_RNIA9V4LZ0Z_15 ;
    wire \ALU.d_RNI9DPVUZ0Z_6 ;
    wire \ALU.rshift_3_cascade_ ;
    wire \ALU.N_293_0 ;
    wire \ALU.d_RNI3V2CP1Z0Z_3_cascade_ ;
    wire \ALU.aluOut_3 ;
    wire \ALU.a_15_m2_ns_1Z0Z_3 ;
    wire \ALU.N_237_0 ;
    wire \ALU.a_15_m2_3_cascade_ ;
    wire \ALU.lshift_1_3 ;
    wire \ALU.d_RNI95MLPZ0Z_3 ;
    wire \ALU.mult_3 ;
    wire \ALU.a_15_m5_3 ;
    wire RXbuffer_2;
    wire testStateZ0Z_1;
    wire \ALU.N_58_0 ;
    wire testWordZ0Z_10;
    wire testState_i_g_2;
    wire \ALU.un9_addsub_cry_0_c_RNI2UZ0Z096 ;
    wire \ALU.un2_addsub_cry_0_c_RNI5MA0EZ0 ;
    wire \ALU.un9_addsub_cry_0_c_RNIEMTLKZ0 ;
    wire \ALU.un9_addsub_cry_1_c_RNI6TDZ0Z17 ;
    wire \ALU.un2_addsub_cry_1_c_RNI966GEZ0 ;
    wire \ALU.un9_addsub_cry_2_c_RNIA3LGZ0Z7 ;
    wire \ALU.un2_addsub_cry_2_c_RNI5IV5FZ0 ;
    wire \ALU.un2_addsub_cry_3_c_RNIOGGJGZ0 ;
    wire \ALU.un9_addsub_cry_3_c_RNI525RZ0Z7 ;
    wire \ALU.un9_addsub_cry_4_c_RNIL4NZ0Z97 ;
    wire \ALU.un2_addsub_cry_4_c_RNI284VEZ0 ;
    wire \ALU.un9_addsub_cry_5_c_RNI6SCFZ0Z7 ;
    wire \ALU.addsub_0_sqmuxa ;
    wire \ALU.un2_addsub_cry_5_c_RNIL7IGFZ0 ;
    wire \ALU.N_422 ;
    wire \ALU.d_RNIP43E91Z0Z_7_cascade_ ;
    wire \ALU.d_RNIT87FA1Z0Z_7 ;
    wire \ALU.madd_cry_5_THRU_CO ;
    wire \ALU.a_15_m5_7_cascade_ ;
    wire \ALU.madd_axb_6 ;
    wire \ALU.d_RNIO75MAZ0Z_0 ;
    wire \ALU.d_RNI9BO713Z0Z_0 ;
    wire \ALU.dZ0Z_0 ;
    wire \ALU.un9_addsub_cry_1_c_RNIM56ULZ0 ;
    wire \ALU.d_RNIIFMN04Z0Z_2 ;
    wire \ALU.dZ0Z_2 ;
    wire \ALU.dZ0Z_5 ;
    wire \ALU.dZ0Z_6 ;
    wire \ALU.d_cnvZ0Z_0 ;
    wire \ALU.fZ0Z_3 ;
    wire \ALU.f_RNIHUEJZ0Z_3 ;
    wire \ALU.rshift_1_12 ;
    wire \ALU.N_532 ;
    wire aluOperation_4;
    wire \ALU.rshift_4_cascade_ ;
    wire \ALU.N_289_0 ;
    wire \ALU.a_15_m3_4_cascade_ ;
    wire \ALU.aluOut_4 ;
    wire \ALU.a_15_m2_ns_1Z0Z_4 ;
    wire \ALU.N_231_0 ;
    wire \ALU.a_15_m2_4_cascade_ ;
    wire \ALU.N_419 ;
    wire \ALU.a_15_m4_4 ;
    wire \ALU.mult_4 ;
    wire \ALU.a_15_m5_4 ;
    wire a_3;
    wire \ALU.a_cnvZ0Z_0 ;
    wire \FTDI.TXshiftZ0Z_2 ;
    wire \FTDI.TXstateZ0Z_3 ;
    wire \FTDI.TXshiftZ0Z_1 ;
    wire \INVFTDI.TXshift_1C_net ;
    wire \FTDI.un1_TXstate_0_sqmuxa_0_i ;
    wire a_5;
    wire TXbufferZ0Z_5;
    wire a_1;
    wire TXbufferZ0Z_1;
    wire m326dup;
    wire aluParams_3;
    wire \ALU.N_308 ;
    wire aluOperation_2;
    wire \ALU.log_0_sqmuxa ;
    wire aluParams_0;
    wire \ALU.aluOut_6 ;
    wire \ALU.a_15_m2_ns_1Z0Z_6_cascade_ ;
    wire \ALU.N_219_0 ;
    wire \ALU.a_15_m2_6 ;
    wire \ALU.a_15_sm3 ;
    wire \ALU.d_RNIL01TD1Z0Z_6 ;
    wire \ALU.d_RNIJ75U41Z0Z_6 ;
    wire aluOperation_1;
    wire \ALU.a_15_m5_6_cascade_ ;
    wire \ALU.mult_6 ;
    wire \ALU.d_RNILPR7TQZ0Z_6_cascade_ ;
    wire \ALU.hZ0Z_6 ;
    wire \ALU.h_cnvZ0Z_0 ;
    wire \ALU.fZ0Z_4 ;
    wire \ALU.f_RNIJ0FJZ0Z_4 ;
    wire \ALU.hZ0Z_7 ;
    wire \ALU.dZ0Z_7 ;
    wire aluOperand2_2;
    wire \ALU.d_RNIU60LZ0Z_7 ;
    wire \ALU.hZ0Z_3 ;
    wire \ALU.dZ0Z_3 ;
    wire aluOperand2_2_rep2;
    wire \ALU.d_RNILAR7Z0Z_3 ;
    wire \ALU.un9_addsub_cry_2_c_RNIMN63NZ0 ;
    wire \ALU.d_RNIE8SJN5Z0Z_3 ;
    wire \ALU.bZ0Z_3 ;
    wire \ALU.un9_addsub_cry_3_c_RNI4L7ROZ0 ;
    wire \ALU.d_RNIMA3938Z0Z_4 ;
    wire \ALU.bZ0Z_4 ;
    wire \ALU.un9_addsub_cry_4_c_RNIUEDLMZ0 ;
    wire \ALU.d_RNIH1NE6FZ0Z_5 ;
    wire \ALU.bZ0Z_5 ;
    wire \ALU.d_RNILPR7TQZ0Z_6 ;
    wire \ALU.un9_addsub_cry_5_c_RNI26HCNZ0 ;
    wire \ALU.bZ0Z_6 ;
    wire \ALU.un9_addsub_cry_6_c_RNIUKMKRZ0 ;
    wire \ALU.d_RNIIIPM081Z0Z_7 ;
    wire \ALU.bZ0Z_7 ;
    wire aluOperation_0;
    wire \ALU.un9_addsub_cry_7_c_RNIQIKVOZ0 ;
    wire \ALU.d_RNI7GCMD22Z0Z_8 ;
    wire \ALU.bZ0Z_8 ;
    wire CLK_0_c_g;
    wire \ALU.b_cnvZ0Z_0 ;
    wire \ALU.a_15_sm0 ;
    wire \ALU.N_213_0 ;
    wire \ALU.a_15_m2_ns_1Z0Z_7 ;
    wire \ALU.aluOut_7 ;
    wire \ALU.a_15_m2_7 ;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__49533),
            .GLOBALBUFFEROUTPUT(CLK_0_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__49535),
            .DIN(N__49534),
            .DOUT(N__49533),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__49535),
            .PADOUT(N__49534),
            .PADIN(N__49533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO11_obuf_iopad (
            .OE(N__49524),
            .DIN(N__49523),
            .DOUT(N__49522),
            .PACKAGEPIN(GPIO11));
    defparam GPIO11_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO11_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO11_obuf_preio (
            .PADOEN(N__49524),
            .PADOUT(N__49523),
            .PADIN(N__49522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO9_obuf_iopad (
            .OE(N__49515),
            .DIN(N__49514),
            .DOUT(N__49513),
            .PACKAGEPIN(GPIO9));
    defparam GPIO9_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO9_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO9_obuf_preio (
            .PADOEN(N__49515),
            .PADOUT(N__49514),
            .PADIN(N__49513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32362),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TX_obuf_iopad (
            .OE(N__49506),
            .DIN(N__49505),
            .DOUT(N__49504),
            .PACKAGEPIN(TX));
    defparam TX_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TX_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TX_obuf_preio (
            .PADOEN(N__49506),
            .PADOUT(N__49505),
            .PADIN(N__49504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36485),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO3_obuf_iopad (
            .OE(N__49497),
            .DIN(N__49496),
            .DOUT(N__49495),
            .PACKAGEPIN(GPIO3));
    defparam GPIO3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO GPIO3_obuf_preio (
            .PADOEN(N__49497),
            .PADOUT(N__49496),
            .PADIN(N__49495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15686),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RX_ibuf_iopad (
            .OE(N__49488),
            .DIN(N__49487),
            .DOUT(N__49486),
            .PACKAGEPIN(RX));
    defparam RX_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RX_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RX_ibuf_preio (
            .PADOEN(N__49488),
            .PADOUT(N__49487),
            .PADIN(N__49486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RX_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__12697 (
            .O(N__49469),
            .I(N__49464));
    InMux I__12696 (
            .O(N__49468),
            .I(N__49461));
    InMux I__12695 (
            .O(N__49467),
            .I(N__49457));
    LocalMux I__12694 (
            .O(N__49464),
            .I(N__49454));
    LocalMux I__12693 (
            .O(N__49461),
            .I(N__49451));
    InMux I__12692 (
            .O(N__49460),
            .I(N__49447));
    LocalMux I__12691 (
            .O(N__49457),
            .I(N__49444));
    Span4Mux_h I__12690 (
            .O(N__49454),
            .I(N__49438));
    Span4Mux_h I__12689 (
            .O(N__49451),
            .I(N__49435));
    InMux I__12688 (
            .O(N__49450),
            .I(N__49432));
    LocalMux I__12687 (
            .O(N__49447),
            .I(N__49429));
    Span4Mux_v I__12686 (
            .O(N__49444),
            .I(N__49426));
    InMux I__12685 (
            .O(N__49443),
            .I(N__49423));
    InMux I__12684 (
            .O(N__49442),
            .I(N__49420));
    InMux I__12683 (
            .O(N__49441),
            .I(N__49417));
    Sp12to4 I__12682 (
            .O(N__49438),
            .I(N__49410));
    Sp12to4 I__12681 (
            .O(N__49435),
            .I(N__49410));
    LocalMux I__12680 (
            .O(N__49432),
            .I(N__49410));
    Span4Mux_h I__12679 (
            .O(N__49429),
            .I(N__49407));
    Span4Mux_h I__12678 (
            .O(N__49426),
            .I(N__49402));
    LocalMux I__12677 (
            .O(N__49423),
            .I(N__49402));
    LocalMux I__12676 (
            .O(N__49420),
            .I(N__49397));
    LocalMux I__12675 (
            .O(N__49417),
            .I(N__49397));
    Odrv12 I__12674 (
            .O(N__49410),
            .I(\ALU.un9_addsub_cry_2_c_RNIMN63NZ0 ));
    Odrv4 I__12673 (
            .O(N__49407),
            .I(\ALU.un9_addsub_cry_2_c_RNIMN63NZ0 ));
    Odrv4 I__12672 (
            .O(N__49402),
            .I(\ALU.un9_addsub_cry_2_c_RNIMN63NZ0 ));
    Odrv4 I__12671 (
            .O(N__49397),
            .I(\ALU.un9_addsub_cry_2_c_RNIMN63NZ0 ));
    InMux I__12670 (
            .O(N__49388),
            .I(N__49384));
    InMux I__12669 (
            .O(N__49387),
            .I(N__49379));
    LocalMux I__12668 (
            .O(N__49384),
            .I(N__49375));
    InMux I__12667 (
            .O(N__49383),
            .I(N__49372));
    InMux I__12666 (
            .O(N__49382),
            .I(N__49369));
    LocalMux I__12665 (
            .O(N__49379),
            .I(N__49365));
    InMux I__12664 (
            .O(N__49378),
            .I(N__49362));
    Sp12to4 I__12663 (
            .O(N__49375),
            .I(N__49355));
    LocalMux I__12662 (
            .O(N__49372),
            .I(N__49355));
    LocalMux I__12661 (
            .O(N__49369),
            .I(N__49352));
    InMux I__12660 (
            .O(N__49368),
            .I(N__49349));
    Span4Mux_h I__12659 (
            .O(N__49365),
            .I(N__49346));
    LocalMux I__12658 (
            .O(N__49362),
            .I(N__49343));
    InMux I__12657 (
            .O(N__49361),
            .I(N__49340));
    InMux I__12656 (
            .O(N__49360),
            .I(N__49337));
    Span12Mux_v I__12655 (
            .O(N__49355),
            .I(N__49334));
    Span4Mux_h I__12654 (
            .O(N__49352),
            .I(N__49331));
    LocalMux I__12653 (
            .O(N__49349),
            .I(N__49328));
    Span4Mux_h I__12652 (
            .O(N__49346),
            .I(N__49319));
    Span4Mux_v I__12651 (
            .O(N__49343),
            .I(N__49319));
    LocalMux I__12650 (
            .O(N__49340),
            .I(N__49319));
    LocalMux I__12649 (
            .O(N__49337),
            .I(N__49319));
    Odrv12 I__12648 (
            .O(N__49334),
            .I(\ALU.d_RNIE8SJN5Z0Z_3 ));
    Odrv4 I__12647 (
            .O(N__49331),
            .I(\ALU.d_RNIE8SJN5Z0Z_3 ));
    Odrv4 I__12646 (
            .O(N__49328),
            .I(\ALU.d_RNIE8SJN5Z0Z_3 ));
    Odrv4 I__12645 (
            .O(N__49319),
            .I(\ALU.d_RNIE8SJN5Z0Z_3 ));
    InMux I__12644 (
            .O(N__49310),
            .I(N__49307));
    LocalMux I__12643 (
            .O(N__49307),
            .I(N__49304));
    Span4Mux_h I__12642 (
            .O(N__49304),
            .I(N__49300));
    InMux I__12641 (
            .O(N__49303),
            .I(N__49297));
    Span4Mux_h I__12640 (
            .O(N__49300),
            .I(N__49294));
    LocalMux I__12639 (
            .O(N__49297),
            .I(\ALU.bZ0Z_3 ));
    Odrv4 I__12638 (
            .O(N__49294),
            .I(\ALU.bZ0Z_3 ));
    InMux I__12637 (
            .O(N__49289),
            .I(N__49282));
    InMux I__12636 (
            .O(N__49288),
            .I(N__49278));
    InMux I__12635 (
            .O(N__49287),
            .I(N__49275));
    InMux I__12634 (
            .O(N__49286),
            .I(N__49272));
    InMux I__12633 (
            .O(N__49285),
            .I(N__49269));
    LocalMux I__12632 (
            .O(N__49282),
            .I(N__49266));
    InMux I__12631 (
            .O(N__49281),
            .I(N__49263));
    LocalMux I__12630 (
            .O(N__49278),
            .I(N__49259));
    LocalMux I__12629 (
            .O(N__49275),
            .I(N__49248));
    LocalMux I__12628 (
            .O(N__49272),
            .I(N__49248));
    LocalMux I__12627 (
            .O(N__49269),
            .I(N__49248));
    Span4Mux_h I__12626 (
            .O(N__49266),
            .I(N__49248));
    LocalMux I__12625 (
            .O(N__49263),
            .I(N__49248));
    InMux I__12624 (
            .O(N__49262),
            .I(N__49245));
    Span4Mux_h I__12623 (
            .O(N__49259),
            .I(N__49241));
    Span4Mux_v I__12622 (
            .O(N__49248),
            .I(N__49236));
    LocalMux I__12621 (
            .O(N__49245),
            .I(N__49236));
    InMux I__12620 (
            .O(N__49244),
            .I(N__49233));
    Span4Mux_v I__12619 (
            .O(N__49241),
            .I(N__49230));
    Span4Mux_h I__12618 (
            .O(N__49236),
            .I(N__49225));
    LocalMux I__12617 (
            .O(N__49233),
            .I(N__49225));
    Odrv4 I__12616 (
            .O(N__49230),
            .I(\ALU.un9_addsub_cry_3_c_RNI4L7ROZ0 ));
    Odrv4 I__12615 (
            .O(N__49225),
            .I(\ALU.un9_addsub_cry_3_c_RNI4L7ROZ0 ));
    InMux I__12614 (
            .O(N__49220),
            .I(N__49214));
    InMux I__12613 (
            .O(N__49219),
            .I(N__49208));
    InMux I__12612 (
            .O(N__49218),
            .I(N__49205));
    InMux I__12611 (
            .O(N__49217),
            .I(N__49201));
    LocalMux I__12610 (
            .O(N__49214),
            .I(N__49198));
    InMux I__12609 (
            .O(N__49213),
            .I(N__49195));
    InMux I__12608 (
            .O(N__49212),
            .I(N__49192));
    InMux I__12607 (
            .O(N__49211),
            .I(N__49189));
    LocalMux I__12606 (
            .O(N__49208),
            .I(N__49184));
    LocalMux I__12605 (
            .O(N__49205),
            .I(N__49184));
    InMux I__12604 (
            .O(N__49204),
            .I(N__49181));
    LocalMux I__12603 (
            .O(N__49201),
            .I(N__49178));
    Span4Mux_h I__12602 (
            .O(N__49198),
            .I(N__49173));
    LocalMux I__12601 (
            .O(N__49195),
            .I(N__49173));
    LocalMux I__12600 (
            .O(N__49192),
            .I(N__49170));
    LocalMux I__12599 (
            .O(N__49189),
            .I(N__49167));
    Span4Mux_v I__12598 (
            .O(N__49184),
            .I(N__49162));
    LocalMux I__12597 (
            .O(N__49181),
            .I(N__49162));
    Odrv12 I__12596 (
            .O(N__49178),
            .I(\ALU.d_RNIMA3938Z0Z_4 ));
    Odrv4 I__12595 (
            .O(N__49173),
            .I(\ALU.d_RNIMA3938Z0Z_4 ));
    Odrv4 I__12594 (
            .O(N__49170),
            .I(\ALU.d_RNIMA3938Z0Z_4 ));
    Odrv4 I__12593 (
            .O(N__49167),
            .I(\ALU.d_RNIMA3938Z0Z_4 ));
    Odrv4 I__12592 (
            .O(N__49162),
            .I(\ALU.d_RNIMA3938Z0Z_4 ));
    InMux I__12591 (
            .O(N__49151),
            .I(N__49148));
    LocalMux I__12590 (
            .O(N__49148),
            .I(N__49145));
    Span4Mux_v I__12589 (
            .O(N__49145),
            .I(N__49141));
    InMux I__12588 (
            .O(N__49144),
            .I(N__49138));
    Span4Mux_h I__12587 (
            .O(N__49141),
            .I(N__49133));
    LocalMux I__12586 (
            .O(N__49138),
            .I(N__49133));
    Odrv4 I__12585 (
            .O(N__49133),
            .I(\ALU.bZ0Z_4 ));
    InMux I__12584 (
            .O(N__49130),
            .I(N__49127));
    LocalMux I__12583 (
            .O(N__49127),
            .I(N__49124));
    Span4Mux_h I__12582 (
            .O(N__49124),
            .I(N__49119));
    InMux I__12581 (
            .O(N__49123),
            .I(N__49116));
    InMux I__12580 (
            .O(N__49122),
            .I(N__49113));
    Span4Mux_h I__12579 (
            .O(N__49119),
            .I(N__49105));
    LocalMux I__12578 (
            .O(N__49116),
            .I(N__49105));
    LocalMux I__12577 (
            .O(N__49113),
            .I(N__49105));
    InMux I__12576 (
            .O(N__49112),
            .I(N__49102));
    Span4Mux_v I__12575 (
            .O(N__49105),
            .I(N__49098));
    LocalMux I__12574 (
            .O(N__49102),
            .I(N__49095));
    InMux I__12573 (
            .O(N__49101),
            .I(N__49091));
    Span4Mux_h I__12572 (
            .O(N__49098),
            .I(N__49086));
    Span4Mux_v I__12571 (
            .O(N__49095),
            .I(N__49083));
    InMux I__12570 (
            .O(N__49094),
            .I(N__49080));
    LocalMux I__12569 (
            .O(N__49091),
            .I(N__49077));
    InMux I__12568 (
            .O(N__49090),
            .I(N__49074));
    InMux I__12567 (
            .O(N__49089),
            .I(N__49071));
    Sp12to4 I__12566 (
            .O(N__49086),
            .I(N__49068));
    Span4Mux_h I__12565 (
            .O(N__49083),
            .I(N__49063));
    LocalMux I__12564 (
            .O(N__49080),
            .I(N__49063));
    Span4Mux_h I__12563 (
            .O(N__49077),
            .I(N__49056));
    LocalMux I__12562 (
            .O(N__49074),
            .I(N__49056));
    LocalMux I__12561 (
            .O(N__49071),
            .I(N__49056));
    Odrv12 I__12560 (
            .O(N__49068),
            .I(\ALU.un9_addsub_cry_4_c_RNIUEDLMZ0 ));
    Odrv4 I__12559 (
            .O(N__49063),
            .I(\ALU.un9_addsub_cry_4_c_RNIUEDLMZ0 ));
    Odrv4 I__12558 (
            .O(N__49056),
            .I(\ALU.un9_addsub_cry_4_c_RNIUEDLMZ0 ));
    InMux I__12557 (
            .O(N__49049),
            .I(N__49040));
    InMux I__12556 (
            .O(N__49048),
            .I(N__49037));
    InMux I__12555 (
            .O(N__49047),
            .I(N__49034));
    InMux I__12554 (
            .O(N__49046),
            .I(N__49031));
    InMux I__12553 (
            .O(N__49045),
            .I(N__49028));
    InMux I__12552 (
            .O(N__49044),
            .I(N__49024));
    InMux I__12551 (
            .O(N__49043),
            .I(N__49021));
    LocalMux I__12550 (
            .O(N__49040),
            .I(N__49018));
    LocalMux I__12549 (
            .O(N__49037),
            .I(N__49013));
    LocalMux I__12548 (
            .O(N__49034),
            .I(N__49013));
    LocalMux I__12547 (
            .O(N__49031),
            .I(N__49010));
    LocalMux I__12546 (
            .O(N__49028),
            .I(N__49007));
    InMux I__12545 (
            .O(N__49027),
            .I(N__49004));
    LocalMux I__12544 (
            .O(N__49024),
            .I(N__48999));
    LocalMux I__12543 (
            .O(N__49021),
            .I(N__48999));
    Span4Mux_v I__12542 (
            .O(N__49018),
            .I(N__48996));
    Span4Mux_v I__12541 (
            .O(N__49013),
            .I(N__48991));
    Span4Mux_h I__12540 (
            .O(N__49010),
            .I(N__48991));
    Span4Mux_v I__12539 (
            .O(N__49007),
            .I(N__48986));
    LocalMux I__12538 (
            .O(N__49004),
            .I(N__48986));
    Span4Mux_v I__12537 (
            .O(N__48999),
            .I(N__48983));
    Span4Mux_h I__12536 (
            .O(N__48996),
            .I(N__48976));
    Span4Mux_v I__12535 (
            .O(N__48991),
            .I(N__48976));
    Span4Mux_v I__12534 (
            .O(N__48986),
            .I(N__48976));
    Span4Mux_v I__12533 (
            .O(N__48983),
            .I(N__48973));
    Span4Mux_v I__12532 (
            .O(N__48976),
            .I(N__48970));
    Odrv4 I__12531 (
            .O(N__48973),
            .I(\ALU.d_RNIH1NE6FZ0Z_5 ));
    Odrv4 I__12530 (
            .O(N__48970),
            .I(\ALU.d_RNIH1NE6FZ0Z_5 ));
    InMux I__12529 (
            .O(N__48965),
            .I(N__48961));
    InMux I__12528 (
            .O(N__48964),
            .I(N__48958));
    LocalMux I__12527 (
            .O(N__48961),
            .I(N__48955));
    LocalMux I__12526 (
            .O(N__48958),
            .I(N__48950));
    Span4Mux_h I__12525 (
            .O(N__48955),
            .I(N__48950));
    Odrv4 I__12524 (
            .O(N__48950),
            .I(\ALU.bZ0Z_5 ));
    InMux I__12523 (
            .O(N__48947),
            .I(N__48944));
    LocalMux I__12522 (
            .O(N__48944),
            .I(N__48939));
    InMux I__12521 (
            .O(N__48943),
            .I(N__48936));
    InMux I__12520 (
            .O(N__48942),
            .I(N__48933));
    Span4Mux_v I__12519 (
            .O(N__48939),
            .I(N__48924));
    LocalMux I__12518 (
            .O(N__48936),
            .I(N__48924));
    LocalMux I__12517 (
            .O(N__48933),
            .I(N__48924));
    InMux I__12516 (
            .O(N__48932),
            .I(N__48921));
    InMux I__12515 (
            .O(N__48931),
            .I(N__48918));
    Span4Mux_v I__12514 (
            .O(N__48924),
            .I(N__48909));
    LocalMux I__12513 (
            .O(N__48921),
            .I(N__48909));
    LocalMux I__12512 (
            .O(N__48918),
            .I(N__48909));
    InMux I__12511 (
            .O(N__48917),
            .I(N__48906));
    InMux I__12510 (
            .O(N__48916),
            .I(N__48903));
    Span4Mux_h I__12509 (
            .O(N__48909),
            .I(N__48896));
    LocalMux I__12508 (
            .O(N__48906),
            .I(N__48896));
    LocalMux I__12507 (
            .O(N__48903),
            .I(N__48896));
    Odrv4 I__12506 (
            .O(N__48896),
            .I(\ALU.d_RNILPR7TQZ0Z_6 ));
    InMux I__12505 (
            .O(N__48893),
            .I(N__48888));
    InMux I__12504 (
            .O(N__48892),
            .I(N__48885));
    InMux I__12503 (
            .O(N__48891),
            .I(N__48882));
    LocalMux I__12502 (
            .O(N__48888),
            .I(N__48877));
    LocalMux I__12501 (
            .O(N__48885),
            .I(N__48874));
    LocalMux I__12500 (
            .O(N__48882),
            .I(N__48871));
    InMux I__12499 (
            .O(N__48881),
            .I(N__48868));
    InMux I__12498 (
            .O(N__48880),
            .I(N__48864));
    Span4Mux_h I__12497 (
            .O(N__48877),
            .I(N__48860));
    Span4Mux_h I__12496 (
            .O(N__48874),
            .I(N__48857));
    Span4Mux_v I__12495 (
            .O(N__48871),
            .I(N__48851));
    LocalMux I__12494 (
            .O(N__48868),
            .I(N__48851));
    InMux I__12493 (
            .O(N__48867),
            .I(N__48848));
    LocalMux I__12492 (
            .O(N__48864),
            .I(N__48845));
    InMux I__12491 (
            .O(N__48863),
            .I(N__48842));
    Span4Mux_v I__12490 (
            .O(N__48860),
            .I(N__48839));
    Span4Mux_v I__12489 (
            .O(N__48857),
            .I(N__48836));
    InMux I__12488 (
            .O(N__48856),
            .I(N__48833));
    Span4Mux_h I__12487 (
            .O(N__48851),
            .I(N__48824));
    LocalMux I__12486 (
            .O(N__48848),
            .I(N__48824));
    Span4Mux_h I__12485 (
            .O(N__48845),
            .I(N__48824));
    LocalMux I__12484 (
            .O(N__48842),
            .I(N__48824));
    Odrv4 I__12483 (
            .O(N__48839),
            .I(\ALU.un9_addsub_cry_5_c_RNI26HCNZ0 ));
    Odrv4 I__12482 (
            .O(N__48836),
            .I(\ALU.un9_addsub_cry_5_c_RNI26HCNZ0 ));
    LocalMux I__12481 (
            .O(N__48833),
            .I(\ALU.un9_addsub_cry_5_c_RNI26HCNZ0 ));
    Odrv4 I__12480 (
            .O(N__48824),
            .I(\ALU.un9_addsub_cry_5_c_RNI26HCNZ0 ));
    InMux I__12479 (
            .O(N__48815),
            .I(N__48812));
    LocalMux I__12478 (
            .O(N__48812),
            .I(N__48808));
    InMux I__12477 (
            .O(N__48811),
            .I(N__48805));
    Span4Mux_h I__12476 (
            .O(N__48808),
            .I(N__48802));
    LocalMux I__12475 (
            .O(N__48805),
            .I(N__48799));
    Span4Mux_h I__12474 (
            .O(N__48802),
            .I(N__48796));
    Odrv12 I__12473 (
            .O(N__48799),
            .I(\ALU.bZ0Z_6 ));
    Odrv4 I__12472 (
            .O(N__48796),
            .I(\ALU.bZ0Z_6 ));
    InMux I__12471 (
            .O(N__48791),
            .I(N__48784));
    InMux I__12470 (
            .O(N__48790),
            .I(N__48781));
    InMux I__12469 (
            .O(N__48789),
            .I(N__48778));
    InMux I__12468 (
            .O(N__48788),
            .I(N__48774));
    InMux I__12467 (
            .O(N__48787),
            .I(N__48771));
    LocalMux I__12466 (
            .O(N__48784),
            .I(N__48765));
    LocalMux I__12465 (
            .O(N__48781),
            .I(N__48765));
    LocalMux I__12464 (
            .O(N__48778),
            .I(N__48762));
    InMux I__12463 (
            .O(N__48777),
            .I(N__48759));
    LocalMux I__12462 (
            .O(N__48774),
            .I(N__48756));
    LocalMux I__12461 (
            .O(N__48771),
            .I(N__48753));
    InMux I__12460 (
            .O(N__48770),
            .I(N__48750));
    Span4Mux_h I__12459 (
            .O(N__48765),
            .I(N__48742));
    Span4Mux_h I__12458 (
            .O(N__48762),
            .I(N__48742));
    LocalMux I__12457 (
            .O(N__48759),
            .I(N__48742));
    Span4Mux_v I__12456 (
            .O(N__48756),
            .I(N__48735));
    Span4Mux_v I__12455 (
            .O(N__48753),
            .I(N__48735));
    LocalMux I__12454 (
            .O(N__48750),
            .I(N__48735));
    InMux I__12453 (
            .O(N__48749),
            .I(N__48732));
    Span4Mux_h I__12452 (
            .O(N__48742),
            .I(N__48729));
    Span4Mux_h I__12451 (
            .O(N__48735),
            .I(N__48726));
    LocalMux I__12450 (
            .O(N__48732),
            .I(N__48723));
    Odrv4 I__12449 (
            .O(N__48729),
            .I(\ALU.un9_addsub_cry_6_c_RNIUKMKRZ0 ));
    Odrv4 I__12448 (
            .O(N__48726),
            .I(\ALU.un9_addsub_cry_6_c_RNIUKMKRZ0 ));
    Odrv12 I__12447 (
            .O(N__48723),
            .I(\ALU.un9_addsub_cry_6_c_RNIUKMKRZ0 ));
    InMux I__12446 (
            .O(N__48716),
            .I(N__48710));
    InMux I__12445 (
            .O(N__48715),
            .I(N__48707));
    InMux I__12444 (
            .O(N__48714),
            .I(N__48704));
    InMux I__12443 (
            .O(N__48713),
            .I(N__48701));
    LocalMux I__12442 (
            .O(N__48710),
            .I(N__48697));
    LocalMux I__12441 (
            .O(N__48707),
            .I(N__48688));
    LocalMux I__12440 (
            .O(N__48704),
            .I(N__48688));
    LocalMux I__12439 (
            .O(N__48701),
            .I(N__48688));
    InMux I__12438 (
            .O(N__48700),
            .I(N__48685));
    Span4Mux_h I__12437 (
            .O(N__48697),
            .I(N__48681));
    InMux I__12436 (
            .O(N__48696),
            .I(N__48678));
    InMux I__12435 (
            .O(N__48695),
            .I(N__48675));
    Span4Mux_v I__12434 (
            .O(N__48688),
            .I(N__48670));
    LocalMux I__12433 (
            .O(N__48685),
            .I(N__48670));
    InMux I__12432 (
            .O(N__48684),
            .I(N__48667));
    Odrv4 I__12431 (
            .O(N__48681),
            .I(\ALU.d_RNIIIPM081Z0Z_7 ));
    LocalMux I__12430 (
            .O(N__48678),
            .I(\ALU.d_RNIIIPM081Z0Z_7 ));
    LocalMux I__12429 (
            .O(N__48675),
            .I(\ALU.d_RNIIIPM081Z0Z_7 ));
    Odrv4 I__12428 (
            .O(N__48670),
            .I(\ALU.d_RNIIIPM081Z0Z_7 ));
    LocalMux I__12427 (
            .O(N__48667),
            .I(\ALU.d_RNIIIPM081Z0Z_7 ));
    InMux I__12426 (
            .O(N__48656),
            .I(N__48650));
    InMux I__12425 (
            .O(N__48655),
            .I(N__48650));
    LocalMux I__12424 (
            .O(N__48650),
            .I(N__48647));
    Span4Mux_h I__12423 (
            .O(N__48647),
            .I(N__48644));
    Odrv4 I__12422 (
            .O(N__48644),
            .I(\ALU.bZ0Z_7 ));
    InMux I__12421 (
            .O(N__48641),
            .I(N__48606));
    InMux I__12420 (
            .O(N__48640),
            .I(N__48606));
    InMux I__12419 (
            .O(N__48639),
            .I(N__48606));
    InMux I__12418 (
            .O(N__48638),
            .I(N__48606));
    InMux I__12417 (
            .O(N__48637),
            .I(N__48599));
    InMux I__12416 (
            .O(N__48636),
            .I(N__48599));
    InMux I__12415 (
            .O(N__48635),
            .I(N__48599));
    CascadeMux I__12414 (
            .O(N__48634),
            .I(N__48557));
    InMux I__12413 (
            .O(N__48633),
            .I(N__48548));
    InMux I__12412 (
            .O(N__48632),
            .I(N__48548));
    InMux I__12411 (
            .O(N__48631),
            .I(N__48548));
    InMux I__12410 (
            .O(N__48630),
            .I(N__48545));
    InMux I__12409 (
            .O(N__48629),
            .I(N__48542));
    InMux I__12408 (
            .O(N__48628),
            .I(N__48535));
    InMux I__12407 (
            .O(N__48627),
            .I(N__48535));
    InMux I__12406 (
            .O(N__48626),
            .I(N__48535));
    InMux I__12405 (
            .O(N__48625),
            .I(N__48526));
    InMux I__12404 (
            .O(N__48624),
            .I(N__48526));
    InMux I__12403 (
            .O(N__48623),
            .I(N__48526));
    InMux I__12402 (
            .O(N__48622),
            .I(N__48526));
    InMux I__12401 (
            .O(N__48621),
            .I(N__48517));
    InMux I__12400 (
            .O(N__48620),
            .I(N__48517));
    InMux I__12399 (
            .O(N__48619),
            .I(N__48517));
    InMux I__12398 (
            .O(N__48618),
            .I(N__48517));
    InMux I__12397 (
            .O(N__48617),
            .I(N__48510));
    InMux I__12396 (
            .O(N__48616),
            .I(N__48510));
    InMux I__12395 (
            .O(N__48615),
            .I(N__48510));
    LocalMux I__12394 (
            .O(N__48606),
            .I(N__48504));
    LocalMux I__12393 (
            .O(N__48599),
            .I(N__48504));
    InMux I__12392 (
            .O(N__48598),
            .I(N__48501));
    InMux I__12391 (
            .O(N__48597),
            .I(N__48498));
    InMux I__12390 (
            .O(N__48596),
            .I(N__48472));
    InMux I__12389 (
            .O(N__48595),
            .I(N__48472));
    InMux I__12388 (
            .O(N__48594),
            .I(N__48472));
    InMux I__12387 (
            .O(N__48593),
            .I(N__48472));
    InMux I__12386 (
            .O(N__48592),
            .I(N__48472));
    InMux I__12385 (
            .O(N__48591),
            .I(N__48469));
    InMux I__12384 (
            .O(N__48590),
            .I(N__48464));
    InMux I__12383 (
            .O(N__48589),
            .I(N__48464));
    InMux I__12382 (
            .O(N__48588),
            .I(N__48461));
    InMux I__12381 (
            .O(N__48587),
            .I(N__48454));
    InMux I__12380 (
            .O(N__48586),
            .I(N__48454));
    InMux I__12379 (
            .O(N__48585),
            .I(N__48454));
    InMux I__12378 (
            .O(N__48584),
            .I(N__48447));
    InMux I__12377 (
            .O(N__48583),
            .I(N__48447));
    InMux I__12376 (
            .O(N__48582),
            .I(N__48447));
    InMux I__12375 (
            .O(N__48581),
            .I(N__48444));
    InMux I__12374 (
            .O(N__48580),
            .I(N__48437));
    InMux I__12373 (
            .O(N__48579),
            .I(N__48437));
    InMux I__12372 (
            .O(N__48578),
            .I(N__48437));
    InMux I__12371 (
            .O(N__48577),
            .I(N__48427));
    CascadeMux I__12370 (
            .O(N__48576),
            .I(N__48416));
    CascadeMux I__12369 (
            .O(N__48575),
            .I(N__48413));
    InMux I__12368 (
            .O(N__48574),
            .I(N__48406));
    InMux I__12367 (
            .O(N__48573),
            .I(N__48401));
    InMux I__12366 (
            .O(N__48572),
            .I(N__48401));
    InMux I__12365 (
            .O(N__48571),
            .I(N__48396));
    InMux I__12364 (
            .O(N__48570),
            .I(N__48396));
    InMux I__12363 (
            .O(N__48569),
            .I(N__48389));
    InMux I__12362 (
            .O(N__48568),
            .I(N__48389));
    InMux I__12361 (
            .O(N__48567),
            .I(N__48389));
    InMux I__12360 (
            .O(N__48566),
            .I(N__48384));
    InMux I__12359 (
            .O(N__48565),
            .I(N__48384));
    InMux I__12358 (
            .O(N__48564),
            .I(N__48375));
    InMux I__12357 (
            .O(N__48563),
            .I(N__48375));
    InMux I__12356 (
            .O(N__48562),
            .I(N__48375));
    InMux I__12355 (
            .O(N__48561),
            .I(N__48375));
    InMux I__12354 (
            .O(N__48560),
            .I(N__48366));
    InMux I__12353 (
            .O(N__48557),
            .I(N__48366));
    InMux I__12352 (
            .O(N__48556),
            .I(N__48366));
    InMux I__12351 (
            .O(N__48555),
            .I(N__48366));
    LocalMux I__12350 (
            .O(N__48548),
            .I(N__48363));
    LocalMux I__12349 (
            .O(N__48545),
            .I(N__48354));
    LocalMux I__12348 (
            .O(N__48542),
            .I(N__48354));
    LocalMux I__12347 (
            .O(N__48535),
            .I(N__48354));
    LocalMux I__12346 (
            .O(N__48526),
            .I(N__48354));
    LocalMux I__12345 (
            .O(N__48517),
            .I(N__48349));
    LocalMux I__12344 (
            .O(N__48510),
            .I(N__48349));
    InMux I__12343 (
            .O(N__48509),
            .I(N__48341));
    Span4Mux_h I__12342 (
            .O(N__48504),
            .I(N__48334));
    LocalMux I__12341 (
            .O(N__48501),
            .I(N__48334));
    LocalMux I__12340 (
            .O(N__48498),
            .I(N__48331));
    InMux I__12339 (
            .O(N__48497),
            .I(N__48317));
    InMux I__12338 (
            .O(N__48496),
            .I(N__48317));
    InMux I__12337 (
            .O(N__48495),
            .I(N__48317));
    InMux I__12336 (
            .O(N__48494),
            .I(N__48317));
    InMux I__12335 (
            .O(N__48493),
            .I(N__48317));
    InMux I__12334 (
            .O(N__48492),
            .I(N__48310));
    InMux I__12333 (
            .O(N__48491),
            .I(N__48310));
    InMux I__12332 (
            .O(N__48490),
            .I(N__48310));
    InMux I__12331 (
            .O(N__48489),
            .I(N__48301));
    InMux I__12330 (
            .O(N__48488),
            .I(N__48301));
    InMux I__12329 (
            .O(N__48487),
            .I(N__48301));
    InMux I__12328 (
            .O(N__48486),
            .I(N__48301));
    InMux I__12327 (
            .O(N__48485),
            .I(N__48294));
    InMux I__12326 (
            .O(N__48484),
            .I(N__48294));
    InMux I__12325 (
            .O(N__48483),
            .I(N__48294));
    LocalMux I__12324 (
            .O(N__48472),
            .I(N__48291));
    LocalMux I__12323 (
            .O(N__48469),
            .I(N__48284));
    LocalMux I__12322 (
            .O(N__48464),
            .I(N__48284));
    LocalMux I__12321 (
            .O(N__48461),
            .I(N__48284));
    LocalMux I__12320 (
            .O(N__48454),
            .I(N__48275));
    LocalMux I__12319 (
            .O(N__48447),
            .I(N__48275));
    LocalMux I__12318 (
            .O(N__48444),
            .I(N__48275));
    LocalMux I__12317 (
            .O(N__48437),
            .I(N__48275));
    InMux I__12316 (
            .O(N__48436),
            .I(N__48262));
    InMux I__12315 (
            .O(N__48435),
            .I(N__48258));
    InMux I__12314 (
            .O(N__48434),
            .I(N__48255));
    InMux I__12313 (
            .O(N__48433),
            .I(N__48252));
    InMux I__12312 (
            .O(N__48432),
            .I(N__48244));
    InMux I__12311 (
            .O(N__48431),
            .I(N__48244));
    InMux I__12310 (
            .O(N__48430),
            .I(N__48244));
    LocalMux I__12309 (
            .O(N__48427),
            .I(N__48241));
    InMux I__12308 (
            .O(N__48426),
            .I(N__48238));
    InMux I__12307 (
            .O(N__48425),
            .I(N__48227));
    InMux I__12306 (
            .O(N__48424),
            .I(N__48227));
    InMux I__12305 (
            .O(N__48423),
            .I(N__48227));
    InMux I__12304 (
            .O(N__48422),
            .I(N__48227));
    InMux I__12303 (
            .O(N__48421),
            .I(N__48227));
    InMux I__12302 (
            .O(N__48420),
            .I(N__48222));
    InMux I__12301 (
            .O(N__48419),
            .I(N__48222));
    InMux I__12300 (
            .O(N__48416),
            .I(N__48215));
    InMux I__12299 (
            .O(N__48413),
            .I(N__48215));
    InMux I__12298 (
            .O(N__48412),
            .I(N__48215));
    InMux I__12297 (
            .O(N__48411),
            .I(N__48208));
    InMux I__12296 (
            .O(N__48410),
            .I(N__48208));
    InMux I__12295 (
            .O(N__48409),
            .I(N__48208));
    LocalMux I__12294 (
            .O(N__48406),
            .I(N__48203));
    LocalMux I__12293 (
            .O(N__48401),
            .I(N__48203));
    LocalMux I__12292 (
            .O(N__48396),
            .I(N__48186));
    LocalMux I__12291 (
            .O(N__48389),
            .I(N__48186));
    LocalMux I__12290 (
            .O(N__48384),
            .I(N__48186));
    LocalMux I__12289 (
            .O(N__48375),
            .I(N__48186));
    LocalMux I__12288 (
            .O(N__48366),
            .I(N__48186));
    Span4Mux_v I__12287 (
            .O(N__48363),
            .I(N__48186));
    Span4Mux_v I__12286 (
            .O(N__48354),
            .I(N__48186));
    Span4Mux_h I__12285 (
            .O(N__48349),
            .I(N__48186));
    InMux I__12284 (
            .O(N__48348),
            .I(N__48183));
    InMux I__12283 (
            .O(N__48347),
            .I(N__48174));
    InMux I__12282 (
            .O(N__48346),
            .I(N__48174));
    InMux I__12281 (
            .O(N__48345),
            .I(N__48174));
    InMux I__12280 (
            .O(N__48344),
            .I(N__48174));
    LocalMux I__12279 (
            .O(N__48341),
            .I(N__48171));
    InMux I__12278 (
            .O(N__48340),
            .I(N__48166));
    InMux I__12277 (
            .O(N__48339),
            .I(N__48166));
    Span4Mux_h I__12276 (
            .O(N__48334),
            .I(N__48161));
    Span4Mux_v I__12275 (
            .O(N__48331),
            .I(N__48161));
    InMux I__12274 (
            .O(N__48330),
            .I(N__48156));
    InMux I__12273 (
            .O(N__48329),
            .I(N__48156));
    InMux I__12272 (
            .O(N__48328),
            .I(N__48153));
    LocalMux I__12271 (
            .O(N__48317),
            .I(N__48146));
    LocalMux I__12270 (
            .O(N__48310),
            .I(N__48146));
    LocalMux I__12269 (
            .O(N__48301),
            .I(N__48146));
    LocalMux I__12268 (
            .O(N__48294),
            .I(N__48137));
    Span4Mux_h I__12267 (
            .O(N__48291),
            .I(N__48137));
    Span4Mux_v I__12266 (
            .O(N__48284),
            .I(N__48137));
    Span4Mux_h I__12265 (
            .O(N__48275),
            .I(N__48137));
    InMux I__12264 (
            .O(N__48274),
            .I(N__48132));
    InMux I__12263 (
            .O(N__48273),
            .I(N__48132));
    InMux I__12262 (
            .O(N__48272),
            .I(N__48127));
    InMux I__12261 (
            .O(N__48271),
            .I(N__48127));
    InMux I__12260 (
            .O(N__48270),
            .I(N__48122));
    InMux I__12259 (
            .O(N__48269),
            .I(N__48122));
    InMux I__12258 (
            .O(N__48268),
            .I(N__48113));
    InMux I__12257 (
            .O(N__48267),
            .I(N__48113));
    InMux I__12256 (
            .O(N__48266),
            .I(N__48113));
    InMux I__12255 (
            .O(N__48265),
            .I(N__48113));
    LocalMux I__12254 (
            .O(N__48262),
            .I(N__48110));
    InMux I__12253 (
            .O(N__48261),
            .I(N__48106));
    LocalMux I__12252 (
            .O(N__48258),
            .I(N__48100));
    LocalMux I__12251 (
            .O(N__48255),
            .I(N__48100));
    LocalMux I__12250 (
            .O(N__48252),
            .I(N__48097));
    InMux I__12249 (
            .O(N__48251),
            .I(N__48089));
    LocalMux I__12248 (
            .O(N__48244),
            .I(N__48078));
    Span4Mux_h I__12247 (
            .O(N__48241),
            .I(N__48078));
    LocalMux I__12246 (
            .O(N__48238),
            .I(N__48078));
    LocalMux I__12245 (
            .O(N__48227),
            .I(N__48078));
    LocalMux I__12244 (
            .O(N__48222),
            .I(N__48078));
    LocalMux I__12243 (
            .O(N__48215),
            .I(N__48065));
    LocalMux I__12242 (
            .O(N__48208),
            .I(N__48065));
    Span4Mux_v I__12241 (
            .O(N__48203),
            .I(N__48065));
    Span4Mux_v I__12240 (
            .O(N__48186),
            .I(N__48065));
    LocalMux I__12239 (
            .O(N__48183),
            .I(N__48060));
    LocalMux I__12238 (
            .O(N__48174),
            .I(N__48060));
    Span4Mux_h I__12237 (
            .O(N__48171),
            .I(N__48055));
    LocalMux I__12236 (
            .O(N__48166),
            .I(N__48055));
    Span4Mux_v I__12235 (
            .O(N__48161),
            .I(N__48049));
    LocalMux I__12234 (
            .O(N__48156),
            .I(N__48049));
    LocalMux I__12233 (
            .O(N__48153),
            .I(N__48034));
    Span4Mux_v I__12232 (
            .O(N__48146),
            .I(N__48034));
    Span4Mux_v I__12231 (
            .O(N__48137),
            .I(N__48034));
    LocalMux I__12230 (
            .O(N__48132),
            .I(N__48034));
    LocalMux I__12229 (
            .O(N__48127),
            .I(N__48034));
    LocalMux I__12228 (
            .O(N__48122),
            .I(N__48034));
    LocalMux I__12227 (
            .O(N__48113),
            .I(N__48034));
    Span4Mux_h I__12226 (
            .O(N__48110),
            .I(N__48031));
    InMux I__12225 (
            .O(N__48109),
            .I(N__48026));
    LocalMux I__12224 (
            .O(N__48106),
            .I(N__48023));
    InMux I__12223 (
            .O(N__48105),
            .I(N__48020));
    Span4Mux_v I__12222 (
            .O(N__48100),
            .I(N__48017));
    Span4Mux_h I__12221 (
            .O(N__48097),
            .I(N__48014));
    InMux I__12220 (
            .O(N__48096),
            .I(N__48007));
    InMux I__12219 (
            .O(N__48095),
            .I(N__48007));
    InMux I__12218 (
            .O(N__48094),
            .I(N__48007));
    InMux I__12217 (
            .O(N__48093),
            .I(N__48002));
    InMux I__12216 (
            .O(N__48092),
            .I(N__48002));
    LocalMux I__12215 (
            .O(N__48089),
            .I(N__47997));
    Span4Mux_v I__12214 (
            .O(N__48078),
            .I(N__47997));
    InMux I__12213 (
            .O(N__48077),
            .I(N__47990));
    InMux I__12212 (
            .O(N__48076),
            .I(N__47990));
    InMux I__12211 (
            .O(N__48075),
            .I(N__47990));
    InMux I__12210 (
            .O(N__48074),
            .I(N__47987));
    Span4Mux_v I__12209 (
            .O(N__48065),
            .I(N__47984));
    Span4Mux_v I__12208 (
            .O(N__48060),
            .I(N__47979));
    Span4Mux_v I__12207 (
            .O(N__48055),
            .I(N__47979));
    CascadeMux I__12206 (
            .O(N__48054),
            .I(N__47976));
    Span4Mux_v I__12205 (
            .O(N__48049),
            .I(N__47971));
    Span4Mux_v I__12204 (
            .O(N__48034),
            .I(N__47971));
    Span4Mux_h I__12203 (
            .O(N__48031),
            .I(N__47968));
    InMux I__12202 (
            .O(N__48030),
            .I(N__47963));
    InMux I__12201 (
            .O(N__48029),
            .I(N__47963));
    LocalMux I__12200 (
            .O(N__48026),
            .I(N__47958));
    Span4Mux_s1_h I__12199 (
            .O(N__48023),
            .I(N__47958));
    LocalMux I__12198 (
            .O(N__48020),
            .I(N__47953));
    Span4Mux_v I__12197 (
            .O(N__48017),
            .I(N__47953));
    Sp12to4 I__12196 (
            .O(N__48014),
            .I(N__47950));
    LocalMux I__12195 (
            .O(N__48007),
            .I(N__47941));
    LocalMux I__12194 (
            .O(N__48002),
            .I(N__47941));
    Sp12to4 I__12193 (
            .O(N__47997),
            .I(N__47941));
    LocalMux I__12192 (
            .O(N__47990),
            .I(N__47941));
    LocalMux I__12191 (
            .O(N__47987),
            .I(N__47934));
    Span4Mux_v I__12190 (
            .O(N__47984),
            .I(N__47934));
    Span4Mux_v I__12189 (
            .O(N__47979),
            .I(N__47934));
    InMux I__12188 (
            .O(N__47976),
            .I(N__47931));
    Span4Mux_h I__12187 (
            .O(N__47971),
            .I(N__47928));
    Span4Mux_v I__12186 (
            .O(N__47968),
            .I(N__47925));
    LocalMux I__12185 (
            .O(N__47963),
            .I(N__47918));
    Span4Mux_v I__12184 (
            .O(N__47958),
            .I(N__47918));
    Span4Mux_h I__12183 (
            .O(N__47953),
            .I(N__47918));
    Span12Mux_v I__12182 (
            .O(N__47950),
            .I(N__47913));
    Span12Mux_h I__12181 (
            .O(N__47941),
            .I(N__47913));
    Span4Mux_h I__12180 (
            .O(N__47934),
            .I(N__47908));
    LocalMux I__12179 (
            .O(N__47931),
            .I(N__47908));
    Span4Mux_h I__12178 (
            .O(N__47928),
            .I(N__47905));
    Odrv4 I__12177 (
            .O(N__47925),
            .I(aluOperation_0));
    Odrv4 I__12176 (
            .O(N__47918),
            .I(aluOperation_0));
    Odrv12 I__12175 (
            .O(N__47913),
            .I(aluOperation_0));
    Odrv4 I__12174 (
            .O(N__47908),
            .I(aluOperation_0));
    Odrv4 I__12173 (
            .O(N__47905),
            .I(aluOperation_0));
    InMux I__12172 (
            .O(N__47894),
            .I(N__47889));
    InMux I__12171 (
            .O(N__47893),
            .I(N__47883));
    InMux I__12170 (
            .O(N__47892),
            .I(N__47880));
    LocalMux I__12169 (
            .O(N__47889),
            .I(N__47877));
    InMux I__12168 (
            .O(N__47888),
            .I(N__47874));
    InMux I__12167 (
            .O(N__47887),
            .I(N__47871));
    InMux I__12166 (
            .O(N__47886),
            .I(N__47868));
    LocalMux I__12165 (
            .O(N__47883),
            .I(N__47865));
    LocalMux I__12164 (
            .O(N__47880),
            .I(N__47861));
    Span4Mux_h I__12163 (
            .O(N__47877),
            .I(N__47858));
    LocalMux I__12162 (
            .O(N__47874),
            .I(N__47853));
    LocalMux I__12161 (
            .O(N__47871),
            .I(N__47853));
    LocalMux I__12160 (
            .O(N__47868),
            .I(N__47850));
    Span4Mux_v I__12159 (
            .O(N__47865),
            .I(N__47847));
    InMux I__12158 (
            .O(N__47864),
            .I(N__47844));
    Span4Mux_v I__12157 (
            .O(N__47861),
            .I(N__47841));
    Span4Mux_h I__12156 (
            .O(N__47858),
            .I(N__47836));
    Span4Mux_s2_v I__12155 (
            .O(N__47853),
            .I(N__47836));
    Span4Mux_v I__12154 (
            .O(N__47850),
            .I(N__47833));
    Span4Mux_h I__12153 (
            .O(N__47847),
            .I(N__47828));
    LocalMux I__12152 (
            .O(N__47844),
            .I(N__47828));
    Span4Mux_v I__12151 (
            .O(N__47841),
            .I(N__47818));
    Span4Mux_v I__12150 (
            .O(N__47836),
            .I(N__47818));
    Span4Mux_v I__12149 (
            .O(N__47833),
            .I(N__47818));
    Span4Mux_h I__12148 (
            .O(N__47828),
            .I(N__47818));
    InMux I__12147 (
            .O(N__47827),
            .I(N__47815));
    Odrv4 I__12146 (
            .O(N__47818),
            .I(\ALU.un9_addsub_cry_7_c_RNIQIKVOZ0 ));
    LocalMux I__12145 (
            .O(N__47815),
            .I(\ALU.un9_addsub_cry_7_c_RNIQIKVOZ0 ));
    InMux I__12144 (
            .O(N__47810),
            .I(N__47805));
    InMux I__12143 (
            .O(N__47809),
            .I(N__47802));
    InMux I__12142 (
            .O(N__47808),
            .I(N__47799));
    LocalMux I__12141 (
            .O(N__47805),
            .I(N__47795));
    LocalMux I__12140 (
            .O(N__47802),
            .I(N__47791));
    LocalMux I__12139 (
            .O(N__47799),
            .I(N__47788));
    InMux I__12138 (
            .O(N__47798),
            .I(N__47785));
    Span4Mux_v I__12137 (
            .O(N__47795),
            .I(N__47782));
    InMux I__12136 (
            .O(N__47794),
            .I(N__47779));
    Span4Mux_h I__12135 (
            .O(N__47791),
            .I(N__47774));
    Span4Mux_h I__12134 (
            .O(N__47788),
            .I(N__47771));
    LocalMux I__12133 (
            .O(N__47785),
            .I(N__47768));
    Span4Mux_h I__12132 (
            .O(N__47782),
            .I(N__47763));
    LocalMux I__12131 (
            .O(N__47779),
            .I(N__47763));
    InMux I__12130 (
            .O(N__47778),
            .I(N__47760));
    InMux I__12129 (
            .O(N__47777),
            .I(N__47757));
    Span4Mux_h I__12128 (
            .O(N__47774),
            .I(N__47753));
    Span4Mux_h I__12127 (
            .O(N__47771),
            .I(N__47750));
    Span4Mux_s3_v I__12126 (
            .O(N__47768),
            .I(N__47747));
    Span4Mux_v I__12125 (
            .O(N__47763),
            .I(N__47744));
    LocalMux I__12124 (
            .O(N__47760),
            .I(N__47741));
    LocalMux I__12123 (
            .O(N__47757),
            .I(N__47738));
    InMux I__12122 (
            .O(N__47756),
            .I(N__47735));
    Odrv4 I__12121 (
            .O(N__47753),
            .I(\ALU.d_RNI7GCMD22Z0Z_8 ));
    Odrv4 I__12120 (
            .O(N__47750),
            .I(\ALU.d_RNI7GCMD22Z0Z_8 ));
    Odrv4 I__12119 (
            .O(N__47747),
            .I(\ALU.d_RNI7GCMD22Z0Z_8 ));
    Odrv4 I__12118 (
            .O(N__47744),
            .I(\ALU.d_RNI7GCMD22Z0Z_8 ));
    Odrv12 I__12117 (
            .O(N__47741),
            .I(\ALU.d_RNI7GCMD22Z0Z_8 ));
    Odrv12 I__12116 (
            .O(N__47738),
            .I(\ALU.d_RNI7GCMD22Z0Z_8 ));
    LocalMux I__12115 (
            .O(N__47735),
            .I(\ALU.d_RNI7GCMD22Z0Z_8 ));
    InMux I__12114 (
            .O(N__47720),
            .I(N__47716));
    InMux I__12113 (
            .O(N__47719),
            .I(N__47713));
    LocalMux I__12112 (
            .O(N__47716),
            .I(N__47710));
    LocalMux I__12111 (
            .O(N__47713),
            .I(N__47707));
    Span4Mux_v I__12110 (
            .O(N__47710),
            .I(N__47702));
    Span4Mux_v I__12109 (
            .O(N__47707),
            .I(N__47702));
    Span4Mux_h I__12108 (
            .O(N__47702),
            .I(N__47699));
    Span4Mux_h I__12107 (
            .O(N__47699),
            .I(N__47696));
    Odrv4 I__12106 (
            .O(N__47696),
            .I(\ALU.bZ0Z_8 ));
    ClkMux I__12105 (
            .O(N__47693),
            .I(N__47408));
    ClkMux I__12104 (
            .O(N__47692),
            .I(N__47408));
    ClkMux I__12103 (
            .O(N__47691),
            .I(N__47408));
    ClkMux I__12102 (
            .O(N__47690),
            .I(N__47408));
    ClkMux I__12101 (
            .O(N__47689),
            .I(N__47408));
    ClkMux I__12100 (
            .O(N__47688),
            .I(N__47408));
    ClkMux I__12099 (
            .O(N__47687),
            .I(N__47408));
    ClkMux I__12098 (
            .O(N__47686),
            .I(N__47408));
    ClkMux I__12097 (
            .O(N__47685),
            .I(N__47408));
    ClkMux I__12096 (
            .O(N__47684),
            .I(N__47408));
    ClkMux I__12095 (
            .O(N__47683),
            .I(N__47408));
    ClkMux I__12094 (
            .O(N__47682),
            .I(N__47408));
    ClkMux I__12093 (
            .O(N__47681),
            .I(N__47408));
    ClkMux I__12092 (
            .O(N__47680),
            .I(N__47408));
    ClkMux I__12091 (
            .O(N__47679),
            .I(N__47408));
    ClkMux I__12090 (
            .O(N__47678),
            .I(N__47408));
    ClkMux I__12089 (
            .O(N__47677),
            .I(N__47408));
    ClkMux I__12088 (
            .O(N__47676),
            .I(N__47408));
    ClkMux I__12087 (
            .O(N__47675),
            .I(N__47408));
    ClkMux I__12086 (
            .O(N__47674),
            .I(N__47408));
    ClkMux I__12085 (
            .O(N__47673),
            .I(N__47408));
    ClkMux I__12084 (
            .O(N__47672),
            .I(N__47408));
    ClkMux I__12083 (
            .O(N__47671),
            .I(N__47408));
    ClkMux I__12082 (
            .O(N__47670),
            .I(N__47408));
    ClkMux I__12081 (
            .O(N__47669),
            .I(N__47408));
    ClkMux I__12080 (
            .O(N__47668),
            .I(N__47408));
    ClkMux I__12079 (
            .O(N__47667),
            .I(N__47408));
    ClkMux I__12078 (
            .O(N__47666),
            .I(N__47408));
    ClkMux I__12077 (
            .O(N__47665),
            .I(N__47408));
    ClkMux I__12076 (
            .O(N__47664),
            .I(N__47408));
    ClkMux I__12075 (
            .O(N__47663),
            .I(N__47408));
    ClkMux I__12074 (
            .O(N__47662),
            .I(N__47408));
    ClkMux I__12073 (
            .O(N__47661),
            .I(N__47408));
    ClkMux I__12072 (
            .O(N__47660),
            .I(N__47408));
    ClkMux I__12071 (
            .O(N__47659),
            .I(N__47408));
    ClkMux I__12070 (
            .O(N__47658),
            .I(N__47408));
    ClkMux I__12069 (
            .O(N__47657),
            .I(N__47408));
    ClkMux I__12068 (
            .O(N__47656),
            .I(N__47408));
    ClkMux I__12067 (
            .O(N__47655),
            .I(N__47408));
    ClkMux I__12066 (
            .O(N__47654),
            .I(N__47408));
    ClkMux I__12065 (
            .O(N__47653),
            .I(N__47408));
    ClkMux I__12064 (
            .O(N__47652),
            .I(N__47408));
    ClkMux I__12063 (
            .O(N__47651),
            .I(N__47408));
    ClkMux I__12062 (
            .O(N__47650),
            .I(N__47408));
    ClkMux I__12061 (
            .O(N__47649),
            .I(N__47408));
    ClkMux I__12060 (
            .O(N__47648),
            .I(N__47408));
    ClkMux I__12059 (
            .O(N__47647),
            .I(N__47408));
    ClkMux I__12058 (
            .O(N__47646),
            .I(N__47408));
    ClkMux I__12057 (
            .O(N__47645),
            .I(N__47408));
    ClkMux I__12056 (
            .O(N__47644),
            .I(N__47408));
    ClkMux I__12055 (
            .O(N__47643),
            .I(N__47408));
    ClkMux I__12054 (
            .O(N__47642),
            .I(N__47408));
    ClkMux I__12053 (
            .O(N__47641),
            .I(N__47408));
    ClkMux I__12052 (
            .O(N__47640),
            .I(N__47408));
    ClkMux I__12051 (
            .O(N__47639),
            .I(N__47408));
    ClkMux I__12050 (
            .O(N__47638),
            .I(N__47408));
    ClkMux I__12049 (
            .O(N__47637),
            .I(N__47408));
    ClkMux I__12048 (
            .O(N__47636),
            .I(N__47408));
    ClkMux I__12047 (
            .O(N__47635),
            .I(N__47408));
    ClkMux I__12046 (
            .O(N__47634),
            .I(N__47408));
    ClkMux I__12045 (
            .O(N__47633),
            .I(N__47408));
    ClkMux I__12044 (
            .O(N__47632),
            .I(N__47408));
    ClkMux I__12043 (
            .O(N__47631),
            .I(N__47408));
    ClkMux I__12042 (
            .O(N__47630),
            .I(N__47408));
    ClkMux I__12041 (
            .O(N__47629),
            .I(N__47408));
    ClkMux I__12040 (
            .O(N__47628),
            .I(N__47408));
    ClkMux I__12039 (
            .O(N__47627),
            .I(N__47408));
    ClkMux I__12038 (
            .O(N__47626),
            .I(N__47408));
    ClkMux I__12037 (
            .O(N__47625),
            .I(N__47408));
    ClkMux I__12036 (
            .O(N__47624),
            .I(N__47408));
    ClkMux I__12035 (
            .O(N__47623),
            .I(N__47408));
    ClkMux I__12034 (
            .O(N__47622),
            .I(N__47408));
    ClkMux I__12033 (
            .O(N__47621),
            .I(N__47408));
    ClkMux I__12032 (
            .O(N__47620),
            .I(N__47408));
    ClkMux I__12031 (
            .O(N__47619),
            .I(N__47408));
    ClkMux I__12030 (
            .O(N__47618),
            .I(N__47408));
    ClkMux I__12029 (
            .O(N__47617),
            .I(N__47408));
    ClkMux I__12028 (
            .O(N__47616),
            .I(N__47408));
    ClkMux I__12027 (
            .O(N__47615),
            .I(N__47408));
    ClkMux I__12026 (
            .O(N__47614),
            .I(N__47408));
    ClkMux I__12025 (
            .O(N__47613),
            .I(N__47408));
    ClkMux I__12024 (
            .O(N__47612),
            .I(N__47408));
    ClkMux I__12023 (
            .O(N__47611),
            .I(N__47408));
    ClkMux I__12022 (
            .O(N__47610),
            .I(N__47408));
    ClkMux I__12021 (
            .O(N__47609),
            .I(N__47408));
    ClkMux I__12020 (
            .O(N__47608),
            .I(N__47408));
    ClkMux I__12019 (
            .O(N__47607),
            .I(N__47408));
    ClkMux I__12018 (
            .O(N__47606),
            .I(N__47408));
    ClkMux I__12017 (
            .O(N__47605),
            .I(N__47408));
    ClkMux I__12016 (
            .O(N__47604),
            .I(N__47408));
    ClkMux I__12015 (
            .O(N__47603),
            .I(N__47408));
    ClkMux I__12014 (
            .O(N__47602),
            .I(N__47408));
    ClkMux I__12013 (
            .O(N__47601),
            .I(N__47408));
    ClkMux I__12012 (
            .O(N__47600),
            .I(N__47408));
    ClkMux I__12011 (
            .O(N__47599),
            .I(N__47408));
    GlobalMux I__12010 (
            .O(N__47408),
            .I(N__47405));
    gio2CtrlBuf I__12009 (
            .O(N__47405),
            .I(CLK_0_c_g));
    CEMux I__12008 (
            .O(N__47402),
            .I(N__47398));
    CEMux I__12007 (
            .O(N__47401),
            .I(N__47394));
    LocalMux I__12006 (
            .O(N__47398),
            .I(N__47390));
    CEMux I__12005 (
            .O(N__47397),
            .I(N__47387));
    LocalMux I__12004 (
            .O(N__47394),
            .I(N__47384));
    CEMux I__12003 (
            .O(N__47393),
            .I(N__47381));
    Span4Mux_h I__12002 (
            .O(N__47390),
            .I(N__47378));
    LocalMux I__12001 (
            .O(N__47387),
            .I(N__47375));
    Span4Mux_v I__12000 (
            .O(N__47384),
            .I(N__47372));
    LocalMux I__11999 (
            .O(N__47381),
            .I(N__47369));
    Span4Mux_h I__11998 (
            .O(N__47378),
            .I(N__47366));
    Span4Mux_h I__11997 (
            .O(N__47375),
            .I(N__47363));
    Span4Mux_v I__11996 (
            .O(N__47372),
            .I(N__47360));
    Span4Mux_h I__11995 (
            .O(N__47369),
            .I(N__47357));
    Span4Mux_v I__11994 (
            .O(N__47366),
            .I(N__47354));
    Span4Mux_v I__11993 (
            .O(N__47363),
            .I(N__47351));
    Span4Mux_v I__11992 (
            .O(N__47360),
            .I(N__47348));
    Sp12to4 I__11991 (
            .O(N__47357),
            .I(N__47343));
    Sp12to4 I__11990 (
            .O(N__47354),
            .I(N__47343));
    Span4Mux_v I__11989 (
            .O(N__47351),
            .I(N__47340));
    Sp12to4 I__11988 (
            .O(N__47348),
            .I(N__47337));
    Span12Mux_h I__11987 (
            .O(N__47343),
            .I(N__47334));
    Span4Mux_h I__11986 (
            .O(N__47340),
            .I(N__47331));
    Odrv12 I__11985 (
            .O(N__47337),
            .I(\ALU.b_cnvZ0Z_0 ));
    Odrv12 I__11984 (
            .O(N__47334),
            .I(\ALU.b_cnvZ0Z_0 ));
    Odrv4 I__11983 (
            .O(N__47331),
            .I(\ALU.b_cnvZ0Z_0 ));
    InMux I__11982 (
            .O(N__47324),
            .I(N__47315));
    InMux I__11981 (
            .O(N__47323),
            .I(N__47315));
    InMux I__11980 (
            .O(N__47322),
            .I(N__47311));
    CascadeMux I__11979 (
            .O(N__47321),
            .I(N__47305));
    InMux I__11978 (
            .O(N__47320),
            .I(N__47300));
    LocalMux I__11977 (
            .O(N__47315),
            .I(N__47297));
    InMux I__11976 (
            .O(N__47314),
            .I(N__47294));
    LocalMux I__11975 (
            .O(N__47311),
            .I(N__47289));
    InMux I__11974 (
            .O(N__47310),
            .I(N__47286));
    InMux I__11973 (
            .O(N__47309),
            .I(N__47283));
    InMux I__11972 (
            .O(N__47308),
            .I(N__47280));
    InMux I__11971 (
            .O(N__47305),
            .I(N__47274));
    InMux I__11970 (
            .O(N__47304),
            .I(N__47269));
    InMux I__11969 (
            .O(N__47303),
            .I(N__47269));
    LocalMux I__11968 (
            .O(N__47300),
            .I(N__47264));
    Span4Mux_v I__11967 (
            .O(N__47297),
            .I(N__47264));
    LocalMux I__11966 (
            .O(N__47294),
            .I(N__47261));
    InMux I__11965 (
            .O(N__47293),
            .I(N__47256));
    InMux I__11964 (
            .O(N__47292),
            .I(N__47253));
    Span4Mux_v I__11963 (
            .O(N__47289),
            .I(N__47246));
    LocalMux I__11962 (
            .O(N__47286),
            .I(N__47246));
    LocalMux I__11961 (
            .O(N__47283),
            .I(N__47246));
    LocalMux I__11960 (
            .O(N__47280),
            .I(N__47243));
    InMux I__11959 (
            .O(N__47279),
            .I(N__47238));
    InMux I__11958 (
            .O(N__47278),
            .I(N__47238));
    InMux I__11957 (
            .O(N__47277),
            .I(N__47235));
    LocalMux I__11956 (
            .O(N__47274),
            .I(N__47224));
    LocalMux I__11955 (
            .O(N__47269),
            .I(N__47224));
    Span4Mux_v I__11954 (
            .O(N__47264),
            .I(N__47221));
    Span4Mux_v I__11953 (
            .O(N__47261),
            .I(N__47217));
    InMux I__11952 (
            .O(N__47260),
            .I(N__47212));
    InMux I__11951 (
            .O(N__47259),
            .I(N__47212));
    LocalMux I__11950 (
            .O(N__47256),
            .I(N__47205));
    LocalMux I__11949 (
            .O(N__47253),
            .I(N__47205));
    Span4Mux_v I__11948 (
            .O(N__47246),
            .I(N__47202));
    Span4Mux_v I__11947 (
            .O(N__47243),
            .I(N__47199));
    LocalMux I__11946 (
            .O(N__47238),
            .I(N__47194));
    LocalMux I__11945 (
            .O(N__47235),
            .I(N__47194));
    InMux I__11944 (
            .O(N__47234),
            .I(N__47185));
    InMux I__11943 (
            .O(N__47233),
            .I(N__47185));
    InMux I__11942 (
            .O(N__47232),
            .I(N__47185));
    InMux I__11941 (
            .O(N__47231),
            .I(N__47185));
    InMux I__11940 (
            .O(N__47230),
            .I(N__47180));
    InMux I__11939 (
            .O(N__47229),
            .I(N__47180));
    Span4Mux_v I__11938 (
            .O(N__47224),
            .I(N__47173));
    Span4Mux_h I__11937 (
            .O(N__47221),
            .I(N__47173));
    InMux I__11936 (
            .O(N__47220),
            .I(N__47170));
    Span4Mux_h I__11935 (
            .O(N__47217),
            .I(N__47165));
    LocalMux I__11934 (
            .O(N__47212),
            .I(N__47165));
    InMux I__11933 (
            .O(N__47211),
            .I(N__47160));
    InMux I__11932 (
            .O(N__47210),
            .I(N__47160));
    Span4Mux_v I__11931 (
            .O(N__47205),
            .I(N__47157));
    Span4Mux_v I__11930 (
            .O(N__47202),
            .I(N__47154));
    Span4Mux_v I__11929 (
            .O(N__47199),
            .I(N__47151));
    Span4Mux_v I__11928 (
            .O(N__47194),
            .I(N__47146));
    LocalMux I__11927 (
            .O(N__47185),
            .I(N__47146));
    LocalMux I__11926 (
            .O(N__47180),
            .I(N__47143));
    InMux I__11925 (
            .O(N__47179),
            .I(N__47140));
    InMux I__11924 (
            .O(N__47178),
            .I(N__47137));
    Span4Mux_v I__11923 (
            .O(N__47173),
            .I(N__47134));
    LocalMux I__11922 (
            .O(N__47170),
            .I(N__47125));
    Span4Mux_v I__11921 (
            .O(N__47165),
            .I(N__47125));
    LocalMux I__11920 (
            .O(N__47160),
            .I(N__47125));
    Span4Mux_h I__11919 (
            .O(N__47157),
            .I(N__47125));
    Span4Mux_h I__11918 (
            .O(N__47154),
            .I(N__47116));
    Span4Mux_h I__11917 (
            .O(N__47151),
            .I(N__47116));
    Span4Mux_v I__11916 (
            .O(N__47146),
            .I(N__47116));
    Span4Mux_s2_v I__11915 (
            .O(N__47143),
            .I(N__47116));
    LocalMux I__11914 (
            .O(N__47140),
            .I(\ALU.a_15_sm0 ));
    LocalMux I__11913 (
            .O(N__47137),
            .I(\ALU.a_15_sm0 ));
    Odrv4 I__11912 (
            .O(N__47134),
            .I(\ALU.a_15_sm0 ));
    Odrv4 I__11911 (
            .O(N__47125),
            .I(\ALU.a_15_sm0 ));
    Odrv4 I__11910 (
            .O(N__47116),
            .I(\ALU.a_15_sm0 ));
    InMux I__11909 (
            .O(N__47105),
            .I(N__47102));
    LocalMux I__11908 (
            .O(N__47102),
            .I(N__47093));
    InMux I__11907 (
            .O(N__47101),
            .I(N__47090));
    InMux I__11906 (
            .O(N__47100),
            .I(N__47084));
    InMux I__11905 (
            .O(N__47099),
            .I(N__47077));
    InMux I__11904 (
            .O(N__47098),
            .I(N__47077));
    InMux I__11903 (
            .O(N__47097),
            .I(N__47077));
    InMux I__11902 (
            .O(N__47096),
            .I(N__47074));
    Span4Mux_v I__11901 (
            .O(N__47093),
            .I(N__47071));
    LocalMux I__11900 (
            .O(N__47090),
            .I(N__47068));
    InMux I__11899 (
            .O(N__47089),
            .I(N__47064));
    InMux I__11898 (
            .O(N__47088),
            .I(N__47061));
    InMux I__11897 (
            .O(N__47087),
            .I(N__47058));
    LocalMux I__11896 (
            .O(N__47084),
            .I(N__47055));
    LocalMux I__11895 (
            .O(N__47077),
            .I(N__47052));
    LocalMux I__11894 (
            .O(N__47074),
            .I(N__47046));
    Span4Mux_h I__11893 (
            .O(N__47071),
            .I(N__47043));
    Span4Mux_v I__11892 (
            .O(N__47068),
            .I(N__47040));
    InMux I__11891 (
            .O(N__47067),
            .I(N__47037));
    LocalMux I__11890 (
            .O(N__47064),
            .I(N__47032));
    LocalMux I__11889 (
            .O(N__47061),
            .I(N__47032));
    LocalMux I__11888 (
            .O(N__47058),
            .I(N__47025));
    Span4Mux_h I__11887 (
            .O(N__47055),
            .I(N__47025));
    Span4Mux_v I__11886 (
            .O(N__47052),
            .I(N__47025));
    InMux I__11885 (
            .O(N__47051),
            .I(N__47022));
    InMux I__11884 (
            .O(N__47050),
            .I(N__47017));
    InMux I__11883 (
            .O(N__47049),
            .I(N__47017));
    Span4Mux_v I__11882 (
            .O(N__47046),
            .I(N__47014));
    Span4Mux_h I__11881 (
            .O(N__47043),
            .I(N__47005));
    Span4Mux_v I__11880 (
            .O(N__47040),
            .I(N__47005));
    LocalMux I__11879 (
            .O(N__47037),
            .I(N__47005));
    Span4Mux_v I__11878 (
            .O(N__47032),
            .I(N__47005));
    Span4Mux_v I__11877 (
            .O(N__47025),
            .I(N__47002));
    LocalMux I__11876 (
            .O(N__47022),
            .I(\ALU.N_213_0 ));
    LocalMux I__11875 (
            .O(N__47017),
            .I(\ALU.N_213_0 ));
    Odrv4 I__11874 (
            .O(N__47014),
            .I(\ALU.N_213_0 ));
    Odrv4 I__11873 (
            .O(N__47005),
            .I(\ALU.N_213_0 ));
    Odrv4 I__11872 (
            .O(N__47002),
            .I(\ALU.N_213_0 ));
    CascadeMux I__11871 (
            .O(N__46991),
            .I(N__46988));
    InMux I__11870 (
            .O(N__46988),
            .I(N__46985));
    LocalMux I__11869 (
            .O(N__46985),
            .I(N__46982));
    Span4Mux_h I__11868 (
            .O(N__46982),
            .I(N__46979));
    Odrv4 I__11867 (
            .O(N__46979),
            .I(\ALU.a_15_m2_ns_1Z0Z_7 ));
    InMux I__11866 (
            .O(N__46976),
            .I(N__46970));
    InMux I__11865 (
            .O(N__46975),
            .I(N__46967));
    InMux I__11864 (
            .O(N__46974),
            .I(N__46957));
    CascadeMux I__11863 (
            .O(N__46973),
            .I(N__46953));
    LocalMux I__11862 (
            .O(N__46970),
            .I(N__46950));
    LocalMux I__11861 (
            .O(N__46967),
            .I(N__46947));
    InMux I__11860 (
            .O(N__46966),
            .I(N__46937));
    InMux I__11859 (
            .O(N__46965),
            .I(N__46937));
    InMux I__11858 (
            .O(N__46964),
            .I(N__46934));
    InMux I__11857 (
            .O(N__46963),
            .I(N__46931));
    InMux I__11856 (
            .O(N__46962),
            .I(N__46928));
    InMux I__11855 (
            .O(N__46961),
            .I(N__46925));
    InMux I__11854 (
            .O(N__46960),
            .I(N__46922));
    LocalMux I__11853 (
            .O(N__46957),
            .I(N__46919));
    InMux I__11852 (
            .O(N__46956),
            .I(N__46913));
    InMux I__11851 (
            .O(N__46953),
            .I(N__46913));
    Span4Mux_h I__11850 (
            .O(N__46950),
            .I(N__46908));
    Span4Mux_h I__11849 (
            .O(N__46947),
            .I(N__46904));
    InMux I__11848 (
            .O(N__46946),
            .I(N__46899));
    InMux I__11847 (
            .O(N__46945),
            .I(N__46899));
    InMux I__11846 (
            .O(N__46944),
            .I(N__46896));
    InMux I__11845 (
            .O(N__46943),
            .I(N__46893));
    InMux I__11844 (
            .O(N__46942),
            .I(N__46890));
    LocalMux I__11843 (
            .O(N__46937),
            .I(N__46887));
    LocalMux I__11842 (
            .O(N__46934),
            .I(N__46884));
    LocalMux I__11841 (
            .O(N__46931),
            .I(N__46877));
    LocalMux I__11840 (
            .O(N__46928),
            .I(N__46877));
    LocalMux I__11839 (
            .O(N__46925),
            .I(N__46877));
    LocalMux I__11838 (
            .O(N__46922),
            .I(N__46873));
    Span4Mux_h I__11837 (
            .O(N__46919),
            .I(N__46870));
    InMux I__11836 (
            .O(N__46918),
            .I(N__46867));
    LocalMux I__11835 (
            .O(N__46913),
            .I(N__46864));
    InMux I__11834 (
            .O(N__46912),
            .I(N__46861));
    InMux I__11833 (
            .O(N__46911),
            .I(N__46858));
    Span4Mux_h I__11832 (
            .O(N__46908),
            .I(N__46855));
    InMux I__11831 (
            .O(N__46907),
            .I(N__46852));
    Span4Mux_h I__11830 (
            .O(N__46904),
            .I(N__46847));
    LocalMux I__11829 (
            .O(N__46899),
            .I(N__46847));
    LocalMux I__11828 (
            .O(N__46896),
            .I(N__46840));
    LocalMux I__11827 (
            .O(N__46893),
            .I(N__46840));
    LocalMux I__11826 (
            .O(N__46890),
            .I(N__46840));
    Span4Mux_h I__11825 (
            .O(N__46887),
            .I(N__46834));
    Span4Mux_h I__11824 (
            .O(N__46884),
            .I(N__46831));
    Span4Mux_v I__11823 (
            .O(N__46877),
            .I(N__46828));
    InMux I__11822 (
            .O(N__46876),
            .I(N__46825));
    Span4Mux_v I__11821 (
            .O(N__46873),
            .I(N__46820));
    Span4Mux_v I__11820 (
            .O(N__46870),
            .I(N__46820));
    LocalMux I__11819 (
            .O(N__46867),
            .I(N__46817));
    Span4Mux_v I__11818 (
            .O(N__46864),
            .I(N__46814));
    LocalMux I__11817 (
            .O(N__46861),
            .I(N__46808));
    LocalMux I__11816 (
            .O(N__46858),
            .I(N__46808));
    Span4Mux_h I__11815 (
            .O(N__46855),
            .I(N__46799));
    LocalMux I__11814 (
            .O(N__46852),
            .I(N__46799));
    Span4Mux_v I__11813 (
            .O(N__46847),
            .I(N__46799));
    Span4Mux_h I__11812 (
            .O(N__46840),
            .I(N__46799));
    InMux I__11811 (
            .O(N__46839),
            .I(N__46794));
    InMux I__11810 (
            .O(N__46838),
            .I(N__46794));
    InMux I__11809 (
            .O(N__46837),
            .I(N__46791));
    Span4Mux_v I__11808 (
            .O(N__46834),
            .I(N__46788));
    Span4Mux_h I__11807 (
            .O(N__46831),
            .I(N__46783));
    Span4Mux_s2_h I__11806 (
            .O(N__46828),
            .I(N__46783));
    LocalMux I__11805 (
            .O(N__46825),
            .I(N__46780));
    Span4Mux_v I__11804 (
            .O(N__46820),
            .I(N__46773));
    Span4Mux_h I__11803 (
            .O(N__46817),
            .I(N__46773));
    Span4Mux_h I__11802 (
            .O(N__46814),
            .I(N__46773));
    InMux I__11801 (
            .O(N__46813),
            .I(N__46770));
    Span4Mux_h I__11800 (
            .O(N__46808),
            .I(N__46763));
    Span4Mux_v I__11799 (
            .O(N__46799),
            .I(N__46763));
    LocalMux I__11798 (
            .O(N__46794),
            .I(N__46763));
    LocalMux I__11797 (
            .O(N__46791),
            .I(\ALU.aluOut_7 ));
    Odrv4 I__11796 (
            .O(N__46788),
            .I(\ALU.aluOut_7 ));
    Odrv4 I__11795 (
            .O(N__46783),
            .I(\ALU.aluOut_7 ));
    Odrv12 I__11794 (
            .O(N__46780),
            .I(\ALU.aluOut_7 ));
    Odrv4 I__11793 (
            .O(N__46773),
            .I(\ALU.aluOut_7 ));
    LocalMux I__11792 (
            .O(N__46770),
            .I(\ALU.aluOut_7 ));
    Odrv4 I__11791 (
            .O(N__46763),
            .I(\ALU.aluOut_7 ));
    CascadeMux I__11790 (
            .O(N__46748),
            .I(N__46745));
    InMux I__11789 (
            .O(N__46745),
            .I(N__46742));
    LocalMux I__11788 (
            .O(N__46742),
            .I(N__46739));
    Odrv4 I__11787 (
            .O(N__46739),
            .I(\ALU.a_15_m2_7 ));
    InMux I__11786 (
            .O(N__46736),
            .I(N__46730));
    InMux I__11785 (
            .O(N__46735),
            .I(N__46724));
    InMux I__11784 (
            .O(N__46734),
            .I(N__46721));
    InMux I__11783 (
            .O(N__46733),
            .I(N__46717));
    LocalMux I__11782 (
            .O(N__46730),
            .I(N__46712));
    InMux I__11781 (
            .O(N__46729),
            .I(N__46709));
    InMux I__11780 (
            .O(N__46728),
            .I(N__46706));
    InMux I__11779 (
            .O(N__46727),
            .I(N__46703));
    LocalMux I__11778 (
            .O(N__46724),
            .I(N__46700));
    LocalMux I__11777 (
            .O(N__46721),
            .I(N__46697));
    InMux I__11776 (
            .O(N__46720),
            .I(N__46694));
    LocalMux I__11775 (
            .O(N__46717),
            .I(N__46690));
    InMux I__11774 (
            .O(N__46716),
            .I(N__46687));
    InMux I__11773 (
            .O(N__46715),
            .I(N__46683));
    Span4Mux_s3_h I__11772 (
            .O(N__46712),
            .I(N__46676));
    LocalMux I__11771 (
            .O(N__46709),
            .I(N__46676));
    LocalMux I__11770 (
            .O(N__46706),
            .I(N__46673));
    LocalMux I__11769 (
            .O(N__46703),
            .I(N__46666));
    Span4Mux_h I__11768 (
            .O(N__46700),
            .I(N__46659));
    Span4Mux_s2_v I__11767 (
            .O(N__46697),
            .I(N__46659));
    LocalMux I__11766 (
            .O(N__46694),
            .I(N__46659));
    InMux I__11765 (
            .O(N__46693),
            .I(N__46654));
    Span4Mux_v I__11764 (
            .O(N__46690),
            .I(N__46649));
    LocalMux I__11763 (
            .O(N__46687),
            .I(N__46649));
    InMux I__11762 (
            .O(N__46686),
            .I(N__46645));
    LocalMux I__11761 (
            .O(N__46683),
            .I(N__46642));
    CascadeMux I__11760 (
            .O(N__46682),
            .I(N__46639));
    InMux I__11759 (
            .O(N__46681),
            .I(N__46635));
    Span4Mux_h I__11758 (
            .O(N__46676),
            .I(N__46630));
    Span4Mux_s3_h I__11757 (
            .O(N__46673),
            .I(N__46630));
    InMux I__11756 (
            .O(N__46672),
            .I(N__46627));
    InMux I__11755 (
            .O(N__46671),
            .I(N__46623));
    InMux I__11754 (
            .O(N__46670),
            .I(N__46617));
    InMux I__11753 (
            .O(N__46669),
            .I(N__46617));
    Span4Mux_v I__11752 (
            .O(N__46666),
            .I(N__46612));
    Span4Mux_v I__11751 (
            .O(N__46659),
            .I(N__46609));
    InMux I__11750 (
            .O(N__46658),
            .I(N__46606));
    InMux I__11749 (
            .O(N__46657),
            .I(N__46603));
    LocalMux I__11748 (
            .O(N__46654),
            .I(N__46600));
    Span4Mux_h I__11747 (
            .O(N__46649),
            .I(N__46597));
    InMux I__11746 (
            .O(N__46648),
            .I(N__46594));
    LocalMux I__11745 (
            .O(N__46645),
            .I(N__46589));
    Span4Mux_v I__11744 (
            .O(N__46642),
            .I(N__46589));
    InMux I__11743 (
            .O(N__46639),
            .I(N__46586));
    InMux I__11742 (
            .O(N__46638),
            .I(N__46583));
    LocalMux I__11741 (
            .O(N__46635),
            .I(N__46576));
    Span4Mux_v I__11740 (
            .O(N__46630),
            .I(N__46576));
    LocalMux I__11739 (
            .O(N__46627),
            .I(N__46576));
    InMux I__11738 (
            .O(N__46626),
            .I(N__46573));
    LocalMux I__11737 (
            .O(N__46623),
            .I(N__46570));
    InMux I__11736 (
            .O(N__46622),
            .I(N__46567));
    LocalMux I__11735 (
            .O(N__46617),
            .I(N__46564));
    InMux I__11734 (
            .O(N__46616),
            .I(N__46559));
    InMux I__11733 (
            .O(N__46615),
            .I(N__46559));
    Span4Mux_v I__11732 (
            .O(N__46612),
            .I(N__46556));
    Span4Mux_v I__11731 (
            .O(N__46609),
            .I(N__46551));
    LocalMux I__11730 (
            .O(N__46606),
            .I(N__46551));
    LocalMux I__11729 (
            .O(N__46603),
            .I(N__46546));
    Span4Mux_h I__11728 (
            .O(N__46600),
            .I(N__46546));
    Span4Mux_v I__11727 (
            .O(N__46597),
            .I(N__46543));
    LocalMux I__11726 (
            .O(N__46594),
            .I(N__46538));
    Span4Mux_h I__11725 (
            .O(N__46589),
            .I(N__46538));
    LocalMux I__11724 (
            .O(N__46586),
            .I(N__46535));
    LocalMux I__11723 (
            .O(N__46583),
            .I(N__46530));
    Span4Mux_v I__11722 (
            .O(N__46576),
            .I(N__46530));
    LocalMux I__11721 (
            .O(N__46573),
            .I(N__46525));
    Span4Mux_v I__11720 (
            .O(N__46570),
            .I(N__46525));
    LocalMux I__11719 (
            .O(N__46567),
            .I(N__46522));
    Span12Mux_v I__11718 (
            .O(N__46564),
            .I(N__46517));
    LocalMux I__11717 (
            .O(N__46559),
            .I(N__46517));
    Span4Mux_h I__11716 (
            .O(N__46556),
            .I(N__46512));
    Span4Mux_v I__11715 (
            .O(N__46551),
            .I(N__46512));
    Span4Mux_h I__11714 (
            .O(N__46546),
            .I(N__46509));
    Span4Mux_v I__11713 (
            .O(N__46543),
            .I(N__46504));
    Span4Mux_h I__11712 (
            .O(N__46538),
            .I(N__46504));
    Span4Mux_v I__11711 (
            .O(N__46535),
            .I(N__46495));
    Span4Mux_h I__11710 (
            .O(N__46530),
            .I(N__46495));
    Span4Mux_h I__11709 (
            .O(N__46525),
            .I(N__46495));
    Span4Mux_v I__11708 (
            .O(N__46522),
            .I(N__46495));
    Odrv12 I__11707 (
            .O(N__46517),
            .I(\ALU.aluOut_6 ));
    Odrv4 I__11706 (
            .O(N__46512),
            .I(\ALU.aluOut_6 ));
    Odrv4 I__11705 (
            .O(N__46509),
            .I(\ALU.aluOut_6 ));
    Odrv4 I__11704 (
            .O(N__46504),
            .I(\ALU.aluOut_6 ));
    Odrv4 I__11703 (
            .O(N__46495),
            .I(\ALU.aluOut_6 ));
    CascadeMux I__11702 (
            .O(N__46484),
            .I(\ALU.a_15_m2_ns_1Z0Z_6_cascade_ ));
    InMux I__11701 (
            .O(N__46481),
            .I(N__46478));
    LocalMux I__11700 (
            .O(N__46478),
            .I(N__46475));
    Span4Mux_v I__11699 (
            .O(N__46475),
            .I(N__46470));
    InMux I__11698 (
            .O(N__46474),
            .I(N__46467));
    InMux I__11697 (
            .O(N__46473),
            .I(N__46464));
    Span4Mux_h I__11696 (
            .O(N__46470),
            .I(N__46459));
    LocalMux I__11695 (
            .O(N__46467),
            .I(N__46456));
    LocalMux I__11694 (
            .O(N__46464),
            .I(N__46453));
    InMux I__11693 (
            .O(N__46463),
            .I(N__46450));
    InMux I__11692 (
            .O(N__46462),
            .I(N__46445));
    Span4Mux_h I__11691 (
            .O(N__46459),
            .I(N__46438));
    Span4Mux_v I__11690 (
            .O(N__46456),
            .I(N__46438));
    Span4Mux_h I__11689 (
            .O(N__46453),
            .I(N__46433));
    LocalMux I__11688 (
            .O(N__46450),
            .I(N__46433));
    InMux I__11687 (
            .O(N__46449),
            .I(N__46430));
    InMux I__11686 (
            .O(N__46448),
            .I(N__46427));
    LocalMux I__11685 (
            .O(N__46445),
            .I(N__46424));
    InMux I__11684 (
            .O(N__46444),
            .I(N__46421));
    InMux I__11683 (
            .O(N__46443),
            .I(N__46418));
    Span4Mux_v I__11682 (
            .O(N__46438),
            .I(N__46413));
    Span4Mux_v I__11681 (
            .O(N__46433),
            .I(N__46413));
    LocalMux I__11680 (
            .O(N__46430),
            .I(\ALU.N_219_0 ));
    LocalMux I__11679 (
            .O(N__46427),
            .I(\ALU.N_219_0 ));
    Odrv4 I__11678 (
            .O(N__46424),
            .I(\ALU.N_219_0 ));
    LocalMux I__11677 (
            .O(N__46421),
            .I(\ALU.N_219_0 ));
    LocalMux I__11676 (
            .O(N__46418),
            .I(\ALU.N_219_0 ));
    Odrv4 I__11675 (
            .O(N__46413),
            .I(\ALU.N_219_0 ));
    InMux I__11674 (
            .O(N__46400),
            .I(N__46397));
    LocalMux I__11673 (
            .O(N__46397),
            .I(\ALU.a_15_m2_6 ));
    InMux I__11672 (
            .O(N__46394),
            .I(N__46388));
    InMux I__11671 (
            .O(N__46393),
            .I(N__46385));
    InMux I__11670 (
            .O(N__46392),
            .I(N__46379));
    InMux I__11669 (
            .O(N__46391),
            .I(N__46376));
    LocalMux I__11668 (
            .O(N__46388),
            .I(N__46373));
    LocalMux I__11667 (
            .O(N__46385),
            .I(N__46370));
    InMux I__11666 (
            .O(N__46384),
            .I(N__46367));
    InMux I__11665 (
            .O(N__46383),
            .I(N__46364));
    InMux I__11664 (
            .O(N__46382),
            .I(N__46359));
    LocalMux I__11663 (
            .O(N__46379),
            .I(N__46354));
    LocalMux I__11662 (
            .O(N__46376),
            .I(N__46354));
    Span4Mux_v I__11661 (
            .O(N__46373),
            .I(N__46349));
    Span4Mux_h I__11660 (
            .O(N__46370),
            .I(N__46346));
    LocalMux I__11659 (
            .O(N__46367),
            .I(N__46343));
    LocalMux I__11658 (
            .O(N__46364),
            .I(N__46340));
    InMux I__11657 (
            .O(N__46363),
            .I(N__46335));
    InMux I__11656 (
            .O(N__46362),
            .I(N__46335));
    LocalMux I__11655 (
            .O(N__46359),
            .I(N__46332));
    Span4Mux_h I__11654 (
            .O(N__46354),
            .I(N__46327));
    InMux I__11653 (
            .O(N__46353),
            .I(N__46323));
    InMux I__11652 (
            .O(N__46352),
            .I(N__46320));
    Span4Mux_v I__11651 (
            .O(N__46349),
            .I(N__46317));
    Sp12to4 I__11650 (
            .O(N__46346),
            .I(N__46312));
    Span12Mux_h I__11649 (
            .O(N__46343),
            .I(N__46312));
    Span4Mux_v I__11648 (
            .O(N__46340),
            .I(N__46305));
    LocalMux I__11647 (
            .O(N__46335),
            .I(N__46305));
    Span4Mux_v I__11646 (
            .O(N__46332),
            .I(N__46302));
    InMux I__11645 (
            .O(N__46331),
            .I(N__46299));
    InMux I__11644 (
            .O(N__46330),
            .I(N__46296));
    Span4Mux_h I__11643 (
            .O(N__46327),
            .I(N__46293));
    InMux I__11642 (
            .O(N__46326),
            .I(N__46290));
    LocalMux I__11641 (
            .O(N__46323),
            .I(N__46285));
    LocalMux I__11640 (
            .O(N__46320),
            .I(N__46285));
    Sp12to4 I__11639 (
            .O(N__46317),
            .I(N__46280));
    Span12Mux_v I__11638 (
            .O(N__46312),
            .I(N__46280));
    InMux I__11637 (
            .O(N__46311),
            .I(N__46277));
    InMux I__11636 (
            .O(N__46310),
            .I(N__46274));
    IoSpan4Mux I__11635 (
            .O(N__46305),
            .I(N__46271));
    Span4Mux_h I__11634 (
            .O(N__46302),
            .I(N__46266));
    LocalMux I__11633 (
            .O(N__46299),
            .I(N__46266));
    LocalMux I__11632 (
            .O(N__46296),
            .I(N__46259));
    Span4Mux_v I__11631 (
            .O(N__46293),
            .I(N__46259));
    LocalMux I__11630 (
            .O(N__46290),
            .I(N__46259));
    Span12Mux_v I__11629 (
            .O(N__46285),
            .I(N__46256));
    Span12Mux_h I__11628 (
            .O(N__46280),
            .I(N__46253));
    LocalMux I__11627 (
            .O(N__46277),
            .I(N__46250));
    LocalMux I__11626 (
            .O(N__46274),
            .I(N__46245));
    IoSpan4Mux I__11625 (
            .O(N__46271),
            .I(N__46245));
    Span4Mux_v I__11624 (
            .O(N__46266),
            .I(N__46240));
    Span4Mux_v I__11623 (
            .O(N__46259),
            .I(N__46240));
    Odrv12 I__11622 (
            .O(N__46256),
            .I(\ALU.a_15_sm3 ));
    Odrv12 I__11621 (
            .O(N__46253),
            .I(\ALU.a_15_sm3 ));
    Odrv4 I__11620 (
            .O(N__46250),
            .I(\ALU.a_15_sm3 ));
    Odrv4 I__11619 (
            .O(N__46245),
            .I(\ALU.a_15_sm3 ));
    Odrv4 I__11618 (
            .O(N__46240),
            .I(\ALU.a_15_sm3 ));
    InMux I__11617 (
            .O(N__46229),
            .I(N__46226));
    LocalMux I__11616 (
            .O(N__46226),
            .I(N__46223));
    Span4Mux_h I__11615 (
            .O(N__46223),
            .I(N__46220));
    Span4Mux_h I__11614 (
            .O(N__46220),
            .I(N__46217));
    Span4Mux_h I__11613 (
            .O(N__46217),
            .I(N__46214));
    Span4Mux_v I__11612 (
            .O(N__46214),
            .I(N__46211));
    Odrv4 I__11611 (
            .O(N__46211),
            .I(\ALU.d_RNIL01TD1Z0Z_6 ));
    InMux I__11610 (
            .O(N__46208),
            .I(N__46205));
    LocalMux I__11609 (
            .O(N__46205),
            .I(\ALU.d_RNIJ75U41Z0Z_6 ));
    CascadeMux I__11608 (
            .O(N__46202),
            .I(N__46197));
    CascadeMux I__11607 (
            .O(N__46201),
            .I(N__46194));
    CascadeMux I__11606 (
            .O(N__46200),
            .I(N__46186));
    InMux I__11605 (
            .O(N__46197),
            .I(N__46181));
    InMux I__11604 (
            .O(N__46194),
            .I(N__46181));
    CascadeMux I__11603 (
            .O(N__46193),
            .I(N__46178));
    CascadeMux I__11602 (
            .O(N__46192),
            .I(N__46175));
    CascadeMux I__11601 (
            .O(N__46191),
            .I(N__46172));
    CascadeMux I__11600 (
            .O(N__46190),
            .I(N__46169));
    CascadeMux I__11599 (
            .O(N__46189),
            .I(N__46166));
    InMux I__11598 (
            .O(N__46186),
            .I(N__46144));
    LocalMux I__11597 (
            .O(N__46181),
            .I(N__46141));
    InMux I__11596 (
            .O(N__46178),
            .I(N__46138));
    InMux I__11595 (
            .O(N__46175),
            .I(N__46123));
    InMux I__11594 (
            .O(N__46172),
            .I(N__46123));
    InMux I__11593 (
            .O(N__46169),
            .I(N__46123));
    InMux I__11592 (
            .O(N__46166),
            .I(N__46123));
    InMux I__11591 (
            .O(N__46165),
            .I(N__46123));
    InMux I__11590 (
            .O(N__46164),
            .I(N__46123));
    InMux I__11589 (
            .O(N__46163),
            .I(N__46123));
    CascadeMux I__11588 (
            .O(N__46162),
            .I(N__46119));
    CascadeMux I__11587 (
            .O(N__46161),
            .I(N__46114));
    CascadeMux I__11586 (
            .O(N__46160),
            .I(N__46111));
    CascadeMux I__11585 (
            .O(N__46159),
            .I(N__46108));
    CascadeMux I__11584 (
            .O(N__46158),
            .I(N__46105));
    CascadeMux I__11583 (
            .O(N__46157),
            .I(N__46102));
    CascadeMux I__11582 (
            .O(N__46156),
            .I(N__46099));
    CascadeMux I__11581 (
            .O(N__46155),
            .I(N__46095));
    CascadeMux I__11580 (
            .O(N__46154),
            .I(N__46092));
    CascadeMux I__11579 (
            .O(N__46153),
            .I(N__46089));
    CascadeMux I__11578 (
            .O(N__46152),
            .I(N__46086));
    CascadeMux I__11577 (
            .O(N__46151),
            .I(N__46073));
    CascadeMux I__11576 (
            .O(N__46150),
            .I(N__46070));
    CascadeMux I__11575 (
            .O(N__46149),
            .I(N__46067));
    CascadeMux I__11574 (
            .O(N__46148),
            .I(N__46064));
    CascadeMux I__11573 (
            .O(N__46147),
            .I(N__46061));
    LocalMux I__11572 (
            .O(N__46144),
            .I(N__46057));
    Span4Mux_h I__11571 (
            .O(N__46141),
            .I(N__46050));
    LocalMux I__11570 (
            .O(N__46138),
            .I(N__46050));
    LocalMux I__11569 (
            .O(N__46123),
            .I(N__46050));
    CascadeMux I__11568 (
            .O(N__46122),
            .I(N__46047));
    InMux I__11567 (
            .O(N__46119),
            .I(N__46042));
    CascadeMux I__11566 (
            .O(N__46118),
            .I(N__46037));
    CascadeMux I__11565 (
            .O(N__46117),
            .I(N__46034));
    InMux I__11564 (
            .O(N__46114),
            .I(N__46024));
    InMux I__11563 (
            .O(N__46111),
            .I(N__46024));
    InMux I__11562 (
            .O(N__46108),
            .I(N__46024));
    InMux I__11561 (
            .O(N__46105),
            .I(N__46024));
    InMux I__11560 (
            .O(N__46102),
            .I(N__46017));
    InMux I__11559 (
            .O(N__46099),
            .I(N__46017));
    InMux I__11558 (
            .O(N__46098),
            .I(N__46017));
    InMux I__11557 (
            .O(N__46095),
            .I(N__46008));
    InMux I__11556 (
            .O(N__46092),
            .I(N__46008));
    InMux I__11555 (
            .O(N__46089),
            .I(N__46008));
    InMux I__11554 (
            .O(N__46086),
            .I(N__46008));
    InMux I__11553 (
            .O(N__46085),
            .I(N__46005));
    CascadeMux I__11552 (
            .O(N__46084),
            .I(N__45997));
    CascadeMux I__11551 (
            .O(N__46083),
            .I(N__45994));
    CascadeMux I__11550 (
            .O(N__46082),
            .I(N__45986));
    CascadeMux I__11549 (
            .O(N__46081),
            .I(N__45983));
    CascadeMux I__11548 (
            .O(N__46080),
            .I(N__45980));
    CascadeMux I__11547 (
            .O(N__46079),
            .I(N__45977));
    CascadeMux I__11546 (
            .O(N__46078),
            .I(N__45974));
    CascadeMux I__11545 (
            .O(N__46077),
            .I(N__45971));
    CascadeMux I__11544 (
            .O(N__46076),
            .I(N__45968));
    InMux I__11543 (
            .O(N__46073),
            .I(N__45962));
    InMux I__11542 (
            .O(N__46070),
            .I(N__45962));
    InMux I__11541 (
            .O(N__46067),
            .I(N__45953));
    InMux I__11540 (
            .O(N__46064),
            .I(N__45953));
    InMux I__11539 (
            .O(N__46061),
            .I(N__45953));
    InMux I__11538 (
            .O(N__46060),
            .I(N__45953));
    Span4Mux_h I__11537 (
            .O(N__46057),
            .I(N__45950));
    Span4Mux_v I__11536 (
            .O(N__46050),
            .I(N__45947));
    InMux I__11535 (
            .O(N__46047),
            .I(N__45940));
    InMux I__11534 (
            .O(N__46046),
            .I(N__45940));
    InMux I__11533 (
            .O(N__46045),
            .I(N__45940));
    LocalMux I__11532 (
            .O(N__46042),
            .I(N__45937));
    InMux I__11531 (
            .O(N__46041),
            .I(N__45934));
    InMux I__11530 (
            .O(N__46040),
            .I(N__45931));
    InMux I__11529 (
            .O(N__46037),
            .I(N__45927));
    InMux I__11528 (
            .O(N__46034),
            .I(N__45924));
    InMux I__11527 (
            .O(N__46033),
            .I(N__45920));
    LocalMux I__11526 (
            .O(N__46024),
            .I(N__45913));
    LocalMux I__11525 (
            .O(N__46017),
            .I(N__45913));
    LocalMux I__11524 (
            .O(N__46008),
            .I(N__45913));
    LocalMux I__11523 (
            .O(N__46005),
            .I(N__45910));
    InMux I__11522 (
            .O(N__46004),
            .I(N__45907));
    InMux I__11521 (
            .O(N__46003),
            .I(N__45904));
    CascadeMux I__11520 (
            .O(N__46002),
            .I(N__45900));
    CascadeMux I__11519 (
            .O(N__46001),
            .I(N__45897));
    CascadeMux I__11518 (
            .O(N__46000),
            .I(N__45894));
    InMux I__11517 (
            .O(N__45997),
            .I(N__45886));
    InMux I__11516 (
            .O(N__45994),
            .I(N__45886));
    InMux I__11515 (
            .O(N__45993),
            .I(N__45886));
    InMux I__11514 (
            .O(N__45992),
            .I(N__45883));
    CascadeMux I__11513 (
            .O(N__45991),
            .I(N__45880));
    InMux I__11512 (
            .O(N__45990),
            .I(N__45877));
    CascadeMux I__11511 (
            .O(N__45989),
            .I(N__45874));
    InMux I__11510 (
            .O(N__45986),
            .I(N__45866));
    InMux I__11509 (
            .O(N__45983),
            .I(N__45866));
    InMux I__11508 (
            .O(N__45980),
            .I(N__45866));
    InMux I__11507 (
            .O(N__45977),
            .I(N__45857));
    InMux I__11506 (
            .O(N__45974),
            .I(N__45857));
    InMux I__11505 (
            .O(N__45971),
            .I(N__45857));
    InMux I__11504 (
            .O(N__45968),
            .I(N__45857));
    InMux I__11503 (
            .O(N__45967),
            .I(N__45854));
    LocalMux I__11502 (
            .O(N__45962),
            .I(N__45843));
    LocalMux I__11501 (
            .O(N__45953),
            .I(N__45843));
    Span4Mux_h I__11500 (
            .O(N__45950),
            .I(N__45843));
    Span4Mux_v I__11499 (
            .O(N__45947),
            .I(N__45843));
    LocalMux I__11498 (
            .O(N__45940),
            .I(N__45843));
    Span4Mux_h I__11497 (
            .O(N__45937),
            .I(N__45837));
    LocalMux I__11496 (
            .O(N__45934),
            .I(N__45837));
    LocalMux I__11495 (
            .O(N__45931),
            .I(N__45833));
    InMux I__11494 (
            .O(N__45930),
            .I(N__45830));
    LocalMux I__11493 (
            .O(N__45927),
            .I(N__45825));
    LocalMux I__11492 (
            .O(N__45924),
            .I(N__45825));
    InMux I__11491 (
            .O(N__45923),
            .I(N__45822));
    LocalMux I__11490 (
            .O(N__45920),
            .I(N__45819));
    Span4Mux_h I__11489 (
            .O(N__45913),
            .I(N__45816));
    Span4Mux_v I__11488 (
            .O(N__45910),
            .I(N__45813));
    LocalMux I__11487 (
            .O(N__45907),
            .I(N__45808));
    LocalMux I__11486 (
            .O(N__45904),
            .I(N__45808));
    InMux I__11485 (
            .O(N__45903),
            .I(N__45805));
    InMux I__11484 (
            .O(N__45900),
            .I(N__45798));
    InMux I__11483 (
            .O(N__45897),
            .I(N__45798));
    InMux I__11482 (
            .O(N__45894),
            .I(N__45798));
    InMux I__11481 (
            .O(N__45893),
            .I(N__45795));
    LocalMux I__11480 (
            .O(N__45886),
            .I(N__45790));
    LocalMux I__11479 (
            .O(N__45883),
            .I(N__45790));
    InMux I__11478 (
            .O(N__45880),
            .I(N__45787));
    LocalMux I__11477 (
            .O(N__45877),
            .I(N__45784));
    InMux I__11476 (
            .O(N__45874),
            .I(N__45781));
    CascadeMux I__11475 (
            .O(N__45873),
            .I(N__45778));
    LocalMux I__11474 (
            .O(N__45866),
            .I(N__45769));
    LocalMux I__11473 (
            .O(N__45857),
            .I(N__45769));
    LocalMux I__11472 (
            .O(N__45854),
            .I(N__45769));
    Span4Mux_v I__11471 (
            .O(N__45843),
            .I(N__45769));
    InMux I__11470 (
            .O(N__45842),
            .I(N__45766));
    Span4Mux_v I__11469 (
            .O(N__45837),
            .I(N__45763));
    InMux I__11468 (
            .O(N__45836),
            .I(N__45760));
    Span4Mux_h I__11467 (
            .O(N__45833),
            .I(N__45751));
    LocalMux I__11466 (
            .O(N__45830),
            .I(N__45751));
    Span4Mux_v I__11465 (
            .O(N__45825),
            .I(N__45751));
    LocalMux I__11464 (
            .O(N__45822),
            .I(N__45751));
    Span4Mux_v I__11463 (
            .O(N__45819),
            .I(N__45748));
    Span4Mux_h I__11462 (
            .O(N__45816),
            .I(N__45741));
    Span4Mux_h I__11461 (
            .O(N__45813),
            .I(N__45741));
    Span4Mux_v I__11460 (
            .O(N__45808),
            .I(N__45741));
    LocalMux I__11459 (
            .O(N__45805),
            .I(N__45734));
    LocalMux I__11458 (
            .O(N__45798),
            .I(N__45734));
    LocalMux I__11457 (
            .O(N__45795),
            .I(N__45734));
    Span4Mux_h I__11456 (
            .O(N__45790),
            .I(N__45731));
    LocalMux I__11455 (
            .O(N__45787),
            .I(N__45724));
    Span4Mux_h I__11454 (
            .O(N__45784),
            .I(N__45724));
    LocalMux I__11453 (
            .O(N__45781),
            .I(N__45724));
    InMux I__11452 (
            .O(N__45778),
            .I(N__45721));
    Span4Mux_h I__11451 (
            .O(N__45769),
            .I(N__45718));
    LocalMux I__11450 (
            .O(N__45766),
            .I(N__45713));
    Span4Mux_h I__11449 (
            .O(N__45763),
            .I(N__45713));
    LocalMux I__11448 (
            .O(N__45760),
            .I(N__45710));
    Span4Mux_v I__11447 (
            .O(N__45751),
            .I(N__45705));
    Span4Mux_v I__11446 (
            .O(N__45748),
            .I(N__45705));
    Span4Mux_v I__11445 (
            .O(N__45741),
            .I(N__45700));
    Span4Mux_v I__11444 (
            .O(N__45734),
            .I(N__45700));
    Span4Mux_v I__11443 (
            .O(N__45731),
            .I(N__45692));
    Span4Mux_v I__11442 (
            .O(N__45724),
            .I(N__45692));
    LocalMux I__11441 (
            .O(N__45721),
            .I(N__45685));
    Span4Mux_h I__11440 (
            .O(N__45718),
            .I(N__45685));
    Span4Mux_v I__11439 (
            .O(N__45713),
            .I(N__45685));
    Span4Mux_v I__11438 (
            .O(N__45710),
            .I(N__45680));
    Span4Mux_h I__11437 (
            .O(N__45705),
            .I(N__45680));
    Span4Mux_v I__11436 (
            .O(N__45700),
            .I(N__45677));
    InMux I__11435 (
            .O(N__45699),
            .I(N__45674));
    InMux I__11434 (
            .O(N__45698),
            .I(N__45671));
    InMux I__11433 (
            .O(N__45697),
            .I(N__45668));
    Span4Mux_h I__11432 (
            .O(N__45692),
            .I(N__45665));
    Span4Mux_v I__11431 (
            .O(N__45685),
            .I(N__45662));
    Span4Mux_h I__11430 (
            .O(N__45680),
            .I(N__45659));
    Span4Mux_h I__11429 (
            .O(N__45677),
            .I(N__45656));
    LocalMux I__11428 (
            .O(N__45674),
            .I(N__45653));
    LocalMux I__11427 (
            .O(N__45671),
            .I(aluOperation_1));
    LocalMux I__11426 (
            .O(N__45668),
            .I(aluOperation_1));
    Odrv4 I__11425 (
            .O(N__45665),
            .I(aluOperation_1));
    Odrv4 I__11424 (
            .O(N__45662),
            .I(aluOperation_1));
    Odrv4 I__11423 (
            .O(N__45659),
            .I(aluOperation_1));
    Odrv4 I__11422 (
            .O(N__45656),
            .I(aluOperation_1));
    Odrv4 I__11421 (
            .O(N__45653),
            .I(aluOperation_1));
    CascadeMux I__11420 (
            .O(N__45638),
            .I(\ALU.a_15_m5_6_cascade_ ));
    InMux I__11419 (
            .O(N__45635),
            .I(N__45632));
    LocalMux I__11418 (
            .O(N__45632),
            .I(N__45629));
    Odrv12 I__11417 (
            .O(N__45629),
            .I(\ALU.mult_6 ));
    CascadeMux I__11416 (
            .O(N__45626),
            .I(\ALU.d_RNILPR7TQZ0Z_6_cascade_ ));
    InMux I__11415 (
            .O(N__45623),
            .I(N__45619));
    CascadeMux I__11414 (
            .O(N__45622),
            .I(N__45616));
    LocalMux I__11413 (
            .O(N__45619),
            .I(N__45613));
    InMux I__11412 (
            .O(N__45616),
            .I(N__45610));
    Span4Mux_h I__11411 (
            .O(N__45613),
            .I(N__45607));
    LocalMux I__11410 (
            .O(N__45610),
            .I(N__45604));
    Span4Mux_h I__11409 (
            .O(N__45607),
            .I(N__45601));
    Span4Mux_v I__11408 (
            .O(N__45604),
            .I(N__45598));
    Span4Mux_v I__11407 (
            .O(N__45601),
            .I(N__45595));
    Span4Mux_h I__11406 (
            .O(N__45598),
            .I(N__45592));
    Odrv4 I__11405 (
            .O(N__45595),
            .I(\ALU.hZ0Z_6 ));
    Odrv4 I__11404 (
            .O(N__45592),
            .I(\ALU.hZ0Z_6 ));
    CEMux I__11403 (
            .O(N__45587),
            .I(N__45583));
    CEMux I__11402 (
            .O(N__45586),
            .I(N__45580));
    LocalMux I__11401 (
            .O(N__45583),
            .I(N__45575));
    LocalMux I__11400 (
            .O(N__45580),
            .I(N__45575));
    Span4Mux_v I__11399 (
            .O(N__45575),
            .I(N__45569));
    CEMux I__11398 (
            .O(N__45574),
            .I(N__45564));
    CEMux I__11397 (
            .O(N__45573),
            .I(N__45561));
    CEMux I__11396 (
            .O(N__45572),
            .I(N__45558));
    Span4Mux_h I__11395 (
            .O(N__45569),
            .I(N__45554));
    CEMux I__11394 (
            .O(N__45568),
            .I(N__45551));
    CEMux I__11393 (
            .O(N__45567),
            .I(N__45548));
    LocalMux I__11392 (
            .O(N__45564),
            .I(N__45545));
    LocalMux I__11391 (
            .O(N__45561),
            .I(N__45542));
    LocalMux I__11390 (
            .O(N__45558),
            .I(N__45539));
    CEMux I__11389 (
            .O(N__45557),
            .I(N__45535));
    Span4Mux_v I__11388 (
            .O(N__45554),
            .I(N__45532));
    LocalMux I__11387 (
            .O(N__45551),
            .I(N__45529));
    LocalMux I__11386 (
            .O(N__45548),
            .I(N__45526));
    Span4Mux_h I__11385 (
            .O(N__45545),
            .I(N__45522));
    Span4Mux_v I__11384 (
            .O(N__45542),
            .I(N__45517));
    Span4Mux_h I__11383 (
            .O(N__45539),
            .I(N__45517));
    CEMux I__11382 (
            .O(N__45538),
            .I(N__45514));
    LocalMux I__11381 (
            .O(N__45535),
            .I(N__45511));
    Span4Mux_v I__11380 (
            .O(N__45532),
            .I(N__45508));
    Span4Mux_h I__11379 (
            .O(N__45529),
            .I(N__45505));
    Span4Mux_v I__11378 (
            .O(N__45526),
            .I(N__45502));
    CEMux I__11377 (
            .O(N__45525),
            .I(N__45499));
    Span4Mux_v I__11376 (
            .O(N__45522),
            .I(N__45495));
    Span4Mux_v I__11375 (
            .O(N__45517),
            .I(N__45490));
    LocalMux I__11374 (
            .O(N__45514),
            .I(N__45490));
    Span4Mux_v I__11373 (
            .O(N__45511),
            .I(N__45486));
    IoSpan4Mux I__11372 (
            .O(N__45508),
            .I(N__45483));
    Span4Mux_v I__11371 (
            .O(N__45505),
            .I(N__45476));
    Span4Mux_h I__11370 (
            .O(N__45502),
            .I(N__45476));
    LocalMux I__11369 (
            .O(N__45499),
            .I(N__45476));
    CEMux I__11368 (
            .O(N__45498),
            .I(N__45473));
    Span4Mux_v I__11367 (
            .O(N__45495),
            .I(N__45468));
    Span4Mux_h I__11366 (
            .O(N__45490),
            .I(N__45468));
    CEMux I__11365 (
            .O(N__45489),
            .I(N__45465));
    Span4Mux_v I__11364 (
            .O(N__45486),
            .I(N__45462));
    Span4Mux_s2_v I__11363 (
            .O(N__45483),
            .I(N__45459));
    Span4Mux_h I__11362 (
            .O(N__45476),
            .I(N__45456));
    LocalMux I__11361 (
            .O(N__45473),
            .I(N__45453));
    Span4Mux_h I__11360 (
            .O(N__45468),
            .I(N__45450));
    LocalMux I__11359 (
            .O(N__45465),
            .I(N__45447));
    Span4Mux_h I__11358 (
            .O(N__45462),
            .I(N__45444));
    Span4Mux_s2_h I__11357 (
            .O(N__45459),
            .I(N__45439));
    Span4Mux_v I__11356 (
            .O(N__45456),
            .I(N__45439));
    Span4Mux_v I__11355 (
            .O(N__45453),
            .I(N__45436));
    Span4Mux_s3_h I__11354 (
            .O(N__45450),
            .I(N__45431));
    Span4Mux_h I__11353 (
            .O(N__45447),
            .I(N__45431));
    Span4Mux_h I__11352 (
            .O(N__45444),
            .I(N__45428));
    Span4Mux_h I__11351 (
            .O(N__45439),
            .I(N__45425));
    Span4Mux_h I__11350 (
            .O(N__45436),
            .I(N__45422));
    Span4Mux_v I__11349 (
            .O(N__45431),
            .I(N__45419));
    Odrv4 I__11348 (
            .O(N__45428),
            .I(\ALU.h_cnvZ0Z_0 ));
    Odrv4 I__11347 (
            .O(N__45425),
            .I(\ALU.h_cnvZ0Z_0 ));
    Odrv4 I__11346 (
            .O(N__45422),
            .I(\ALU.h_cnvZ0Z_0 ));
    Odrv4 I__11345 (
            .O(N__45419),
            .I(\ALU.h_cnvZ0Z_0 ));
    InMux I__11344 (
            .O(N__45410),
            .I(N__45406));
    InMux I__11343 (
            .O(N__45409),
            .I(N__45403));
    LocalMux I__11342 (
            .O(N__45406),
            .I(N__45400));
    LocalMux I__11341 (
            .O(N__45403),
            .I(N__45397));
    Span4Mux_h I__11340 (
            .O(N__45400),
            .I(N__45392));
    Span4Mux_h I__11339 (
            .O(N__45397),
            .I(N__45392));
    Odrv4 I__11338 (
            .O(N__45392),
            .I(\ALU.fZ0Z_4 ));
    InMux I__11337 (
            .O(N__45389),
            .I(N__45386));
    LocalMux I__11336 (
            .O(N__45386),
            .I(N__45383));
    Span4Mux_h I__11335 (
            .O(N__45383),
            .I(N__45380));
    Span4Mux_h I__11334 (
            .O(N__45380),
            .I(N__45377));
    Odrv4 I__11333 (
            .O(N__45377),
            .I(\ALU.f_RNIJ0FJZ0Z_4 ));
    InMux I__11332 (
            .O(N__45374),
            .I(N__45370));
    InMux I__11331 (
            .O(N__45373),
            .I(N__45367));
    LocalMux I__11330 (
            .O(N__45370),
            .I(N__45364));
    LocalMux I__11329 (
            .O(N__45367),
            .I(N__45359));
    Span12Mux_v I__11328 (
            .O(N__45364),
            .I(N__45359));
    Odrv12 I__11327 (
            .O(N__45359),
            .I(\ALU.hZ0Z_7 ));
    InMux I__11326 (
            .O(N__45356),
            .I(N__45353));
    LocalMux I__11325 (
            .O(N__45353),
            .I(N__45350));
    Span12Mux_s9_h I__11324 (
            .O(N__45350),
            .I(N__45346));
    InMux I__11323 (
            .O(N__45349),
            .I(N__45343));
    Odrv12 I__11322 (
            .O(N__45346),
            .I(\ALU.dZ0Z_7 ));
    LocalMux I__11321 (
            .O(N__45343),
            .I(\ALU.dZ0Z_7 ));
    InMux I__11320 (
            .O(N__45338),
            .I(N__45330));
    InMux I__11319 (
            .O(N__45337),
            .I(N__45323));
    InMux I__11318 (
            .O(N__45336),
            .I(N__45323));
    InMux I__11317 (
            .O(N__45335),
            .I(N__45323));
    InMux I__11316 (
            .O(N__45334),
            .I(N__45318));
    InMux I__11315 (
            .O(N__45333),
            .I(N__45315));
    LocalMux I__11314 (
            .O(N__45330),
            .I(N__45309));
    LocalMux I__11313 (
            .O(N__45323),
            .I(N__45306));
    InMux I__11312 (
            .O(N__45322),
            .I(N__45303));
    InMux I__11311 (
            .O(N__45321),
            .I(N__45300));
    LocalMux I__11310 (
            .O(N__45318),
            .I(N__45296));
    LocalMux I__11309 (
            .O(N__45315),
            .I(N__45293));
    InMux I__11308 (
            .O(N__45314),
            .I(N__45288));
    InMux I__11307 (
            .O(N__45313),
            .I(N__45288));
    InMux I__11306 (
            .O(N__45312),
            .I(N__45285));
    Span4Mux_v I__11305 (
            .O(N__45309),
            .I(N__45270));
    Span4Mux_v I__11304 (
            .O(N__45306),
            .I(N__45270));
    LocalMux I__11303 (
            .O(N__45303),
            .I(N__45265));
    LocalMux I__11302 (
            .O(N__45300),
            .I(N__45265));
    InMux I__11301 (
            .O(N__45299),
            .I(N__45262));
    Span4Mux_h I__11300 (
            .O(N__45296),
            .I(N__45255));
    Span4Mux_v I__11299 (
            .O(N__45293),
            .I(N__45255));
    LocalMux I__11298 (
            .O(N__45288),
            .I(N__45255));
    LocalMux I__11297 (
            .O(N__45285),
            .I(N__45252));
    InMux I__11296 (
            .O(N__45284),
            .I(N__45247));
    InMux I__11295 (
            .O(N__45283),
            .I(N__45247));
    InMux I__11294 (
            .O(N__45282),
            .I(N__45242));
    InMux I__11293 (
            .O(N__45281),
            .I(N__45242));
    InMux I__11292 (
            .O(N__45280),
            .I(N__45231));
    InMux I__11291 (
            .O(N__45279),
            .I(N__45231));
    InMux I__11290 (
            .O(N__45278),
            .I(N__45231));
    InMux I__11289 (
            .O(N__45277),
            .I(N__45231));
    InMux I__11288 (
            .O(N__45276),
            .I(N__45231));
    InMux I__11287 (
            .O(N__45275),
            .I(N__45228));
    Span4Mux_v I__11286 (
            .O(N__45270),
            .I(N__45223));
    Span4Mux_v I__11285 (
            .O(N__45265),
            .I(N__45223));
    LocalMux I__11284 (
            .O(N__45262),
            .I(N__45216));
    Span4Mux_v I__11283 (
            .O(N__45255),
            .I(N__45216));
    Span4Mux_v I__11282 (
            .O(N__45252),
            .I(N__45216));
    LocalMux I__11281 (
            .O(N__45247),
            .I(aluOperand2_2));
    LocalMux I__11280 (
            .O(N__45242),
            .I(aluOperand2_2));
    LocalMux I__11279 (
            .O(N__45231),
            .I(aluOperand2_2));
    LocalMux I__11278 (
            .O(N__45228),
            .I(aluOperand2_2));
    Odrv4 I__11277 (
            .O(N__45223),
            .I(aluOperand2_2));
    Odrv4 I__11276 (
            .O(N__45216),
            .I(aluOperand2_2));
    InMux I__11275 (
            .O(N__45203),
            .I(N__45200));
    LocalMux I__11274 (
            .O(N__45200),
            .I(N__45197));
    Span4Mux_h I__11273 (
            .O(N__45197),
            .I(N__45194));
    Span4Mux_h I__11272 (
            .O(N__45194),
            .I(N__45191));
    Span4Mux_h I__11271 (
            .O(N__45191),
            .I(N__45188));
    Odrv4 I__11270 (
            .O(N__45188),
            .I(\ALU.d_RNIU60LZ0Z_7 ));
    CascadeMux I__11269 (
            .O(N__45185),
            .I(N__45182));
    InMux I__11268 (
            .O(N__45182),
            .I(N__45179));
    LocalMux I__11267 (
            .O(N__45179),
            .I(N__45176));
    Span4Mux_h I__11266 (
            .O(N__45176),
            .I(N__45172));
    InMux I__11265 (
            .O(N__45175),
            .I(N__45169));
    Span4Mux_h I__11264 (
            .O(N__45172),
            .I(N__45166));
    LocalMux I__11263 (
            .O(N__45169),
            .I(N__45163));
    Odrv4 I__11262 (
            .O(N__45166),
            .I(\ALU.hZ0Z_3 ));
    Odrv4 I__11261 (
            .O(N__45163),
            .I(\ALU.hZ0Z_3 ));
    InMux I__11260 (
            .O(N__45158),
            .I(N__45155));
    LocalMux I__11259 (
            .O(N__45155),
            .I(N__45152));
    Span4Mux_v I__11258 (
            .O(N__45152),
            .I(N__45149));
    Span4Mux_h I__11257 (
            .O(N__45149),
            .I(N__45145));
    InMux I__11256 (
            .O(N__45148),
            .I(N__45142));
    Odrv4 I__11255 (
            .O(N__45145),
            .I(\ALU.dZ0Z_3 ));
    LocalMux I__11254 (
            .O(N__45142),
            .I(\ALU.dZ0Z_3 ));
    InMux I__11253 (
            .O(N__45137),
            .I(N__45130));
    InMux I__11252 (
            .O(N__45136),
            .I(N__45130));
    CascadeMux I__11251 (
            .O(N__45135),
            .I(N__45123));
    LocalMux I__11250 (
            .O(N__45130),
            .I(N__45116));
    InMux I__11249 (
            .O(N__45129),
            .I(N__45113));
    InMux I__11248 (
            .O(N__45128),
            .I(N__45109));
    InMux I__11247 (
            .O(N__45127),
            .I(N__45104));
    InMux I__11246 (
            .O(N__45126),
            .I(N__45104));
    InMux I__11245 (
            .O(N__45123),
            .I(N__45100));
    InMux I__11244 (
            .O(N__45122),
            .I(N__45097));
    InMux I__11243 (
            .O(N__45121),
            .I(N__45094));
    InMux I__11242 (
            .O(N__45120),
            .I(N__45091));
    InMux I__11241 (
            .O(N__45119),
            .I(N__45088));
    Span4Mux_v I__11240 (
            .O(N__45116),
            .I(N__45085));
    LocalMux I__11239 (
            .O(N__45113),
            .I(N__45082));
    InMux I__11238 (
            .O(N__45112),
            .I(N__45073));
    LocalMux I__11237 (
            .O(N__45109),
            .I(N__45070));
    LocalMux I__11236 (
            .O(N__45104),
            .I(N__45067));
    InMux I__11235 (
            .O(N__45103),
            .I(N__45064));
    LocalMux I__11234 (
            .O(N__45100),
            .I(N__45060));
    LocalMux I__11233 (
            .O(N__45097),
            .I(N__45057));
    LocalMux I__11232 (
            .O(N__45094),
            .I(N__45050));
    LocalMux I__11231 (
            .O(N__45091),
            .I(N__45050));
    LocalMux I__11230 (
            .O(N__45088),
            .I(N__45050));
    Span4Mux_s3_h I__11229 (
            .O(N__45085),
            .I(N__45047));
    Span4Mux_h I__11228 (
            .O(N__45082),
            .I(N__45044));
    InMux I__11227 (
            .O(N__45081),
            .I(N__45041));
    InMux I__11226 (
            .O(N__45080),
            .I(N__45030));
    InMux I__11225 (
            .O(N__45079),
            .I(N__45030));
    InMux I__11224 (
            .O(N__45078),
            .I(N__45030));
    InMux I__11223 (
            .O(N__45077),
            .I(N__45030));
    InMux I__11222 (
            .O(N__45076),
            .I(N__45030));
    LocalMux I__11221 (
            .O(N__45073),
            .I(N__45027));
    Span4Mux_v I__11220 (
            .O(N__45070),
            .I(N__45022));
    Span4Mux_h I__11219 (
            .O(N__45067),
            .I(N__45022));
    LocalMux I__11218 (
            .O(N__45064),
            .I(N__45019));
    InMux I__11217 (
            .O(N__45063),
            .I(N__45016));
    Span4Mux_v I__11216 (
            .O(N__45060),
            .I(N__45009));
    Span4Mux_v I__11215 (
            .O(N__45057),
            .I(N__45009));
    Span4Mux_v I__11214 (
            .O(N__45050),
            .I(N__45009));
    Span4Mux_h I__11213 (
            .O(N__45047),
            .I(N__45004));
    Span4Mux_v I__11212 (
            .O(N__45044),
            .I(N__45004));
    LocalMux I__11211 (
            .O(N__45041),
            .I(aluOperand2_2_rep2));
    LocalMux I__11210 (
            .O(N__45030),
            .I(aluOperand2_2_rep2));
    Odrv4 I__11209 (
            .O(N__45027),
            .I(aluOperand2_2_rep2));
    Odrv4 I__11208 (
            .O(N__45022),
            .I(aluOperand2_2_rep2));
    Odrv4 I__11207 (
            .O(N__45019),
            .I(aluOperand2_2_rep2));
    LocalMux I__11206 (
            .O(N__45016),
            .I(aluOperand2_2_rep2));
    Odrv4 I__11205 (
            .O(N__45009),
            .I(aluOperand2_2_rep2));
    Odrv4 I__11204 (
            .O(N__45004),
            .I(aluOperand2_2_rep2));
    InMux I__11203 (
            .O(N__44987),
            .I(N__44984));
    LocalMux I__11202 (
            .O(N__44984),
            .I(N__44981));
    Span4Mux_h I__11201 (
            .O(N__44981),
            .I(N__44978));
    Span4Mux_h I__11200 (
            .O(N__44978),
            .I(N__44975));
    Odrv4 I__11199 (
            .O(N__44975),
            .I(\ALU.d_RNILAR7Z0Z_3 ));
    CascadeMux I__11198 (
            .O(N__44972),
            .I(\ALU.a_15_m2_4_cascade_ ));
    InMux I__11197 (
            .O(N__44969),
            .I(N__44966));
    LocalMux I__11196 (
            .O(N__44966),
            .I(N__44963));
    Span4Mux_v I__11195 (
            .O(N__44963),
            .I(N__44960));
    Span4Mux_v I__11194 (
            .O(N__44960),
            .I(N__44956));
    InMux I__11193 (
            .O(N__44959),
            .I(N__44953));
    Span4Mux_h I__11192 (
            .O(N__44956),
            .I(N__44950));
    LocalMux I__11191 (
            .O(N__44953),
            .I(N__44947));
    Odrv4 I__11190 (
            .O(N__44950),
            .I(\ALU.N_419 ));
    Odrv4 I__11189 (
            .O(N__44947),
            .I(\ALU.N_419 ));
    InMux I__11188 (
            .O(N__44942),
            .I(N__44939));
    LocalMux I__11187 (
            .O(N__44939),
            .I(\ALU.a_15_m4_4 ));
    InMux I__11186 (
            .O(N__44936),
            .I(N__44933));
    LocalMux I__11185 (
            .O(N__44933),
            .I(N__44930));
    Sp12to4 I__11184 (
            .O(N__44930),
            .I(N__44927));
    Span12Mux_v I__11183 (
            .O(N__44927),
            .I(N__44924));
    Odrv12 I__11182 (
            .O(N__44924),
            .I(\ALU.mult_4 ));
    InMux I__11181 (
            .O(N__44921),
            .I(N__44918));
    LocalMux I__11180 (
            .O(N__44918),
            .I(\ALU.a_15_m5_4 ));
    InMux I__11179 (
            .O(N__44915),
            .I(N__44912));
    LocalMux I__11178 (
            .O(N__44912),
            .I(N__44909));
    Span4Mux_h I__11177 (
            .O(N__44909),
            .I(N__44904));
    InMux I__11176 (
            .O(N__44908),
            .I(N__44899));
    InMux I__11175 (
            .O(N__44907),
            .I(N__44899));
    Sp12to4 I__11174 (
            .O(N__44904),
            .I(N__44896));
    LocalMux I__11173 (
            .O(N__44899),
            .I(N__44893));
    Odrv12 I__11172 (
            .O(N__44896),
            .I(a_3));
    Odrv12 I__11171 (
            .O(N__44893),
            .I(a_3));
    CEMux I__11170 (
            .O(N__44888),
            .I(N__44885));
    LocalMux I__11169 (
            .O(N__44885),
            .I(N__44881));
    CEMux I__11168 (
            .O(N__44884),
            .I(N__44878));
    Span4Mux_h I__11167 (
            .O(N__44881),
            .I(N__44873));
    LocalMux I__11166 (
            .O(N__44878),
            .I(N__44873));
    Span4Mux_v I__11165 (
            .O(N__44873),
            .I(N__44867));
    CEMux I__11164 (
            .O(N__44872),
            .I(N__44864));
    CEMux I__11163 (
            .O(N__44871),
            .I(N__44861));
    CEMux I__11162 (
            .O(N__44870),
            .I(N__44858));
    Span4Mux_v I__11161 (
            .O(N__44867),
            .I(N__44853));
    LocalMux I__11160 (
            .O(N__44864),
            .I(N__44853));
    LocalMux I__11159 (
            .O(N__44861),
            .I(N__44850));
    LocalMux I__11158 (
            .O(N__44858),
            .I(N__44846));
    Span4Mux_v I__11157 (
            .O(N__44853),
            .I(N__44841));
    Span4Mux_v I__11156 (
            .O(N__44850),
            .I(N__44841));
    CEMux I__11155 (
            .O(N__44849),
            .I(N__44838));
    Span4Mux_h I__11154 (
            .O(N__44846),
            .I(N__44834));
    IoSpan4Mux I__11153 (
            .O(N__44841),
            .I(N__44831));
    LocalMux I__11152 (
            .O(N__44838),
            .I(N__44828));
    CEMux I__11151 (
            .O(N__44837),
            .I(N__44825));
    Sp12to4 I__11150 (
            .O(N__44834),
            .I(N__44822));
    IoSpan4Mux I__11149 (
            .O(N__44831),
            .I(N__44819));
    Span4Mux_h I__11148 (
            .O(N__44828),
            .I(N__44816));
    LocalMux I__11147 (
            .O(N__44825),
            .I(N__44813));
    Span12Mux_s8_h I__11146 (
            .O(N__44822),
            .I(N__44810));
    Span4Mux_s0_v I__11145 (
            .O(N__44819),
            .I(N__44807));
    Span4Mux_h I__11144 (
            .O(N__44816),
            .I(N__44804));
    Span4Mux_v I__11143 (
            .O(N__44813),
            .I(N__44801));
    Span12Mux_v I__11142 (
            .O(N__44810),
            .I(N__44798));
    Span4Mux_h I__11141 (
            .O(N__44807),
            .I(N__44795));
    Span4Mux_v I__11140 (
            .O(N__44804),
            .I(N__44792));
    Span4Mux_v I__11139 (
            .O(N__44801),
            .I(N__44789));
    Odrv12 I__11138 (
            .O(N__44798),
            .I(\ALU.a_cnvZ0Z_0 ));
    Odrv4 I__11137 (
            .O(N__44795),
            .I(\ALU.a_cnvZ0Z_0 ));
    Odrv4 I__11136 (
            .O(N__44792),
            .I(\ALU.a_cnvZ0Z_0 ));
    Odrv4 I__11135 (
            .O(N__44789),
            .I(\ALU.a_cnvZ0Z_0 ));
    InMux I__11134 (
            .O(N__44780),
            .I(N__44777));
    LocalMux I__11133 (
            .O(N__44777),
            .I(N__44774));
    Odrv4 I__11132 (
            .O(N__44774),
            .I(\FTDI.TXshiftZ0Z_2 ));
    InMux I__11131 (
            .O(N__44771),
            .I(N__44763));
    InMux I__11130 (
            .O(N__44770),
            .I(N__44763));
    InMux I__11129 (
            .O(N__44769),
            .I(N__44760));
    CascadeMux I__11128 (
            .O(N__44768),
            .I(N__44750));
    LocalMux I__11127 (
            .O(N__44763),
            .I(N__44745));
    LocalMux I__11126 (
            .O(N__44760),
            .I(N__44741));
    InMux I__11125 (
            .O(N__44759),
            .I(N__44726));
    InMux I__11124 (
            .O(N__44758),
            .I(N__44726));
    InMux I__11123 (
            .O(N__44757),
            .I(N__44726));
    InMux I__11122 (
            .O(N__44756),
            .I(N__44726));
    InMux I__11121 (
            .O(N__44755),
            .I(N__44726));
    InMux I__11120 (
            .O(N__44754),
            .I(N__44726));
    InMux I__11119 (
            .O(N__44753),
            .I(N__44726));
    InMux I__11118 (
            .O(N__44750),
            .I(N__44723));
    CascadeMux I__11117 (
            .O(N__44749),
            .I(N__44720));
    CascadeMux I__11116 (
            .O(N__44748),
            .I(N__44714));
    Span4Mux_s2_v I__11115 (
            .O(N__44745),
            .I(N__44711));
    InMux I__11114 (
            .O(N__44744),
            .I(N__44708));
    Span4Mux_h I__11113 (
            .O(N__44741),
            .I(N__44701));
    LocalMux I__11112 (
            .O(N__44726),
            .I(N__44701));
    LocalMux I__11111 (
            .O(N__44723),
            .I(N__44701));
    InMux I__11110 (
            .O(N__44720),
            .I(N__44698));
    InMux I__11109 (
            .O(N__44719),
            .I(N__44693));
    InMux I__11108 (
            .O(N__44718),
            .I(N__44693));
    InMux I__11107 (
            .O(N__44717),
            .I(N__44688));
    InMux I__11106 (
            .O(N__44714),
            .I(N__44688));
    Odrv4 I__11105 (
            .O(N__44711),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__11104 (
            .O(N__44708),
            .I(\FTDI.TXstateZ0Z_3 ));
    Odrv4 I__11103 (
            .O(N__44701),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__11102 (
            .O(N__44698),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__11101 (
            .O(N__44693),
            .I(\FTDI.TXstateZ0Z_3 ));
    LocalMux I__11100 (
            .O(N__44688),
            .I(\FTDI.TXstateZ0Z_3 ));
    InMux I__11099 (
            .O(N__44675),
            .I(N__44672));
    LocalMux I__11098 (
            .O(N__44672),
            .I(N__44669));
    Odrv4 I__11097 (
            .O(N__44669),
            .I(\FTDI.TXshiftZ0Z_1 ));
    CEMux I__11096 (
            .O(N__44666),
            .I(N__44663));
    LocalMux I__11095 (
            .O(N__44663),
            .I(N__44660));
    Span4Mux_h I__11094 (
            .O(N__44660),
            .I(N__44656));
    CEMux I__11093 (
            .O(N__44659),
            .I(N__44653));
    Sp12to4 I__11092 (
            .O(N__44656),
            .I(N__44648));
    LocalMux I__11091 (
            .O(N__44653),
            .I(N__44648));
    Odrv12 I__11090 (
            .O(N__44648),
            .I(\FTDI.un1_TXstate_0_sqmuxa_0_i ));
    InMux I__11089 (
            .O(N__44645),
            .I(N__44642));
    LocalMux I__11088 (
            .O(N__44642),
            .I(N__44638));
    InMux I__11087 (
            .O(N__44641),
            .I(N__44635));
    Span4Mux_v I__11086 (
            .O(N__44638),
            .I(N__44632));
    LocalMux I__11085 (
            .O(N__44635),
            .I(N__44629));
    Span4Mux_h I__11084 (
            .O(N__44632),
            .I(N__44625));
    Span4Mux_h I__11083 (
            .O(N__44629),
            .I(N__44622));
    InMux I__11082 (
            .O(N__44628),
            .I(N__44619));
    Odrv4 I__11081 (
            .O(N__44625),
            .I(a_5));
    Odrv4 I__11080 (
            .O(N__44622),
            .I(a_5));
    LocalMux I__11079 (
            .O(N__44619),
            .I(a_5));
    InMux I__11078 (
            .O(N__44612),
            .I(N__44609));
    LocalMux I__11077 (
            .O(N__44609),
            .I(N__44606));
    Span4Mux_h I__11076 (
            .O(N__44606),
            .I(N__44603));
    Odrv4 I__11075 (
            .O(N__44603),
            .I(TXbufferZ0Z_5));
    InMux I__11074 (
            .O(N__44600),
            .I(N__44597));
    LocalMux I__11073 (
            .O(N__44597),
            .I(N__44593));
    InMux I__11072 (
            .O(N__44596),
            .I(N__44590));
    Span4Mux_v I__11071 (
            .O(N__44593),
            .I(N__44587));
    LocalMux I__11070 (
            .O(N__44590),
            .I(N__44583));
    Span4Mux_h I__11069 (
            .O(N__44587),
            .I(N__44580));
    InMux I__11068 (
            .O(N__44586),
            .I(N__44577));
    Span4Mux_h I__11067 (
            .O(N__44583),
            .I(N__44574));
    Odrv4 I__11066 (
            .O(N__44580),
            .I(a_1));
    LocalMux I__11065 (
            .O(N__44577),
            .I(a_1));
    Odrv4 I__11064 (
            .O(N__44574),
            .I(a_1));
    InMux I__11063 (
            .O(N__44567),
            .I(N__44564));
    LocalMux I__11062 (
            .O(N__44564),
            .I(N__44561));
    Odrv4 I__11061 (
            .O(N__44561),
            .I(TXbufferZ0Z_1));
    CEMux I__11060 (
            .O(N__44558),
            .I(N__44555));
    LocalMux I__11059 (
            .O(N__44555),
            .I(N__44552));
    Span4Mux_v I__11058 (
            .O(N__44552),
            .I(N__44548));
    CEMux I__11057 (
            .O(N__44551),
            .I(N__44545));
    Odrv4 I__11056 (
            .O(N__44548),
            .I(m326dup));
    LocalMux I__11055 (
            .O(N__44545),
            .I(m326dup));
    InMux I__11054 (
            .O(N__44540),
            .I(N__44534));
    InMux I__11053 (
            .O(N__44539),
            .I(N__44531));
    CascadeMux I__11052 (
            .O(N__44538),
            .I(N__44528));
    InMux I__11051 (
            .O(N__44537),
            .I(N__44515));
    LocalMux I__11050 (
            .O(N__44534),
            .I(N__44512));
    LocalMux I__11049 (
            .O(N__44531),
            .I(N__44509));
    InMux I__11048 (
            .O(N__44528),
            .I(N__44506));
    InMux I__11047 (
            .O(N__44527),
            .I(N__44501));
    InMux I__11046 (
            .O(N__44526),
            .I(N__44501));
    CascadeMux I__11045 (
            .O(N__44525),
            .I(N__44496));
    CascadeMux I__11044 (
            .O(N__44524),
            .I(N__44493));
    CascadeMux I__11043 (
            .O(N__44523),
            .I(N__44488));
    CascadeMux I__11042 (
            .O(N__44522),
            .I(N__44484));
    CascadeMux I__11041 (
            .O(N__44521),
            .I(N__44481));
    InMux I__11040 (
            .O(N__44520),
            .I(N__44476));
    InMux I__11039 (
            .O(N__44519),
            .I(N__44471));
    InMux I__11038 (
            .O(N__44518),
            .I(N__44471));
    LocalMux I__11037 (
            .O(N__44515),
            .I(N__44466));
    Span4Mux_v I__11036 (
            .O(N__44512),
            .I(N__44466));
    Span4Mux_v I__11035 (
            .O(N__44509),
            .I(N__44459));
    LocalMux I__11034 (
            .O(N__44506),
            .I(N__44459));
    LocalMux I__11033 (
            .O(N__44501),
            .I(N__44459));
    InMux I__11032 (
            .O(N__44500),
            .I(N__44456));
    InMux I__11031 (
            .O(N__44499),
            .I(N__44453));
    InMux I__11030 (
            .O(N__44496),
            .I(N__44450));
    InMux I__11029 (
            .O(N__44493),
            .I(N__44445));
    CascadeMux I__11028 (
            .O(N__44492),
            .I(N__44439));
    InMux I__11027 (
            .O(N__44491),
            .I(N__44434));
    InMux I__11026 (
            .O(N__44488),
            .I(N__44431));
    InMux I__11025 (
            .O(N__44487),
            .I(N__44426));
    InMux I__11024 (
            .O(N__44484),
            .I(N__44426));
    InMux I__11023 (
            .O(N__44481),
            .I(N__44423));
    InMux I__11022 (
            .O(N__44480),
            .I(N__44417));
    InMux I__11021 (
            .O(N__44479),
            .I(N__44414));
    LocalMux I__11020 (
            .O(N__44476),
            .I(N__44409));
    LocalMux I__11019 (
            .O(N__44471),
            .I(N__44409));
    Span4Mux_v I__11018 (
            .O(N__44466),
            .I(N__44404));
    Span4Mux_v I__11017 (
            .O(N__44459),
            .I(N__44404));
    LocalMux I__11016 (
            .O(N__44456),
            .I(N__44396));
    LocalMux I__11015 (
            .O(N__44453),
            .I(N__44396));
    LocalMux I__11014 (
            .O(N__44450),
            .I(N__44396));
    CascadeMux I__11013 (
            .O(N__44449),
            .I(N__44390));
    InMux I__11012 (
            .O(N__44448),
            .I(N__44387));
    LocalMux I__11011 (
            .O(N__44445),
            .I(N__44384));
    InMux I__11010 (
            .O(N__44444),
            .I(N__44381));
    InMux I__11009 (
            .O(N__44443),
            .I(N__44374));
    InMux I__11008 (
            .O(N__44442),
            .I(N__44374));
    InMux I__11007 (
            .O(N__44439),
            .I(N__44374));
    InMux I__11006 (
            .O(N__44438),
            .I(N__44371));
    InMux I__11005 (
            .O(N__44437),
            .I(N__44368));
    LocalMux I__11004 (
            .O(N__44434),
            .I(N__44363));
    LocalMux I__11003 (
            .O(N__44431),
            .I(N__44363));
    LocalMux I__11002 (
            .O(N__44426),
            .I(N__44358));
    LocalMux I__11001 (
            .O(N__44423),
            .I(N__44358));
    InMux I__11000 (
            .O(N__44422),
            .I(N__44355));
    InMux I__10999 (
            .O(N__44421),
            .I(N__44352));
    InMux I__10998 (
            .O(N__44420),
            .I(N__44349));
    LocalMux I__10997 (
            .O(N__44417),
            .I(N__44346));
    LocalMux I__10996 (
            .O(N__44414),
            .I(N__44341));
    Span4Mux_v I__10995 (
            .O(N__44409),
            .I(N__44341));
    Span4Mux_v I__10994 (
            .O(N__44404),
            .I(N__44338));
    CascadeMux I__10993 (
            .O(N__44403),
            .I(N__44335));
    Span4Mux_h I__10992 (
            .O(N__44396),
            .I(N__44331));
    InMux I__10991 (
            .O(N__44395),
            .I(N__44326));
    InMux I__10990 (
            .O(N__44394),
            .I(N__44326));
    InMux I__10989 (
            .O(N__44393),
            .I(N__44318));
    InMux I__10988 (
            .O(N__44390),
            .I(N__44318));
    LocalMux I__10987 (
            .O(N__44387),
            .I(N__44315));
    Span4Mux_s2_v I__10986 (
            .O(N__44384),
            .I(N__44306));
    LocalMux I__10985 (
            .O(N__44381),
            .I(N__44306));
    LocalMux I__10984 (
            .O(N__44374),
            .I(N__44306));
    LocalMux I__10983 (
            .O(N__44371),
            .I(N__44306));
    LocalMux I__10982 (
            .O(N__44368),
            .I(N__44303));
    Span4Mux_v I__10981 (
            .O(N__44363),
            .I(N__44292));
    Span4Mux_v I__10980 (
            .O(N__44358),
            .I(N__44292));
    LocalMux I__10979 (
            .O(N__44355),
            .I(N__44292));
    LocalMux I__10978 (
            .O(N__44352),
            .I(N__44292));
    LocalMux I__10977 (
            .O(N__44349),
            .I(N__44292));
    Span4Mux_s2_v I__10976 (
            .O(N__44346),
            .I(N__44285));
    Span4Mux_s2_v I__10975 (
            .O(N__44341),
            .I(N__44285));
    Span4Mux_h I__10974 (
            .O(N__44338),
            .I(N__44285));
    InMux I__10973 (
            .O(N__44335),
            .I(N__44280));
    InMux I__10972 (
            .O(N__44334),
            .I(N__44280));
    Sp12to4 I__10971 (
            .O(N__44331),
            .I(N__44275));
    LocalMux I__10970 (
            .O(N__44326),
            .I(N__44275));
    InMux I__10969 (
            .O(N__44325),
            .I(N__44270));
    InMux I__10968 (
            .O(N__44324),
            .I(N__44270));
    InMux I__10967 (
            .O(N__44323),
            .I(N__44267));
    LocalMux I__10966 (
            .O(N__44318),
            .I(N__44260));
    Span4Mux_v I__10965 (
            .O(N__44315),
            .I(N__44260));
    Span4Mux_v I__10964 (
            .O(N__44306),
            .I(N__44260));
    Span12Mux_v I__10963 (
            .O(N__44303),
            .I(N__44249));
    Sp12to4 I__10962 (
            .O(N__44292),
            .I(N__44249));
    Sp12to4 I__10961 (
            .O(N__44285),
            .I(N__44249));
    LocalMux I__10960 (
            .O(N__44280),
            .I(N__44249));
    Span12Mux_s2_v I__10959 (
            .O(N__44275),
            .I(N__44249));
    LocalMux I__10958 (
            .O(N__44270),
            .I(aluParams_3));
    LocalMux I__10957 (
            .O(N__44267),
            .I(aluParams_3));
    Odrv4 I__10956 (
            .O(N__44260),
            .I(aluParams_3));
    Odrv12 I__10955 (
            .O(N__44249),
            .I(aluParams_3));
    InMux I__10954 (
            .O(N__44240),
            .I(N__44237));
    LocalMux I__10953 (
            .O(N__44237),
            .I(N__44234));
    Span4Mux_v I__10952 (
            .O(N__44234),
            .I(N__44231));
    Odrv4 I__10951 (
            .O(N__44231),
            .I(\ALU.N_308 ));
    InMux I__10950 (
            .O(N__44228),
            .I(N__44220));
    InMux I__10949 (
            .O(N__44227),
            .I(N__44215));
    InMux I__10948 (
            .O(N__44226),
            .I(N__44212));
    InMux I__10947 (
            .O(N__44225),
            .I(N__44207));
    InMux I__10946 (
            .O(N__44224),
            .I(N__44207));
    InMux I__10945 (
            .O(N__44223),
            .I(N__44199));
    LocalMux I__10944 (
            .O(N__44220),
            .I(N__44195));
    InMux I__10943 (
            .O(N__44219),
            .I(N__44192));
    CascadeMux I__10942 (
            .O(N__44218),
            .I(N__44189));
    LocalMux I__10941 (
            .O(N__44215),
            .I(N__44182));
    LocalMux I__10940 (
            .O(N__44212),
            .I(N__44182));
    LocalMux I__10939 (
            .O(N__44207),
            .I(N__44179));
    InMux I__10938 (
            .O(N__44206),
            .I(N__44174));
    InMux I__10937 (
            .O(N__44205),
            .I(N__44174));
    InMux I__10936 (
            .O(N__44204),
            .I(N__44169));
    InMux I__10935 (
            .O(N__44203),
            .I(N__44169));
    InMux I__10934 (
            .O(N__44202),
            .I(N__44166));
    LocalMux I__10933 (
            .O(N__44199),
            .I(N__44163));
    InMux I__10932 (
            .O(N__44198),
            .I(N__44160));
    Span4Mux_v I__10931 (
            .O(N__44195),
            .I(N__44156));
    LocalMux I__10930 (
            .O(N__44192),
            .I(N__44153));
    InMux I__10929 (
            .O(N__44189),
            .I(N__44143));
    InMux I__10928 (
            .O(N__44188),
            .I(N__44143));
    InMux I__10927 (
            .O(N__44187),
            .I(N__44140));
    Span4Mux_h I__10926 (
            .O(N__44182),
            .I(N__44134));
    Span4Mux_v I__10925 (
            .O(N__44179),
            .I(N__44134));
    LocalMux I__10924 (
            .O(N__44174),
            .I(N__44122));
    LocalMux I__10923 (
            .O(N__44169),
            .I(N__44122));
    LocalMux I__10922 (
            .O(N__44166),
            .I(N__44122));
    Span4Mux_h I__10921 (
            .O(N__44163),
            .I(N__44122));
    LocalMux I__10920 (
            .O(N__44160),
            .I(N__44122));
    InMux I__10919 (
            .O(N__44159),
            .I(N__44118));
    Span4Mux_h I__10918 (
            .O(N__44156),
            .I(N__44113));
    Span4Mux_v I__10917 (
            .O(N__44153),
            .I(N__44113));
    InMux I__10916 (
            .O(N__44152),
            .I(N__44108));
    InMux I__10915 (
            .O(N__44151),
            .I(N__44108));
    InMux I__10914 (
            .O(N__44150),
            .I(N__44105));
    InMux I__10913 (
            .O(N__44149),
            .I(N__44100));
    InMux I__10912 (
            .O(N__44148),
            .I(N__44100));
    LocalMux I__10911 (
            .O(N__44143),
            .I(N__44097));
    LocalMux I__10910 (
            .O(N__44140),
            .I(N__44094));
    InMux I__10909 (
            .O(N__44139),
            .I(N__44091));
    Span4Mux_h I__10908 (
            .O(N__44134),
            .I(N__44086));
    InMux I__10907 (
            .O(N__44133),
            .I(N__44083));
    Span4Mux_v I__10906 (
            .O(N__44122),
            .I(N__44080));
    InMux I__10905 (
            .O(N__44121),
            .I(N__44077));
    LocalMux I__10904 (
            .O(N__44118),
            .I(N__44074));
    Span4Mux_v I__10903 (
            .O(N__44113),
            .I(N__44071));
    LocalMux I__10902 (
            .O(N__44108),
            .I(N__44068));
    LocalMux I__10901 (
            .O(N__44105),
            .I(N__44061));
    LocalMux I__10900 (
            .O(N__44100),
            .I(N__44061));
    Span4Mux_v I__10899 (
            .O(N__44097),
            .I(N__44061));
    Span4Mux_v I__10898 (
            .O(N__44094),
            .I(N__44055));
    LocalMux I__10897 (
            .O(N__44091),
            .I(N__44055));
    InMux I__10896 (
            .O(N__44090),
            .I(N__44050));
    InMux I__10895 (
            .O(N__44089),
            .I(N__44050));
    Span4Mux_v I__10894 (
            .O(N__44086),
            .I(N__44047));
    LocalMux I__10893 (
            .O(N__44083),
            .I(N__44044));
    Span4Mux_h I__10892 (
            .O(N__44080),
            .I(N__44039));
    LocalMux I__10891 (
            .O(N__44077),
            .I(N__44039));
    Span4Mux_v I__10890 (
            .O(N__44074),
            .I(N__44030));
    Span4Mux_h I__10889 (
            .O(N__44071),
            .I(N__44030));
    Span4Mux_v I__10888 (
            .O(N__44068),
            .I(N__44030));
    Span4Mux_v I__10887 (
            .O(N__44061),
            .I(N__44025));
    InMux I__10886 (
            .O(N__44060),
            .I(N__44022));
    Span4Mux_h I__10885 (
            .O(N__44055),
            .I(N__44013));
    LocalMux I__10884 (
            .O(N__44050),
            .I(N__44013));
    Span4Mux_h I__10883 (
            .O(N__44047),
            .I(N__44013));
    Span4Mux_h I__10882 (
            .O(N__44044),
            .I(N__44013));
    Span4Mux_v I__10881 (
            .O(N__44039),
            .I(N__44010));
    InMux I__10880 (
            .O(N__44038),
            .I(N__44007));
    InMux I__10879 (
            .O(N__44037),
            .I(N__44004));
    Span4Mux_h I__10878 (
            .O(N__44030),
            .I(N__44001));
    InMux I__10877 (
            .O(N__44029),
            .I(N__43998));
    InMux I__10876 (
            .O(N__44028),
            .I(N__43995));
    Sp12to4 I__10875 (
            .O(N__44025),
            .I(N__43992));
    LocalMux I__10874 (
            .O(N__44022),
            .I(N__43987));
    Span4Mux_v I__10873 (
            .O(N__44013),
            .I(N__43987));
    Span4Mux_s0_v I__10872 (
            .O(N__44010),
            .I(N__43984));
    LocalMux I__10871 (
            .O(N__44007),
            .I(aluOperation_2));
    LocalMux I__10870 (
            .O(N__44004),
            .I(aluOperation_2));
    Odrv4 I__10869 (
            .O(N__44001),
            .I(aluOperation_2));
    LocalMux I__10868 (
            .O(N__43998),
            .I(aluOperation_2));
    LocalMux I__10867 (
            .O(N__43995),
            .I(aluOperation_2));
    Odrv12 I__10866 (
            .O(N__43992),
            .I(aluOperation_2));
    Odrv4 I__10865 (
            .O(N__43987),
            .I(aluOperation_2));
    Odrv4 I__10864 (
            .O(N__43984),
            .I(aluOperation_2));
    CascadeMux I__10863 (
            .O(N__43967),
            .I(N__43964));
    InMux I__10862 (
            .O(N__43964),
            .I(N__43959));
    CascadeMux I__10861 (
            .O(N__43963),
            .I(N__43956));
    CascadeMux I__10860 (
            .O(N__43962),
            .I(N__43953));
    LocalMux I__10859 (
            .O(N__43959),
            .I(N__43949));
    InMux I__10858 (
            .O(N__43956),
            .I(N__43946));
    InMux I__10857 (
            .O(N__43953),
            .I(N__43943));
    CascadeMux I__10856 (
            .O(N__43952),
            .I(N__43940));
    Span4Mux_h I__10855 (
            .O(N__43949),
            .I(N__43934));
    LocalMux I__10854 (
            .O(N__43946),
            .I(N__43930));
    LocalMux I__10853 (
            .O(N__43943),
            .I(N__43926));
    InMux I__10852 (
            .O(N__43940),
            .I(N__43923));
    CascadeMux I__10851 (
            .O(N__43939),
            .I(N__43920));
    CascadeMux I__10850 (
            .O(N__43938),
            .I(N__43916));
    InMux I__10849 (
            .O(N__43937),
            .I(N__43913));
    Span4Mux_h I__10848 (
            .O(N__43934),
            .I(N__43910));
    InMux I__10847 (
            .O(N__43933),
            .I(N__43907));
    Span4Mux_v I__10846 (
            .O(N__43930),
            .I(N__43904));
    CascadeMux I__10845 (
            .O(N__43929),
            .I(N__43901));
    Span4Mux_h I__10844 (
            .O(N__43926),
            .I(N__43894));
    LocalMux I__10843 (
            .O(N__43923),
            .I(N__43894));
    InMux I__10842 (
            .O(N__43920),
            .I(N__43891));
    CascadeMux I__10841 (
            .O(N__43919),
            .I(N__43888));
    InMux I__10840 (
            .O(N__43916),
            .I(N__43885));
    LocalMux I__10839 (
            .O(N__43913),
            .I(N__43882));
    Span4Mux_v I__10838 (
            .O(N__43910),
            .I(N__43876));
    LocalMux I__10837 (
            .O(N__43907),
            .I(N__43876));
    Span4Mux_v I__10836 (
            .O(N__43904),
            .I(N__43873));
    InMux I__10835 (
            .O(N__43901),
            .I(N__43870));
    InMux I__10834 (
            .O(N__43900),
            .I(N__43865));
    InMux I__10833 (
            .O(N__43899),
            .I(N__43865));
    Span4Mux_h I__10832 (
            .O(N__43894),
            .I(N__43862));
    LocalMux I__10831 (
            .O(N__43891),
            .I(N__43856));
    InMux I__10830 (
            .O(N__43888),
            .I(N__43853));
    LocalMux I__10829 (
            .O(N__43885),
            .I(N__43850));
    Span4Mux_v I__10828 (
            .O(N__43882),
            .I(N__43847));
    CascadeMux I__10827 (
            .O(N__43881),
            .I(N__43844));
    Span4Mux_v I__10826 (
            .O(N__43876),
            .I(N__43841));
    Span4Mux_v I__10825 (
            .O(N__43873),
            .I(N__43838));
    LocalMux I__10824 (
            .O(N__43870),
            .I(N__43833));
    LocalMux I__10823 (
            .O(N__43865),
            .I(N__43833));
    Span4Mux_h I__10822 (
            .O(N__43862),
            .I(N__43830));
    InMux I__10821 (
            .O(N__43861),
            .I(N__43825));
    InMux I__10820 (
            .O(N__43860),
            .I(N__43825));
    InMux I__10819 (
            .O(N__43859),
            .I(N__43822));
    Span4Mux_v I__10818 (
            .O(N__43856),
            .I(N__43819));
    LocalMux I__10817 (
            .O(N__43853),
            .I(N__43816));
    Span4Mux_v I__10816 (
            .O(N__43850),
            .I(N__43811));
    Span4Mux_h I__10815 (
            .O(N__43847),
            .I(N__43811));
    InMux I__10814 (
            .O(N__43844),
            .I(N__43808));
    Span4Mux_v I__10813 (
            .O(N__43841),
            .I(N__43805));
    Span4Mux_h I__10812 (
            .O(N__43838),
            .I(N__43800));
    Span4Mux_v I__10811 (
            .O(N__43833),
            .I(N__43800));
    Span4Mux_v I__10810 (
            .O(N__43830),
            .I(N__43795));
    LocalMux I__10809 (
            .O(N__43825),
            .I(N__43795));
    LocalMux I__10808 (
            .O(N__43822),
            .I(N__43792));
    Span4Mux_h I__10807 (
            .O(N__43819),
            .I(N__43781));
    Span4Mux_v I__10806 (
            .O(N__43816),
            .I(N__43781));
    Span4Mux_v I__10805 (
            .O(N__43811),
            .I(N__43781));
    LocalMux I__10804 (
            .O(N__43808),
            .I(N__43781));
    Span4Mux_s1_v I__10803 (
            .O(N__43805),
            .I(N__43781));
    Span4Mux_h I__10802 (
            .O(N__43800),
            .I(N__43776));
    Span4Mux_v I__10801 (
            .O(N__43795),
            .I(N__43776));
    Odrv4 I__10800 (
            .O(N__43792),
            .I(\ALU.log_0_sqmuxa ));
    Odrv4 I__10799 (
            .O(N__43781),
            .I(\ALU.log_0_sqmuxa ));
    Odrv4 I__10798 (
            .O(N__43776),
            .I(\ALU.log_0_sqmuxa ));
    CascadeMux I__10797 (
            .O(N__43769),
            .I(N__43764));
    InMux I__10796 (
            .O(N__43768),
            .I(N__43758));
    InMux I__10795 (
            .O(N__43767),
            .I(N__43755));
    InMux I__10794 (
            .O(N__43764),
            .I(N__43751));
    InMux I__10793 (
            .O(N__43763),
            .I(N__43748));
    InMux I__10792 (
            .O(N__43762),
            .I(N__43744));
    InMux I__10791 (
            .O(N__43761),
            .I(N__43741));
    LocalMux I__10790 (
            .O(N__43758),
            .I(N__43736));
    LocalMux I__10789 (
            .O(N__43755),
            .I(N__43736));
    InMux I__10788 (
            .O(N__43754),
            .I(N__43733));
    LocalMux I__10787 (
            .O(N__43751),
            .I(N__43730));
    LocalMux I__10786 (
            .O(N__43748),
            .I(N__43723));
    CascadeMux I__10785 (
            .O(N__43747),
            .I(N__43720));
    LocalMux I__10784 (
            .O(N__43744),
            .I(N__43716));
    LocalMux I__10783 (
            .O(N__43741),
            .I(N__43708));
    Span4Mux_v I__10782 (
            .O(N__43736),
            .I(N__43708));
    LocalMux I__10781 (
            .O(N__43733),
            .I(N__43704));
    Span4Mux_v I__10780 (
            .O(N__43730),
            .I(N__43701));
    InMux I__10779 (
            .O(N__43729),
            .I(N__43698));
    InMux I__10778 (
            .O(N__43728),
            .I(N__43694));
    CascadeMux I__10777 (
            .O(N__43727),
            .I(N__43691));
    InMux I__10776 (
            .O(N__43726),
            .I(N__43685));
    Span4Mux_v I__10775 (
            .O(N__43723),
            .I(N__43680));
    InMux I__10774 (
            .O(N__43720),
            .I(N__43677));
    CascadeMux I__10773 (
            .O(N__43719),
            .I(N__43670));
    Span4Mux_v I__10772 (
            .O(N__43716),
            .I(N__43661));
    InMux I__10771 (
            .O(N__43715),
            .I(N__43654));
    InMux I__10770 (
            .O(N__43714),
            .I(N__43654));
    InMux I__10769 (
            .O(N__43713),
            .I(N__43654));
    Span4Mux_v I__10768 (
            .O(N__43708),
            .I(N__43650));
    InMux I__10767 (
            .O(N__43707),
            .I(N__43647));
    Span4Mux_h I__10766 (
            .O(N__43704),
            .I(N__43642));
    Span4Mux_v I__10765 (
            .O(N__43701),
            .I(N__43642));
    LocalMux I__10764 (
            .O(N__43698),
            .I(N__43639));
    InMux I__10763 (
            .O(N__43697),
            .I(N__43635));
    LocalMux I__10762 (
            .O(N__43694),
            .I(N__43632));
    InMux I__10761 (
            .O(N__43691),
            .I(N__43629));
    InMux I__10760 (
            .O(N__43690),
            .I(N__43626));
    InMux I__10759 (
            .O(N__43689),
            .I(N__43623));
    InMux I__10758 (
            .O(N__43688),
            .I(N__43617));
    LocalMux I__10757 (
            .O(N__43685),
            .I(N__43614));
    InMux I__10756 (
            .O(N__43684),
            .I(N__43609));
    InMux I__10755 (
            .O(N__43683),
            .I(N__43609));
    Span4Mux_v I__10754 (
            .O(N__43680),
            .I(N__43604));
    LocalMux I__10753 (
            .O(N__43677),
            .I(N__43604));
    InMux I__10752 (
            .O(N__43676),
            .I(N__43601));
    InMux I__10751 (
            .O(N__43675),
            .I(N__43598));
    InMux I__10750 (
            .O(N__43674),
            .I(N__43595));
    InMux I__10749 (
            .O(N__43673),
            .I(N__43588));
    InMux I__10748 (
            .O(N__43670),
            .I(N__43588));
    InMux I__10747 (
            .O(N__43669),
            .I(N__43588));
    InMux I__10746 (
            .O(N__43668),
            .I(N__43579));
    InMux I__10745 (
            .O(N__43667),
            .I(N__43576));
    InMux I__10744 (
            .O(N__43666),
            .I(N__43573));
    InMux I__10743 (
            .O(N__43665),
            .I(N__43568));
    InMux I__10742 (
            .O(N__43664),
            .I(N__43568));
    Span4Mux_v I__10741 (
            .O(N__43661),
            .I(N__43565));
    LocalMux I__10740 (
            .O(N__43654),
            .I(N__43562));
    InMux I__10739 (
            .O(N__43653),
            .I(N__43559));
    Span4Mux_h I__10738 (
            .O(N__43650),
            .I(N__43552));
    LocalMux I__10737 (
            .O(N__43647),
            .I(N__43552));
    Span4Mux_v I__10736 (
            .O(N__43642),
            .I(N__43552));
    Sp12to4 I__10735 (
            .O(N__43639),
            .I(N__43549));
    CascadeMux I__10734 (
            .O(N__43638),
            .I(N__43546));
    LocalMux I__10733 (
            .O(N__43635),
            .I(N__43542));
    Span4Mux_v I__10732 (
            .O(N__43632),
            .I(N__43533));
    LocalMux I__10731 (
            .O(N__43629),
            .I(N__43533));
    LocalMux I__10730 (
            .O(N__43626),
            .I(N__43533));
    LocalMux I__10729 (
            .O(N__43623),
            .I(N__43533));
    InMux I__10728 (
            .O(N__43622),
            .I(N__43528));
    InMux I__10727 (
            .O(N__43621),
            .I(N__43528));
    InMux I__10726 (
            .O(N__43620),
            .I(N__43525));
    LocalMux I__10725 (
            .O(N__43617),
            .I(N__43522));
    Span4Mux_h I__10724 (
            .O(N__43614),
            .I(N__43517));
    LocalMux I__10723 (
            .O(N__43609),
            .I(N__43517));
    Span4Mux_h I__10722 (
            .O(N__43604),
            .I(N__43512));
    LocalMux I__10721 (
            .O(N__43601),
            .I(N__43512));
    LocalMux I__10720 (
            .O(N__43598),
            .I(N__43507));
    LocalMux I__10719 (
            .O(N__43595),
            .I(N__43502));
    LocalMux I__10718 (
            .O(N__43588),
            .I(N__43502));
    InMux I__10717 (
            .O(N__43587),
            .I(N__43495));
    InMux I__10716 (
            .O(N__43586),
            .I(N__43495));
    InMux I__10715 (
            .O(N__43585),
            .I(N__43495));
    InMux I__10714 (
            .O(N__43584),
            .I(N__43492));
    InMux I__10713 (
            .O(N__43583),
            .I(N__43486));
    InMux I__10712 (
            .O(N__43582),
            .I(N__43486));
    LocalMux I__10711 (
            .O(N__43579),
            .I(N__43471));
    LocalMux I__10710 (
            .O(N__43576),
            .I(N__43471));
    LocalMux I__10709 (
            .O(N__43573),
            .I(N__43471));
    LocalMux I__10708 (
            .O(N__43568),
            .I(N__43471));
    Span4Mux_h I__10707 (
            .O(N__43565),
            .I(N__43471));
    Span4Mux_h I__10706 (
            .O(N__43562),
            .I(N__43471));
    LocalMux I__10705 (
            .O(N__43559),
            .I(N__43471));
    Span4Mux_v I__10704 (
            .O(N__43552),
            .I(N__43468));
    Span12Mux_v I__10703 (
            .O(N__43549),
            .I(N__43465));
    InMux I__10702 (
            .O(N__43546),
            .I(N__43460));
    InMux I__10701 (
            .O(N__43545),
            .I(N__43460));
    Span4Mux_h I__10700 (
            .O(N__43542),
            .I(N__43455));
    Span4Mux_h I__10699 (
            .O(N__43533),
            .I(N__43455));
    LocalMux I__10698 (
            .O(N__43528),
            .I(N__43448));
    LocalMux I__10697 (
            .O(N__43525),
            .I(N__43448));
    Span4Mux_h I__10696 (
            .O(N__43522),
            .I(N__43448));
    Span4Mux_v I__10695 (
            .O(N__43517),
            .I(N__43443));
    Span4Mux_h I__10694 (
            .O(N__43512),
            .I(N__43443));
    InMux I__10693 (
            .O(N__43511),
            .I(N__43438));
    InMux I__10692 (
            .O(N__43510),
            .I(N__43438));
    Span12Mux_h I__10691 (
            .O(N__43507),
            .I(N__43429));
    Sp12to4 I__10690 (
            .O(N__43502),
            .I(N__43429));
    LocalMux I__10689 (
            .O(N__43495),
            .I(N__43429));
    LocalMux I__10688 (
            .O(N__43492),
            .I(N__43429));
    InMux I__10687 (
            .O(N__43491),
            .I(N__43426));
    LocalMux I__10686 (
            .O(N__43486),
            .I(N__43419));
    Span4Mux_v I__10685 (
            .O(N__43471),
            .I(N__43419));
    Span4Mux_s1_v I__10684 (
            .O(N__43468),
            .I(N__43419));
    Odrv12 I__10683 (
            .O(N__43465),
            .I(aluParams_0));
    LocalMux I__10682 (
            .O(N__43460),
            .I(aluParams_0));
    Odrv4 I__10681 (
            .O(N__43455),
            .I(aluParams_0));
    Odrv4 I__10680 (
            .O(N__43448),
            .I(aluParams_0));
    Odrv4 I__10679 (
            .O(N__43443),
            .I(aluParams_0));
    LocalMux I__10678 (
            .O(N__43438),
            .I(aluParams_0));
    Odrv12 I__10677 (
            .O(N__43429),
            .I(aluParams_0));
    LocalMux I__10676 (
            .O(N__43426),
            .I(aluParams_0));
    Odrv4 I__10675 (
            .O(N__43419),
            .I(aluParams_0));
    InMux I__10674 (
            .O(N__43400),
            .I(N__43397));
    LocalMux I__10673 (
            .O(N__43397),
            .I(N__43393));
    InMux I__10672 (
            .O(N__43396),
            .I(N__43390));
    Span4Mux_h I__10671 (
            .O(N__43393),
            .I(N__43387));
    LocalMux I__10670 (
            .O(N__43390),
            .I(N__43384));
    Span4Mux_h I__10669 (
            .O(N__43387),
            .I(N__43381));
    Span4Mux_h I__10668 (
            .O(N__43384),
            .I(N__43378));
    Odrv4 I__10667 (
            .O(N__43381),
            .I(\ALU.dZ0Z_5 ));
    Odrv4 I__10666 (
            .O(N__43378),
            .I(\ALU.dZ0Z_5 ));
    InMux I__10665 (
            .O(N__43373),
            .I(N__43369));
    InMux I__10664 (
            .O(N__43372),
            .I(N__43366));
    LocalMux I__10663 (
            .O(N__43369),
            .I(N__43363));
    LocalMux I__10662 (
            .O(N__43366),
            .I(N__43360));
    Span4Mux_h I__10661 (
            .O(N__43363),
            .I(N__43357));
    Span4Mux_h I__10660 (
            .O(N__43360),
            .I(N__43354));
    Span4Mux_h I__10659 (
            .O(N__43357),
            .I(N__43351));
    Odrv4 I__10658 (
            .O(N__43354),
            .I(\ALU.dZ0Z_6 ));
    Odrv4 I__10657 (
            .O(N__43351),
            .I(\ALU.dZ0Z_6 ));
    CEMux I__10656 (
            .O(N__43346),
            .I(N__43341));
    CEMux I__10655 (
            .O(N__43345),
            .I(N__43337));
    CEMux I__10654 (
            .O(N__43344),
            .I(N__43334));
    LocalMux I__10653 (
            .O(N__43341),
            .I(N__43331));
    CEMux I__10652 (
            .O(N__43340),
            .I(N__43328));
    LocalMux I__10651 (
            .O(N__43337),
            .I(N__43325));
    LocalMux I__10650 (
            .O(N__43334),
            .I(N__43321));
    Span4Mux_h I__10649 (
            .O(N__43331),
            .I(N__43318));
    LocalMux I__10648 (
            .O(N__43328),
            .I(N__43315));
    Span4Mux_v I__10647 (
            .O(N__43325),
            .I(N__43312));
    CEMux I__10646 (
            .O(N__43324),
            .I(N__43309));
    Sp12to4 I__10645 (
            .O(N__43321),
            .I(N__43306));
    Span4Mux_v I__10644 (
            .O(N__43318),
            .I(N__43301));
    Span4Mux_h I__10643 (
            .O(N__43315),
            .I(N__43301));
    Span4Mux_h I__10642 (
            .O(N__43312),
            .I(N__43298));
    LocalMux I__10641 (
            .O(N__43309),
            .I(N__43295));
    Span12Mux_h I__10640 (
            .O(N__43306),
            .I(N__43292));
    Sp12to4 I__10639 (
            .O(N__43301),
            .I(N__43287));
    Sp12to4 I__10638 (
            .O(N__43298),
            .I(N__43287));
    Span4Mux_s1_v I__10637 (
            .O(N__43295),
            .I(N__43284));
    Span12Mux_v I__10636 (
            .O(N__43292),
            .I(N__43281));
    Span12Mux_v I__10635 (
            .O(N__43287),
            .I(N__43278));
    Span4Mux_h I__10634 (
            .O(N__43284),
            .I(N__43275));
    Odrv12 I__10633 (
            .O(N__43281),
            .I(\ALU.d_cnvZ0Z_0 ));
    Odrv12 I__10632 (
            .O(N__43278),
            .I(\ALU.d_cnvZ0Z_0 ));
    Odrv4 I__10631 (
            .O(N__43275),
            .I(\ALU.d_cnvZ0Z_0 ));
    CascadeMux I__10630 (
            .O(N__43268),
            .I(N__43265));
    InMux I__10629 (
            .O(N__43265),
            .I(N__43262));
    LocalMux I__10628 (
            .O(N__43262),
            .I(N__43258));
    InMux I__10627 (
            .O(N__43261),
            .I(N__43255));
    Span4Mux_v I__10626 (
            .O(N__43258),
            .I(N__43252));
    LocalMux I__10625 (
            .O(N__43255),
            .I(\ALU.fZ0Z_3 ));
    Odrv4 I__10624 (
            .O(N__43252),
            .I(\ALU.fZ0Z_3 ));
    InMux I__10623 (
            .O(N__43247),
            .I(N__43244));
    LocalMux I__10622 (
            .O(N__43244),
            .I(N__43241));
    Span4Mux_v I__10621 (
            .O(N__43241),
            .I(N__43238));
    Span4Mux_h I__10620 (
            .O(N__43238),
            .I(N__43235));
    Odrv4 I__10619 (
            .O(N__43235),
            .I(\ALU.f_RNIHUEJZ0Z_3 ));
    InMux I__10618 (
            .O(N__43232),
            .I(N__43228));
    InMux I__10617 (
            .O(N__43231),
            .I(N__43225));
    LocalMux I__10616 (
            .O(N__43228),
            .I(N__43222));
    LocalMux I__10615 (
            .O(N__43225),
            .I(N__43219));
    Span12Mux_v I__10614 (
            .O(N__43222),
            .I(N__43216));
    Odrv12 I__10613 (
            .O(N__43219),
            .I(\ALU.rshift_1_12 ));
    Odrv12 I__10612 (
            .O(N__43216),
            .I(\ALU.rshift_1_12 ));
    InMux I__10611 (
            .O(N__43211),
            .I(N__43208));
    LocalMux I__10610 (
            .O(N__43208),
            .I(N__43205));
    Span4Mux_v I__10609 (
            .O(N__43205),
            .I(N__43202));
    Sp12to4 I__10608 (
            .O(N__43202),
            .I(N__43199));
    Span12Mux_h I__10607 (
            .O(N__43199),
            .I(N__43196));
    Odrv12 I__10606 (
            .O(N__43196),
            .I(\ALU.N_532 ));
    InMux I__10605 (
            .O(N__43193),
            .I(N__43190));
    LocalMux I__10604 (
            .O(N__43190),
            .I(N__43186));
    CascadeMux I__10603 (
            .O(N__43189),
            .I(N__43181));
    Span4Mux_v I__10602 (
            .O(N__43186),
            .I(N__43176));
    InMux I__10601 (
            .O(N__43185),
            .I(N__43173));
    CascadeMux I__10600 (
            .O(N__43184),
            .I(N__43169));
    InMux I__10599 (
            .O(N__43181),
            .I(N__43166));
    CascadeMux I__10598 (
            .O(N__43180),
            .I(N__43162));
    InMux I__10597 (
            .O(N__43179),
            .I(N__43159));
    Span4Mux_v I__10596 (
            .O(N__43176),
            .I(N__43156));
    LocalMux I__10595 (
            .O(N__43173),
            .I(N__43153));
    InMux I__10594 (
            .O(N__43172),
            .I(N__43144));
    InMux I__10593 (
            .O(N__43169),
            .I(N__43144));
    LocalMux I__10592 (
            .O(N__43166),
            .I(N__43141));
    InMux I__10591 (
            .O(N__43165),
            .I(N__43136));
    InMux I__10590 (
            .O(N__43162),
            .I(N__43133));
    LocalMux I__10589 (
            .O(N__43159),
            .I(N__43130));
    Span4Mux_v I__10588 (
            .O(N__43156),
            .I(N__43125));
    Span4Mux_v I__10587 (
            .O(N__43153),
            .I(N__43125));
    InMux I__10586 (
            .O(N__43152),
            .I(N__43120));
    InMux I__10585 (
            .O(N__43151),
            .I(N__43120));
    InMux I__10584 (
            .O(N__43150),
            .I(N__43117));
    InMux I__10583 (
            .O(N__43149),
            .I(N__43114));
    LocalMux I__10582 (
            .O(N__43144),
            .I(N__43111));
    Span4Mux_v I__10581 (
            .O(N__43141),
            .I(N__43106));
    InMux I__10580 (
            .O(N__43140),
            .I(N__43101));
    InMux I__10579 (
            .O(N__43139),
            .I(N__43101));
    LocalMux I__10578 (
            .O(N__43136),
            .I(N__43098));
    LocalMux I__10577 (
            .O(N__43133),
            .I(N__43094));
    Span4Mux_v I__10576 (
            .O(N__43130),
            .I(N__43091));
    Span4Mux_v I__10575 (
            .O(N__43125),
            .I(N__43087));
    LocalMux I__10574 (
            .O(N__43120),
            .I(N__43082));
    LocalMux I__10573 (
            .O(N__43117),
            .I(N__43082));
    LocalMux I__10572 (
            .O(N__43114),
            .I(N__43077));
    Span4Mux_h I__10571 (
            .O(N__43111),
            .I(N__43077));
    InMux I__10570 (
            .O(N__43110),
            .I(N__43072));
    InMux I__10569 (
            .O(N__43109),
            .I(N__43072));
    Span4Mux_h I__10568 (
            .O(N__43106),
            .I(N__43067));
    LocalMux I__10567 (
            .O(N__43101),
            .I(N__43067));
    Span4Mux_v I__10566 (
            .O(N__43098),
            .I(N__43064));
    InMux I__10565 (
            .O(N__43097),
            .I(N__43061));
    Span4Mux_s3_h I__10564 (
            .O(N__43094),
            .I(N__43056));
    Span4Mux_h I__10563 (
            .O(N__43091),
            .I(N__43056));
    InMux I__10562 (
            .O(N__43090),
            .I(N__43053));
    Span4Mux_h I__10561 (
            .O(N__43087),
            .I(N__43048));
    Span4Mux_v I__10560 (
            .O(N__43082),
            .I(N__43048));
    Span4Mux_h I__10559 (
            .O(N__43077),
            .I(N__43043));
    LocalMux I__10558 (
            .O(N__43072),
            .I(N__43043));
    Span4Mux_v I__10557 (
            .O(N__43067),
            .I(N__43038));
    Span4Mux_h I__10556 (
            .O(N__43064),
            .I(N__43038));
    LocalMux I__10555 (
            .O(N__43061),
            .I(aluOperation_4));
    Odrv4 I__10554 (
            .O(N__43056),
            .I(aluOperation_4));
    LocalMux I__10553 (
            .O(N__43053),
            .I(aluOperation_4));
    Odrv4 I__10552 (
            .O(N__43048),
            .I(aluOperation_4));
    Odrv4 I__10551 (
            .O(N__43043),
            .I(aluOperation_4));
    Odrv4 I__10550 (
            .O(N__43038),
            .I(aluOperation_4));
    CascadeMux I__10549 (
            .O(N__43025),
            .I(\ALU.rshift_4_cascade_ ));
    InMux I__10548 (
            .O(N__43022),
            .I(N__43019));
    LocalMux I__10547 (
            .O(N__43019),
            .I(N__43016));
    Span4Mux_v I__10546 (
            .O(N__43016),
            .I(N__43013));
    Span4Mux_v I__10545 (
            .O(N__43013),
            .I(N__43010));
    Span4Mux_h I__10544 (
            .O(N__43010),
            .I(N__43007));
    Span4Mux_h I__10543 (
            .O(N__43007),
            .I(N__43004));
    Odrv4 I__10542 (
            .O(N__43004),
            .I(\ALU.N_289_0 ));
    CascadeMux I__10541 (
            .O(N__43001),
            .I(\ALU.a_15_m3_4_cascade_ ));
    InMux I__10540 (
            .O(N__42998),
            .I(N__42987));
    CascadeMux I__10539 (
            .O(N__42997),
            .I(N__42984));
    InMux I__10538 (
            .O(N__42996),
            .I(N__42981));
    InMux I__10537 (
            .O(N__42995),
            .I(N__42977));
    InMux I__10536 (
            .O(N__42994),
            .I(N__42974));
    InMux I__10535 (
            .O(N__42993),
            .I(N__42966));
    InMux I__10534 (
            .O(N__42992),
            .I(N__42963));
    InMux I__10533 (
            .O(N__42991),
            .I(N__42960));
    CascadeMux I__10532 (
            .O(N__42990),
            .I(N__42954));
    LocalMux I__10531 (
            .O(N__42987),
            .I(N__42951));
    InMux I__10530 (
            .O(N__42984),
            .I(N__42948));
    LocalMux I__10529 (
            .O(N__42981),
            .I(N__42942));
    InMux I__10528 (
            .O(N__42980),
            .I(N__42939));
    LocalMux I__10527 (
            .O(N__42977),
            .I(N__42934));
    LocalMux I__10526 (
            .O(N__42974),
            .I(N__42934));
    InMux I__10525 (
            .O(N__42973),
            .I(N__42928));
    InMux I__10524 (
            .O(N__42972),
            .I(N__42928));
    CascadeMux I__10523 (
            .O(N__42971),
            .I(N__42923));
    CascadeMux I__10522 (
            .O(N__42970),
            .I(N__42920));
    CascadeMux I__10521 (
            .O(N__42969),
            .I(N__42917));
    LocalMux I__10520 (
            .O(N__42966),
            .I(N__42913));
    LocalMux I__10519 (
            .O(N__42963),
            .I(N__42910));
    LocalMux I__10518 (
            .O(N__42960),
            .I(N__42907));
    InMux I__10517 (
            .O(N__42959),
            .I(N__42900));
    InMux I__10516 (
            .O(N__42958),
            .I(N__42897));
    InMux I__10515 (
            .O(N__42957),
            .I(N__42892));
    InMux I__10514 (
            .O(N__42954),
            .I(N__42892));
    Span4Mux_s3_v I__10513 (
            .O(N__42951),
            .I(N__42886));
    LocalMux I__10512 (
            .O(N__42948),
            .I(N__42886));
    InMux I__10511 (
            .O(N__42947),
            .I(N__42879));
    InMux I__10510 (
            .O(N__42946),
            .I(N__42879));
    InMux I__10509 (
            .O(N__42945),
            .I(N__42879));
    Span4Mux_s3_v I__10508 (
            .O(N__42942),
            .I(N__42874));
    LocalMux I__10507 (
            .O(N__42939),
            .I(N__42874));
    Span4Mux_h I__10506 (
            .O(N__42934),
            .I(N__42871));
    InMux I__10505 (
            .O(N__42933),
            .I(N__42868));
    LocalMux I__10504 (
            .O(N__42928),
            .I(N__42865));
    InMux I__10503 (
            .O(N__42927),
            .I(N__42862));
    InMux I__10502 (
            .O(N__42926),
            .I(N__42859));
    InMux I__10501 (
            .O(N__42923),
            .I(N__42856));
    InMux I__10500 (
            .O(N__42920),
            .I(N__42849));
    InMux I__10499 (
            .O(N__42917),
            .I(N__42849));
    InMux I__10498 (
            .O(N__42916),
            .I(N__42849));
    Span4Mux_v I__10497 (
            .O(N__42913),
            .I(N__42844));
    Span4Mux_v I__10496 (
            .O(N__42910),
            .I(N__42844));
    Span4Mux_v I__10495 (
            .O(N__42907),
            .I(N__42841));
    InMux I__10494 (
            .O(N__42906),
            .I(N__42838));
    InMux I__10493 (
            .O(N__42905),
            .I(N__42835));
    InMux I__10492 (
            .O(N__42904),
            .I(N__42830));
    InMux I__10491 (
            .O(N__42903),
            .I(N__42830));
    LocalMux I__10490 (
            .O(N__42900),
            .I(N__42827));
    LocalMux I__10489 (
            .O(N__42897),
            .I(N__42824));
    LocalMux I__10488 (
            .O(N__42892),
            .I(N__42818));
    InMux I__10487 (
            .O(N__42891),
            .I(N__42815));
    Span4Mux_h I__10486 (
            .O(N__42886),
            .I(N__42810));
    LocalMux I__10485 (
            .O(N__42879),
            .I(N__42810));
    Span4Mux_v I__10484 (
            .O(N__42874),
            .I(N__42807));
    Span4Mux_v I__10483 (
            .O(N__42871),
            .I(N__42800));
    LocalMux I__10482 (
            .O(N__42868),
            .I(N__42800));
    Span4Mux_s2_h I__10481 (
            .O(N__42865),
            .I(N__42800));
    LocalMux I__10480 (
            .O(N__42862),
            .I(N__42797));
    LocalMux I__10479 (
            .O(N__42859),
            .I(N__42790));
    LocalMux I__10478 (
            .O(N__42856),
            .I(N__42790));
    LocalMux I__10477 (
            .O(N__42849),
            .I(N__42790));
    Span4Mux_h I__10476 (
            .O(N__42844),
            .I(N__42782));
    Span4Mux_v I__10475 (
            .O(N__42841),
            .I(N__42782));
    LocalMux I__10474 (
            .O(N__42838),
            .I(N__42777));
    LocalMux I__10473 (
            .O(N__42835),
            .I(N__42777));
    LocalMux I__10472 (
            .O(N__42830),
            .I(N__42774));
    Span4Mux_v I__10471 (
            .O(N__42827),
            .I(N__42769));
    Span4Mux_s1_h I__10470 (
            .O(N__42824),
            .I(N__42769));
    InMux I__10469 (
            .O(N__42823),
            .I(N__42764));
    InMux I__10468 (
            .O(N__42822),
            .I(N__42764));
    InMux I__10467 (
            .O(N__42821),
            .I(N__42761));
    Span4Mux_h I__10466 (
            .O(N__42818),
            .I(N__42758));
    LocalMux I__10465 (
            .O(N__42815),
            .I(N__42753));
    Span4Mux_v I__10464 (
            .O(N__42810),
            .I(N__42753));
    Span4Mux_v I__10463 (
            .O(N__42807),
            .I(N__42748));
    Span4Mux_v I__10462 (
            .O(N__42800),
            .I(N__42748));
    Span4Mux_h I__10461 (
            .O(N__42797),
            .I(N__42743));
    Span4Mux_v I__10460 (
            .O(N__42790),
            .I(N__42743));
    InMux I__10459 (
            .O(N__42789),
            .I(N__42738));
    InMux I__10458 (
            .O(N__42788),
            .I(N__42738));
    InMux I__10457 (
            .O(N__42787),
            .I(N__42735));
    Span4Mux_h I__10456 (
            .O(N__42782),
            .I(N__42724));
    Span4Mux_h I__10455 (
            .O(N__42777),
            .I(N__42724));
    Span4Mux_v I__10454 (
            .O(N__42774),
            .I(N__42724));
    Span4Mux_h I__10453 (
            .O(N__42769),
            .I(N__42724));
    LocalMux I__10452 (
            .O(N__42764),
            .I(N__42724));
    LocalMux I__10451 (
            .O(N__42761),
            .I(\ALU.aluOut_4 ));
    Odrv4 I__10450 (
            .O(N__42758),
            .I(\ALU.aluOut_4 ));
    Odrv4 I__10449 (
            .O(N__42753),
            .I(\ALU.aluOut_4 ));
    Odrv4 I__10448 (
            .O(N__42748),
            .I(\ALU.aluOut_4 ));
    Odrv4 I__10447 (
            .O(N__42743),
            .I(\ALU.aluOut_4 ));
    LocalMux I__10446 (
            .O(N__42738),
            .I(\ALU.aluOut_4 ));
    LocalMux I__10445 (
            .O(N__42735),
            .I(\ALU.aluOut_4 ));
    Odrv4 I__10444 (
            .O(N__42724),
            .I(\ALU.aluOut_4 ));
    CascadeMux I__10443 (
            .O(N__42707),
            .I(N__42704));
    InMux I__10442 (
            .O(N__42704),
            .I(N__42701));
    LocalMux I__10441 (
            .O(N__42701),
            .I(\ALU.a_15_m2_ns_1Z0Z_4 ));
    CascadeMux I__10440 (
            .O(N__42698),
            .I(N__42693));
    InMux I__10439 (
            .O(N__42697),
            .I(N__42684));
    InMux I__10438 (
            .O(N__42696),
            .I(N__42680));
    InMux I__10437 (
            .O(N__42693),
            .I(N__42677));
    InMux I__10436 (
            .O(N__42692),
            .I(N__42668));
    InMux I__10435 (
            .O(N__42691),
            .I(N__42668));
    InMux I__10434 (
            .O(N__42690),
            .I(N__42668));
    InMux I__10433 (
            .O(N__42689),
            .I(N__42663));
    InMux I__10432 (
            .O(N__42688),
            .I(N__42657));
    InMux I__10431 (
            .O(N__42687),
            .I(N__42657));
    LocalMux I__10430 (
            .O(N__42684),
            .I(N__42654));
    InMux I__10429 (
            .O(N__42683),
            .I(N__42651));
    LocalMux I__10428 (
            .O(N__42680),
            .I(N__42648));
    LocalMux I__10427 (
            .O(N__42677),
            .I(N__42645));
    InMux I__10426 (
            .O(N__42676),
            .I(N__42639));
    InMux I__10425 (
            .O(N__42675),
            .I(N__42639));
    LocalMux I__10424 (
            .O(N__42668),
            .I(N__42636));
    InMux I__10423 (
            .O(N__42667),
            .I(N__42631));
    InMux I__10422 (
            .O(N__42666),
            .I(N__42631));
    LocalMux I__10421 (
            .O(N__42663),
            .I(N__42628));
    InMux I__10420 (
            .O(N__42662),
            .I(N__42625));
    LocalMux I__10419 (
            .O(N__42657),
            .I(N__42622));
    Span4Mux_v I__10418 (
            .O(N__42654),
            .I(N__42619));
    LocalMux I__10417 (
            .O(N__42651),
            .I(N__42616));
    Span4Mux_h I__10416 (
            .O(N__42648),
            .I(N__42611));
    Span4Mux_h I__10415 (
            .O(N__42645),
            .I(N__42611));
    InMux I__10414 (
            .O(N__42644),
            .I(N__42608));
    LocalMux I__10413 (
            .O(N__42639),
            .I(N__42603));
    Span4Mux_s2_h I__10412 (
            .O(N__42636),
            .I(N__42603));
    LocalMux I__10411 (
            .O(N__42631),
            .I(N__42598));
    Span4Mux_s2_h I__10410 (
            .O(N__42628),
            .I(N__42598));
    LocalMux I__10409 (
            .O(N__42625),
            .I(N__42595));
    Span4Mux_s3_h I__10408 (
            .O(N__42622),
            .I(N__42592));
    Span4Mux_h I__10407 (
            .O(N__42619),
            .I(N__42587));
    Span4Mux_v I__10406 (
            .O(N__42616),
            .I(N__42587));
    Span4Mux_v I__10405 (
            .O(N__42611),
            .I(N__42584));
    LocalMux I__10404 (
            .O(N__42608),
            .I(N__42577));
    Span4Mux_h I__10403 (
            .O(N__42603),
            .I(N__42577));
    Span4Mux_h I__10402 (
            .O(N__42598),
            .I(N__42577));
    Span4Mux_s3_h I__10401 (
            .O(N__42595),
            .I(N__42572));
    Span4Mux_v I__10400 (
            .O(N__42592),
            .I(N__42572));
    Odrv4 I__10399 (
            .O(N__42587),
            .I(\ALU.N_231_0 ));
    Odrv4 I__10398 (
            .O(N__42584),
            .I(\ALU.N_231_0 ));
    Odrv4 I__10397 (
            .O(N__42577),
            .I(\ALU.N_231_0 ));
    Odrv4 I__10396 (
            .O(N__42572),
            .I(\ALU.N_231_0 ));
    InMux I__10395 (
            .O(N__42563),
            .I(N__42560));
    LocalMux I__10394 (
            .O(N__42560),
            .I(N__42557));
    Odrv4 I__10393 (
            .O(N__42557),
            .I(\ALU.un9_addsub_cry_4_c_RNIL4NZ0Z97 ));
    InMux I__10392 (
            .O(N__42554),
            .I(N__42551));
    LocalMux I__10391 (
            .O(N__42551),
            .I(N__42548));
    Span4Mux_v I__10390 (
            .O(N__42548),
            .I(N__42545));
    Span4Mux_h I__10389 (
            .O(N__42545),
            .I(N__42542));
    Odrv4 I__10388 (
            .O(N__42542),
            .I(\ALU.un2_addsub_cry_4_c_RNI284VEZ0 ));
    InMux I__10387 (
            .O(N__42539),
            .I(N__42536));
    LocalMux I__10386 (
            .O(N__42536),
            .I(N__42533));
    Odrv4 I__10385 (
            .O(N__42533),
            .I(\ALU.un9_addsub_cry_5_c_RNI6SCFZ0Z7 ));
    InMux I__10384 (
            .O(N__42530),
            .I(N__42527));
    LocalMux I__10383 (
            .O(N__42527),
            .I(N__42523));
    CascadeMux I__10382 (
            .O(N__42526),
            .I(N__42519));
    Span4Mux_v I__10381 (
            .O(N__42523),
            .I(N__42514));
    InMux I__10380 (
            .O(N__42522),
            .I(N__42511));
    InMux I__10379 (
            .O(N__42519),
            .I(N__42508));
    InMux I__10378 (
            .O(N__42518),
            .I(N__42499));
    InMux I__10377 (
            .O(N__42517),
            .I(N__42496));
    Span4Mux_h I__10376 (
            .O(N__42514),
            .I(N__42490));
    LocalMux I__10375 (
            .O(N__42511),
            .I(N__42490));
    LocalMux I__10374 (
            .O(N__42508),
            .I(N__42487));
    InMux I__10373 (
            .O(N__42507),
            .I(N__42482));
    InMux I__10372 (
            .O(N__42506),
            .I(N__42482));
    InMux I__10371 (
            .O(N__42505),
            .I(N__42473));
    InMux I__10370 (
            .O(N__42504),
            .I(N__42473));
    InMux I__10369 (
            .O(N__42503),
            .I(N__42473));
    InMux I__10368 (
            .O(N__42502),
            .I(N__42473));
    LocalMux I__10367 (
            .O(N__42499),
            .I(N__42470));
    LocalMux I__10366 (
            .O(N__42496),
            .I(N__42467));
    InMux I__10365 (
            .O(N__42495),
            .I(N__42464));
    Span4Mux_v I__10364 (
            .O(N__42490),
            .I(N__42460));
    Span4Mux_v I__10363 (
            .O(N__42487),
            .I(N__42445));
    LocalMux I__10362 (
            .O(N__42482),
            .I(N__42445));
    LocalMux I__10361 (
            .O(N__42473),
            .I(N__42445));
    Span4Mux_h I__10360 (
            .O(N__42470),
            .I(N__42445));
    Span4Mux_v I__10359 (
            .O(N__42467),
            .I(N__42445));
    LocalMux I__10358 (
            .O(N__42464),
            .I(N__42445));
    InMux I__10357 (
            .O(N__42463),
            .I(N__42442));
    Span4Mux_h I__10356 (
            .O(N__42460),
            .I(N__42439));
    InMux I__10355 (
            .O(N__42459),
            .I(N__42436));
    InMux I__10354 (
            .O(N__42458),
            .I(N__42433));
    Span4Mux_v I__10353 (
            .O(N__42445),
            .I(N__42430));
    LocalMux I__10352 (
            .O(N__42442),
            .I(\ALU.addsub_0_sqmuxa ));
    Odrv4 I__10351 (
            .O(N__42439),
            .I(\ALU.addsub_0_sqmuxa ));
    LocalMux I__10350 (
            .O(N__42436),
            .I(\ALU.addsub_0_sqmuxa ));
    LocalMux I__10349 (
            .O(N__42433),
            .I(\ALU.addsub_0_sqmuxa ));
    Odrv4 I__10348 (
            .O(N__42430),
            .I(\ALU.addsub_0_sqmuxa ));
    InMux I__10347 (
            .O(N__42419),
            .I(N__42416));
    LocalMux I__10346 (
            .O(N__42416),
            .I(N__42413));
    Span4Mux_h I__10345 (
            .O(N__42413),
            .I(N__42410));
    Span4Mux_h I__10344 (
            .O(N__42410),
            .I(N__42407));
    Odrv4 I__10343 (
            .O(N__42407),
            .I(\ALU.un2_addsub_cry_5_c_RNIL7IGFZ0 ));
    InMux I__10342 (
            .O(N__42404),
            .I(N__42401));
    LocalMux I__10341 (
            .O(N__42401),
            .I(N__42398));
    Span4Mux_v I__10340 (
            .O(N__42398),
            .I(N__42395));
    Span4Mux_h I__10339 (
            .O(N__42395),
            .I(N__42392));
    Odrv4 I__10338 (
            .O(N__42392),
            .I(\ALU.N_422 ));
    CascadeMux I__10337 (
            .O(N__42389),
            .I(\ALU.d_RNIP43E91Z0Z_7_cascade_ ));
    InMux I__10336 (
            .O(N__42386),
            .I(N__42383));
    LocalMux I__10335 (
            .O(N__42383),
            .I(N__42380));
    Span4Mux_v I__10334 (
            .O(N__42380),
            .I(N__42377));
    Span4Mux_h I__10333 (
            .O(N__42377),
            .I(N__42374));
    Odrv4 I__10332 (
            .O(N__42374),
            .I(\ALU.d_RNIT87FA1Z0Z_7 ));
    InMux I__10331 (
            .O(N__42371),
            .I(N__42368));
    LocalMux I__10330 (
            .O(N__42368),
            .I(N__42365));
    Span4Mux_v I__10329 (
            .O(N__42365),
            .I(N__42362));
    Span4Mux_h I__10328 (
            .O(N__42362),
            .I(N__42359));
    Odrv4 I__10327 (
            .O(N__42359),
            .I(\ALU.madd_cry_5_THRU_CO ));
    CascadeMux I__10326 (
            .O(N__42356),
            .I(\ALU.a_15_m5_7_cascade_ ));
    InMux I__10325 (
            .O(N__42353),
            .I(N__42350));
    LocalMux I__10324 (
            .O(N__42350),
            .I(N__42346));
    InMux I__10323 (
            .O(N__42349),
            .I(N__42343));
    Span4Mux_v I__10322 (
            .O(N__42346),
            .I(N__42340));
    LocalMux I__10321 (
            .O(N__42343),
            .I(N__42337));
    Span4Mux_h I__10320 (
            .O(N__42340),
            .I(N__42332));
    Span4Mux_v I__10319 (
            .O(N__42337),
            .I(N__42332));
    Span4Mux_h I__10318 (
            .O(N__42332),
            .I(N__42329));
    Odrv4 I__10317 (
            .O(N__42329),
            .I(\ALU.madd_axb_6 ));
    InMux I__10316 (
            .O(N__42326),
            .I(N__42323));
    LocalMux I__10315 (
            .O(N__42323),
            .I(N__42318));
    InMux I__10314 (
            .O(N__42322),
            .I(N__42315));
    InMux I__10313 (
            .O(N__42321),
            .I(N__42312));
    Span4Mux_h I__10312 (
            .O(N__42318),
            .I(N__42308));
    LocalMux I__10311 (
            .O(N__42315),
            .I(N__42305));
    LocalMux I__10310 (
            .O(N__42312),
            .I(N__42302));
    InMux I__10309 (
            .O(N__42311),
            .I(N__42299));
    Span4Mux_h I__10308 (
            .O(N__42308),
            .I(N__42289));
    Span4Mux_v I__10307 (
            .O(N__42305),
            .I(N__42289));
    Span4Mux_v I__10306 (
            .O(N__42302),
            .I(N__42289));
    LocalMux I__10305 (
            .O(N__42299),
            .I(N__42286));
    InMux I__10304 (
            .O(N__42298),
            .I(N__42283));
    InMux I__10303 (
            .O(N__42297),
            .I(N__42280));
    InMux I__10302 (
            .O(N__42296),
            .I(N__42277));
    Odrv4 I__10301 (
            .O(N__42289),
            .I(\ALU.d_RNIO75MAZ0Z_0 ));
    Odrv12 I__10300 (
            .O(N__42286),
            .I(\ALU.d_RNIO75MAZ0Z_0 ));
    LocalMux I__10299 (
            .O(N__42283),
            .I(\ALU.d_RNIO75MAZ0Z_0 ));
    LocalMux I__10298 (
            .O(N__42280),
            .I(\ALU.d_RNIO75MAZ0Z_0 ));
    LocalMux I__10297 (
            .O(N__42277),
            .I(\ALU.d_RNIO75MAZ0Z_0 ));
    InMux I__10296 (
            .O(N__42266),
            .I(N__42261));
    InMux I__10295 (
            .O(N__42265),
            .I(N__42258));
    InMux I__10294 (
            .O(N__42264),
            .I(N__42255));
    LocalMux I__10293 (
            .O(N__42261),
            .I(N__42249));
    LocalMux I__10292 (
            .O(N__42258),
            .I(N__42246));
    LocalMux I__10291 (
            .O(N__42255),
            .I(N__42243));
    InMux I__10290 (
            .O(N__42254),
            .I(N__42240));
    InMux I__10289 (
            .O(N__42253),
            .I(N__42237));
    InMux I__10288 (
            .O(N__42252),
            .I(N__42234));
    Span4Mux_v I__10287 (
            .O(N__42249),
            .I(N__42228));
    Span4Mux_v I__10286 (
            .O(N__42246),
            .I(N__42228));
    Span4Mux_v I__10285 (
            .O(N__42243),
            .I(N__42225));
    LocalMux I__10284 (
            .O(N__42240),
            .I(N__42222));
    LocalMux I__10283 (
            .O(N__42237),
            .I(N__42219));
    LocalMux I__10282 (
            .O(N__42234),
            .I(N__42216));
    InMux I__10281 (
            .O(N__42233),
            .I(N__42213));
    Span4Mux_h I__10280 (
            .O(N__42228),
            .I(N__42210));
    Span4Mux_h I__10279 (
            .O(N__42225),
            .I(N__42199));
    Span4Mux_v I__10278 (
            .O(N__42222),
            .I(N__42199));
    Span4Mux_h I__10277 (
            .O(N__42219),
            .I(N__42199));
    Span4Mux_v I__10276 (
            .O(N__42216),
            .I(N__42199));
    LocalMux I__10275 (
            .O(N__42213),
            .I(N__42199));
    Odrv4 I__10274 (
            .O(N__42210),
            .I(\ALU.d_RNI9BO713Z0Z_0 ));
    Odrv4 I__10273 (
            .O(N__42199),
            .I(\ALU.d_RNI9BO713Z0Z_0 ));
    InMux I__10272 (
            .O(N__42194),
            .I(N__42190));
    InMux I__10271 (
            .O(N__42193),
            .I(N__42187));
    LocalMux I__10270 (
            .O(N__42190),
            .I(N__42184));
    LocalMux I__10269 (
            .O(N__42187),
            .I(N__42181));
    Span4Mux_h I__10268 (
            .O(N__42184),
            .I(N__42178));
    Span4Mux_h I__10267 (
            .O(N__42181),
            .I(N__42175));
    Span4Mux_h I__10266 (
            .O(N__42178),
            .I(N__42172));
    Span4Mux_h I__10265 (
            .O(N__42175),
            .I(N__42169));
    Odrv4 I__10264 (
            .O(N__42172),
            .I(\ALU.dZ0Z_0 ));
    Odrv4 I__10263 (
            .O(N__42169),
            .I(\ALU.dZ0Z_0 ));
    InMux I__10262 (
            .O(N__42164),
            .I(N__42158));
    InMux I__10261 (
            .O(N__42163),
            .I(N__42155));
    InMux I__10260 (
            .O(N__42162),
            .I(N__42152));
    InMux I__10259 (
            .O(N__42161),
            .I(N__42147));
    LocalMux I__10258 (
            .O(N__42158),
            .I(N__42139));
    LocalMux I__10257 (
            .O(N__42155),
            .I(N__42139));
    LocalMux I__10256 (
            .O(N__42152),
            .I(N__42139));
    InMux I__10255 (
            .O(N__42151),
            .I(N__42136));
    InMux I__10254 (
            .O(N__42150),
            .I(N__42133));
    LocalMux I__10253 (
            .O(N__42147),
            .I(N__42130));
    InMux I__10252 (
            .O(N__42146),
            .I(N__42127));
    Span4Mux_v I__10251 (
            .O(N__42139),
            .I(N__42119));
    LocalMux I__10250 (
            .O(N__42136),
            .I(N__42119));
    LocalMux I__10249 (
            .O(N__42133),
            .I(N__42119));
    Span4Mux_h I__10248 (
            .O(N__42130),
            .I(N__42114));
    LocalMux I__10247 (
            .O(N__42127),
            .I(N__42114));
    InMux I__10246 (
            .O(N__42126),
            .I(N__42111));
    Span4Mux_h I__10245 (
            .O(N__42119),
            .I(N__42108));
    Sp12to4 I__10244 (
            .O(N__42114),
            .I(N__42103));
    LocalMux I__10243 (
            .O(N__42111),
            .I(N__42103));
    Odrv4 I__10242 (
            .O(N__42108),
            .I(\ALU.un9_addsub_cry_1_c_RNIM56ULZ0 ));
    Odrv12 I__10241 (
            .O(N__42103),
            .I(\ALU.un9_addsub_cry_1_c_RNIM56ULZ0 ));
    InMux I__10240 (
            .O(N__42098),
            .I(N__42093));
    InMux I__10239 (
            .O(N__42097),
            .I(N__42089));
    InMux I__10238 (
            .O(N__42096),
            .I(N__42086));
    LocalMux I__10237 (
            .O(N__42093),
            .I(N__42083));
    InMux I__10236 (
            .O(N__42092),
            .I(N__42080));
    LocalMux I__10235 (
            .O(N__42089),
            .I(N__42073));
    LocalMux I__10234 (
            .O(N__42086),
            .I(N__42073));
    Span4Mux_v I__10233 (
            .O(N__42083),
            .I(N__42069));
    LocalMux I__10232 (
            .O(N__42080),
            .I(N__42066));
    InMux I__10231 (
            .O(N__42079),
            .I(N__42063));
    InMux I__10230 (
            .O(N__42078),
            .I(N__42060));
    Span4Mux_v I__10229 (
            .O(N__42073),
            .I(N__42057));
    InMux I__10228 (
            .O(N__42072),
            .I(N__42054));
    Span4Mux_h I__10227 (
            .O(N__42069),
            .I(N__42045));
    Span4Mux_v I__10226 (
            .O(N__42066),
            .I(N__42045));
    LocalMux I__10225 (
            .O(N__42063),
            .I(N__42045));
    LocalMux I__10224 (
            .O(N__42060),
            .I(N__42045));
    Odrv4 I__10223 (
            .O(N__42057),
            .I(\ALU.d_RNIIFMN04Z0Z_2 ));
    LocalMux I__10222 (
            .O(N__42054),
            .I(\ALU.d_RNIIFMN04Z0Z_2 ));
    Odrv4 I__10221 (
            .O(N__42045),
            .I(\ALU.d_RNIIFMN04Z0Z_2 ));
    InMux I__10220 (
            .O(N__42038),
            .I(N__42035));
    LocalMux I__10219 (
            .O(N__42035),
            .I(N__42031));
    InMux I__10218 (
            .O(N__42034),
            .I(N__42028));
    Span4Mux_v I__10217 (
            .O(N__42031),
            .I(N__42023));
    LocalMux I__10216 (
            .O(N__42028),
            .I(N__42023));
    Span4Mux_v I__10215 (
            .O(N__42023),
            .I(N__42020));
    Odrv4 I__10214 (
            .O(N__42020),
            .I(\ALU.dZ0Z_2 ));
    InMux I__10213 (
            .O(N__42017),
            .I(N__42006));
    InMux I__10212 (
            .O(N__42016),
            .I(N__42006));
    InMux I__10211 (
            .O(N__42015),
            .I(N__42002));
    InMux I__10210 (
            .O(N__42014),
            .I(N__41999));
    InMux I__10209 (
            .O(N__42013),
            .I(N__41996));
    InMux I__10208 (
            .O(N__42012),
            .I(N__41989));
    InMux I__10207 (
            .O(N__42011),
            .I(N__41986));
    LocalMux I__10206 (
            .O(N__42006),
            .I(N__41983));
    InMux I__10205 (
            .O(N__42005),
            .I(N__41980));
    LocalMux I__10204 (
            .O(N__42002),
            .I(N__41966));
    LocalMux I__10203 (
            .O(N__41999),
            .I(N__41966));
    LocalMux I__10202 (
            .O(N__41996),
            .I(N__41966));
    InMux I__10201 (
            .O(N__41995),
            .I(N__41963));
    InMux I__10200 (
            .O(N__41994),
            .I(N__41960));
    InMux I__10199 (
            .O(N__41993),
            .I(N__41956));
    InMux I__10198 (
            .O(N__41992),
            .I(N__41952));
    LocalMux I__10197 (
            .O(N__41989),
            .I(N__41947));
    LocalMux I__10196 (
            .O(N__41986),
            .I(N__41947));
    Span4Mux_v I__10195 (
            .O(N__41983),
            .I(N__41944));
    LocalMux I__10194 (
            .O(N__41980),
            .I(N__41938));
    InMux I__10193 (
            .O(N__41979),
            .I(N__41931));
    InMux I__10192 (
            .O(N__41978),
            .I(N__41931));
    InMux I__10191 (
            .O(N__41977),
            .I(N__41931));
    InMux I__10190 (
            .O(N__41976),
            .I(N__41928));
    CascadeMux I__10189 (
            .O(N__41975),
            .I(N__41923));
    InMux I__10188 (
            .O(N__41974),
            .I(N__41920));
    InMux I__10187 (
            .O(N__41973),
            .I(N__41916));
    Span4Mux_h I__10186 (
            .O(N__41966),
            .I(N__41911));
    LocalMux I__10185 (
            .O(N__41963),
            .I(N__41911));
    LocalMux I__10184 (
            .O(N__41960),
            .I(N__41908));
    InMux I__10183 (
            .O(N__41959),
            .I(N__41905));
    LocalMux I__10182 (
            .O(N__41956),
            .I(N__41902));
    InMux I__10181 (
            .O(N__41955),
            .I(N__41899));
    LocalMux I__10180 (
            .O(N__41952),
            .I(N__41892));
    Span4Mux_v I__10179 (
            .O(N__41947),
            .I(N__41892));
    Span4Mux_v I__10178 (
            .O(N__41944),
            .I(N__41892));
    InMux I__10177 (
            .O(N__41943),
            .I(N__41887));
    InMux I__10176 (
            .O(N__41942),
            .I(N__41887));
    InMux I__10175 (
            .O(N__41941),
            .I(N__41884));
    Span4Mux_h I__10174 (
            .O(N__41938),
            .I(N__41879));
    LocalMux I__10173 (
            .O(N__41931),
            .I(N__41874));
    LocalMux I__10172 (
            .O(N__41928),
            .I(N__41874));
    InMux I__10171 (
            .O(N__41927),
            .I(N__41871));
    InMux I__10170 (
            .O(N__41926),
            .I(N__41868));
    InMux I__10169 (
            .O(N__41923),
            .I(N__41865));
    LocalMux I__10168 (
            .O(N__41920),
            .I(N__41857));
    InMux I__10167 (
            .O(N__41919),
            .I(N__41854));
    LocalMux I__10166 (
            .O(N__41916),
            .I(N__41851));
    Span4Mux_v I__10165 (
            .O(N__41911),
            .I(N__41848));
    Span4Mux_s2_h I__10164 (
            .O(N__41908),
            .I(N__41843));
    LocalMux I__10163 (
            .O(N__41905),
            .I(N__41843));
    Span4Mux_h I__10162 (
            .O(N__41902),
            .I(N__41840));
    LocalMux I__10161 (
            .O(N__41899),
            .I(N__41833));
    Sp12to4 I__10160 (
            .O(N__41892),
            .I(N__41833));
    LocalMux I__10159 (
            .O(N__41887),
            .I(N__41833));
    LocalMux I__10158 (
            .O(N__41884),
            .I(N__41830));
    InMux I__10157 (
            .O(N__41883),
            .I(N__41825));
    InMux I__10156 (
            .O(N__41882),
            .I(N__41825));
    Span4Mux_h I__10155 (
            .O(N__41879),
            .I(N__41820));
    Span4Mux_v I__10154 (
            .O(N__41874),
            .I(N__41820));
    LocalMux I__10153 (
            .O(N__41871),
            .I(N__41813));
    LocalMux I__10152 (
            .O(N__41868),
            .I(N__41813));
    LocalMux I__10151 (
            .O(N__41865),
            .I(N__41813));
    InMux I__10150 (
            .O(N__41864),
            .I(N__41810));
    InMux I__10149 (
            .O(N__41863),
            .I(N__41804));
    InMux I__10148 (
            .O(N__41862),
            .I(N__41804));
    InMux I__10147 (
            .O(N__41861),
            .I(N__41799));
    InMux I__10146 (
            .O(N__41860),
            .I(N__41799));
    Span12Mux_v I__10145 (
            .O(N__41857),
            .I(N__41794));
    LocalMux I__10144 (
            .O(N__41854),
            .I(N__41794));
    Span4Mux_h I__10143 (
            .O(N__41851),
            .I(N__41787));
    Span4Mux_v I__10142 (
            .O(N__41848),
            .I(N__41787));
    Span4Mux_h I__10141 (
            .O(N__41843),
            .I(N__41787));
    Sp12to4 I__10140 (
            .O(N__41840),
            .I(N__41782));
    Span12Mux_s6_h I__10139 (
            .O(N__41833),
            .I(N__41782));
    Span4Mux_h I__10138 (
            .O(N__41830),
            .I(N__41779));
    LocalMux I__10137 (
            .O(N__41825),
            .I(N__41776));
    Span4Mux_v I__10136 (
            .O(N__41820),
            .I(N__41769));
    Span4Mux_h I__10135 (
            .O(N__41813),
            .I(N__41769));
    LocalMux I__10134 (
            .O(N__41810),
            .I(N__41769));
    InMux I__10133 (
            .O(N__41809),
            .I(N__41766));
    LocalMux I__10132 (
            .O(N__41804),
            .I(\ALU.aluOut_3 ));
    LocalMux I__10131 (
            .O(N__41799),
            .I(\ALU.aluOut_3 ));
    Odrv12 I__10130 (
            .O(N__41794),
            .I(\ALU.aluOut_3 ));
    Odrv4 I__10129 (
            .O(N__41787),
            .I(\ALU.aluOut_3 ));
    Odrv12 I__10128 (
            .O(N__41782),
            .I(\ALU.aluOut_3 ));
    Odrv4 I__10127 (
            .O(N__41779),
            .I(\ALU.aluOut_3 ));
    Odrv4 I__10126 (
            .O(N__41776),
            .I(\ALU.aluOut_3 ));
    Odrv4 I__10125 (
            .O(N__41769),
            .I(\ALU.aluOut_3 ));
    LocalMux I__10124 (
            .O(N__41766),
            .I(\ALU.aluOut_3 ));
    CascadeMux I__10123 (
            .O(N__41747),
            .I(N__41744));
    InMux I__10122 (
            .O(N__41744),
            .I(N__41741));
    LocalMux I__10121 (
            .O(N__41741),
            .I(\ALU.a_15_m2_ns_1Z0Z_3 ));
    InMux I__10120 (
            .O(N__41738),
            .I(N__41730));
    InMux I__10119 (
            .O(N__41737),
            .I(N__41730));
    InMux I__10118 (
            .O(N__41736),
            .I(N__41727));
    InMux I__10117 (
            .O(N__41735),
            .I(N__41723));
    LocalMux I__10116 (
            .O(N__41730),
            .I(N__41716));
    LocalMux I__10115 (
            .O(N__41727),
            .I(N__41713));
    InMux I__10114 (
            .O(N__41726),
            .I(N__41710));
    LocalMux I__10113 (
            .O(N__41723),
            .I(N__41707));
    InMux I__10112 (
            .O(N__41722),
            .I(N__41701));
    InMux I__10111 (
            .O(N__41721),
            .I(N__41696));
    InMux I__10110 (
            .O(N__41720),
            .I(N__41696));
    InMux I__10109 (
            .O(N__41719),
            .I(N__41691));
    Span4Mux_s2_h I__10108 (
            .O(N__41716),
            .I(N__41688));
    Span4Mux_v I__10107 (
            .O(N__41713),
            .I(N__41685));
    LocalMux I__10106 (
            .O(N__41710),
            .I(N__41682));
    Span4Mux_v I__10105 (
            .O(N__41707),
            .I(N__41679));
    InMux I__10104 (
            .O(N__41706),
            .I(N__41676));
    InMux I__10103 (
            .O(N__41705),
            .I(N__41671));
    InMux I__10102 (
            .O(N__41704),
            .I(N__41671));
    LocalMux I__10101 (
            .O(N__41701),
            .I(N__41668));
    LocalMux I__10100 (
            .O(N__41696),
            .I(N__41664));
    InMux I__10099 (
            .O(N__41695),
            .I(N__41659));
    InMux I__10098 (
            .O(N__41694),
            .I(N__41659));
    LocalMux I__10097 (
            .O(N__41691),
            .I(N__41654));
    Span4Mux_h I__10096 (
            .O(N__41688),
            .I(N__41654));
    Span4Mux_v I__10095 (
            .O(N__41685),
            .I(N__41649));
    Span4Mux_v I__10094 (
            .O(N__41682),
            .I(N__41649));
    Span4Mux_v I__10093 (
            .O(N__41679),
            .I(N__41646));
    LocalMux I__10092 (
            .O(N__41676),
            .I(N__41641));
    LocalMux I__10091 (
            .O(N__41671),
            .I(N__41641));
    Span12Mux_s6_h I__10090 (
            .O(N__41668),
            .I(N__41638));
    InMux I__10089 (
            .O(N__41667),
            .I(N__41635));
    Span4Mux_h I__10088 (
            .O(N__41664),
            .I(N__41628));
    LocalMux I__10087 (
            .O(N__41659),
            .I(N__41628));
    Span4Mux_v I__10086 (
            .O(N__41654),
            .I(N__41628));
    Span4Mux_h I__10085 (
            .O(N__41649),
            .I(N__41625));
    Span4Mux_h I__10084 (
            .O(N__41646),
            .I(N__41620));
    Span4Mux_v I__10083 (
            .O(N__41641),
            .I(N__41620));
    Odrv12 I__10082 (
            .O(N__41638),
            .I(\ALU.N_237_0 ));
    LocalMux I__10081 (
            .O(N__41635),
            .I(\ALU.N_237_0 ));
    Odrv4 I__10080 (
            .O(N__41628),
            .I(\ALU.N_237_0 ));
    Odrv4 I__10079 (
            .O(N__41625),
            .I(\ALU.N_237_0 ));
    Odrv4 I__10078 (
            .O(N__41620),
            .I(\ALU.N_237_0 ));
    CascadeMux I__10077 (
            .O(N__41609),
            .I(\ALU.a_15_m2_3_cascade_ ));
    InMux I__10076 (
            .O(N__41606),
            .I(N__41603));
    LocalMux I__10075 (
            .O(N__41603),
            .I(N__41600));
    Span4Mux_h I__10074 (
            .O(N__41600),
            .I(N__41597));
    Span4Mux_h I__10073 (
            .O(N__41597),
            .I(N__41594));
    Span4Mux_v I__10072 (
            .O(N__41594),
            .I(N__41591));
    Odrv4 I__10071 (
            .O(N__41591),
            .I(\ALU.lshift_1_3 ));
    InMux I__10070 (
            .O(N__41588),
            .I(N__41585));
    LocalMux I__10069 (
            .O(N__41585),
            .I(\ALU.d_RNI95MLPZ0Z_3 ));
    InMux I__10068 (
            .O(N__41582),
            .I(N__41579));
    LocalMux I__10067 (
            .O(N__41579),
            .I(N__41576));
    Odrv12 I__10066 (
            .O(N__41576),
            .I(\ALU.mult_3 ));
    InMux I__10065 (
            .O(N__41573),
            .I(N__41570));
    LocalMux I__10064 (
            .O(N__41570),
            .I(\ALU.a_15_m5_3 ));
    InMux I__10063 (
            .O(N__41567),
            .I(N__41564));
    LocalMux I__10062 (
            .O(N__41564),
            .I(N__41560));
    CascadeMux I__10061 (
            .O(N__41563),
            .I(N__41557));
    Span4Mux_v I__10060 (
            .O(N__41560),
            .I(N__41554));
    InMux I__10059 (
            .O(N__41557),
            .I(N__41551));
    Span4Mux_h I__10058 (
            .O(N__41554),
            .I(N__41548));
    LocalMux I__10057 (
            .O(N__41551),
            .I(N__41545));
    Span4Mux_h I__10056 (
            .O(N__41548),
            .I(N__41539));
    Span4Mux_v I__10055 (
            .O(N__41545),
            .I(N__41539));
    CascadeMux I__10054 (
            .O(N__41544),
            .I(N__41535));
    Span4Mux_h I__10053 (
            .O(N__41539),
            .I(N__41531));
    InMux I__10052 (
            .O(N__41538),
            .I(N__41526));
    InMux I__10051 (
            .O(N__41535),
            .I(N__41526));
    InMux I__10050 (
            .O(N__41534),
            .I(N__41523));
    Span4Mux_v I__10049 (
            .O(N__41531),
            .I(N__41520));
    LocalMux I__10048 (
            .O(N__41526),
            .I(N__41517));
    LocalMux I__10047 (
            .O(N__41523),
            .I(RXbuffer_2));
    Odrv4 I__10046 (
            .O(N__41520),
            .I(RXbuffer_2));
    Odrv4 I__10045 (
            .O(N__41517),
            .I(RXbuffer_2));
    CascadeMux I__10044 (
            .O(N__41510),
            .I(N__41503));
    CascadeMux I__10043 (
            .O(N__41509),
            .I(N__41497));
    CascadeMux I__10042 (
            .O(N__41508),
            .I(N__41494));
    CascadeMux I__10041 (
            .O(N__41507),
            .I(N__41491));
    InMux I__10040 (
            .O(N__41506),
            .I(N__41479));
    InMux I__10039 (
            .O(N__41503),
            .I(N__41479));
    InMux I__10038 (
            .O(N__41502),
            .I(N__41479));
    InMux I__10037 (
            .O(N__41501),
            .I(N__41471));
    InMux I__10036 (
            .O(N__41500),
            .I(N__41468));
    InMux I__10035 (
            .O(N__41497),
            .I(N__41458));
    InMux I__10034 (
            .O(N__41494),
            .I(N__41458));
    InMux I__10033 (
            .O(N__41491),
            .I(N__41458));
    InMux I__10032 (
            .O(N__41490),
            .I(N__41458));
    InMux I__10031 (
            .O(N__41489),
            .I(N__41455));
    InMux I__10030 (
            .O(N__41488),
            .I(N__41448));
    InMux I__10029 (
            .O(N__41487),
            .I(N__41448));
    InMux I__10028 (
            .O(N__41486),
            .I(N__41448));
    LocalMux I__10027 (
            .O(N__41479),
            .I(N__41445));
    CascadeMux I__10026 (
            .O(N__41478),
            .I(N__41442));
    CascadeMux I__10025 (
            .O(N__41477),
            .I(N__41439));
    CascadeMux I__10024 (
            .O(N__41476),
            .I(N__41435));
    CascadeMux I__10023 (
            .O(N__41475),
            .I(N__41432));
    InMux I__10022 (
            .O(N__41474),
            .I(N__41420));
    LocalMux I__10021 (
            .O(N__41471),
            .I(N__41417));
    LocalMux I__10020 (
            .O(N__41468),
            .I(N__41414));
    InMux I__10019 (
            .O(N__41467),
            .I(N__41410));
    LocalMux I__10018 (
            .O(N__41458),
            .I(N__41400));
    LocalMux I__10017 (
            .O(N__41455),
            .I(N__41400));
    LocalMux I__10016 (
            .O(N__41448),
            .I(N__41400));
    Span4Mux_v I__10015 (
            .O(N__41445),
            .I(N__41400));
    InMux I__10014 (
            .O(N__41442),
            .I(N__41396));
    InMux I__10013 (
            .O(N__41439),
            .I(N__41391));
    InMux I__10012 (
            .O(N__41438),
            .I(N__41391));
    InMux I__10011 (
            .O(N__41435),
            .I(N__41382));
    InMux I__10010 (
            .O(N__41432),
            .I(N__41382));
    InMux I__10009 (
            .O(N__41431),
            .I(N__41382));
    InMux I__10008 (
            .O(N__41430),
            .I(N__41382));
    InMux I__10007 (
            .O(N__41429),
            .I(N__41375));
    InMux I__10006 (
            .O(N__41428),
            .I(N__41375));
    InMux I__10005 (
            .O(N__41427),
            .I(N__41375));
    InMux I__10004 (
            .O(N__41426),
            .I(N__41366));
    InMux I__10003 (
            .O(N__41425),
            .I(N__41366));
    InMux I__10002 (
            .O(N__41424),
            .I(N__41366));
    InMux I__10001 (
            .O(N__41423),
            .I(N__41366));
    LocalMux I__10000 (
            .O(N__41420),
            .I(N__41363));
    Span4Mux_h I__9999 (
            .O(N__41417),
            .I(N__41360));
    Span4Mux_v I__9998 (
            .O(N__41414),
            .I(N__41356));
    InMux I__9997 (
            .O(N__41413),
            .I(N__41353));
    LocalMux I__9996 (
            .O(N__41410),
            .I(N__41350));
    InMux I__9995 (
            .O(N__41409),
            .I(N__41347));
    Span4Mux_v I__9994 (
            .O(N__41400),
            .I(N__41344));
    InMux I__9993 (
            .O(N__41399),
            .I(N__41341));
    LocalMux I__9992 (
            .O(N__41396),
            .I(N__41335));
    LocalMux I__9991 (
            .O(N__41391),
            .I(N__41332));
    LocalMux I__9990 (
            .O(N__41382),
            .I(N__41329));
    LocalMux I__9989 (
            .O(N__41375),
            .I(N__41324));
    LocalMux I__9988 (
            .O(N__41366),
            .I(N__41324));
    Span4Mux_h I__9987 (
            .O(N__41363),
            .I(N__41319));
    Span4Mux_h I__9986 (
            .O(N__41360),
            .I(N__41319));
    InMux I__9985 (
            .O(N__41359),
            .I(N__41316));
    Span4Mux_h I__9984 (
            .O(N__41356),
            .I(N__41313));
    LocalMux I__9983 (
            .O(N__41353),
            .I(N__41306));
    Span4Mux_v I__9982 (
            .O(N__41350),
            .I(N__41306));
    LocalMux I__9981 (
            .O(N__41347),
            .I(N__41306));
    Span4Mux_h I__9980 (
            .O(N__41344),
            .I(N__41301));
    LocalMux I__9979 (
            .O(N__41341),
            .I(N__41301));
    InMux I__9978 (
            .O(N__41340),
            .I(N__41294));
    InMux I__9977 (
            .O(N__41339),
            .I(N__41294));
    InMux I__9976 (
            .O(N__41338),
            .I(N__41294));
    Span4Mux_h I__9975 (
            .O(N__41335),
            .I(N__41289));
    Span4Mux_h I__9974 (
            .O(N__41332),
            .I(N__41286));
    Span4Mux_s3_v I__9973 (
            .O(N__41329),
            .I(N__41281));
    Span4Mux_s2_h I__9972 (
            .O(N__41324),
            .I(N__41281));
    Span4Mux_v I__9971 (
            .O(N__41319),
            .I(N__41278));
    LocalMux I__9970 (
            .O(N__41316),
            .I(N__41271));
    Span4Mux_v I__9969 (
            .O(N__41313),
            .I(N__41271));
    Span4Mux_h I__9968 (
            .O(N__41306),
            .I(N__41271));
    Span4Mux_v I__9967 (
            .O(N__41301),
            .I(N__41266));
    LocalMux I__9966 (
            .O(N__41294),
            .I(N__41266));
    InMux I__9965 (
            .O(N__41293),
            .I(N__41261));
    InMux I__9964 (
            .O(N__41292),
            .I(N__41261));
    Span4Mux_v I__9963 (
            .O(N__41289),
            .I(N__41258));
    Span4Mux_v I__9962 (
            .O(N__41286),
            .I(N__41255));
    Span4Mux_h I__9961 (
            .O(N__41281),
            .I(N__41252));
    Span4Mux_v I__9960 (
            .O(N__41278),
            .I(N__41249));
    Span4Mux_v I__9959 (
            .O(N__41271),
            .I(N__41244));
    Span4Mux_s0_v I__9958 (
            .O(N__41266),
            .I(N__41244));
    LocalMux I__9957 (
            .O(N__41261),
            .I(testStateZ0Z_1));
    Odrv4 I__9956 (
            .O(N__41258),
            .I(testStateZ0Z_1));
    Odrv4 I__9955 (
            .O(N__41255),
            .I(testStateZ0Z_1));
    Odrv4 I__9954 (
            .O(N__41252),
            .I(testStateZ0Z_1));
    Odrv4 I__9953 (
            .O(N__41249),
            .I(testStateZ0Z_1));
    Odrv4 I__9952 (
            .O(N__41244),
            .I(testStateZ0Z_1));
    InMux I__9951 (
            .O(N__41231),
            .I(N__41227));
    InMux I__9950 (
            .O(N__41230),
            .I(N__41224));
    LocalMux I__9949 (
            .O(N__41227),
            .I(N__41221));
    LocalMux I__9948 (
            .O(N__41224),
            .I(N__41215));
    Span4Mux_v I__9947 (
            .O(N__41221),
            .I(N__41211));
    InMux I__9946 (
            .O(N__41220),
            .I(N__41208));
    InMux I__9945 (
            .O(N__41219),
            .I(N__41194));
    InMux I__9944 (
            .O(N__41218),
            .I(N__41194));
    Span4Mux_v I__9943 (
            .O(N__41215),
            .I(N__41191));
    InMux I__9942 (
            .O(N__41214),
            .I(N__41188));
    Span4Mux_v I__9941 (
            .O(N__41211),
            .I(N__41183));
    LocalMux I__9940 (
            .O(N__41208),
            .I(N__41183));
    InMux I__9939 (
            .O(N__41207),
            .I(N__41178));
    InMux I__9938 (
            .O(N__41206),
            .I(N__41178));
    InMux I__9937 (
            .O(N__41205),
            .I(N__41163));
    InMux I__9936 (
            .O(N__41204),
            .I(N__41163));
    InMux I__9935 (
            .O(N__41203),
            .I(N__41163));
    InMux I__9934 (
            .O(N__41202),
            .I(N__41163));
    InMux I__9933 (
            .O(N__41201),
            .I(N__41163));
    InMux I__9932 (
            .O(N__41200),
            .I(N__41163));
    InMux I__9931 (
            .O(N__41199),
            .I(N__41163));
    LocalMux I__9930 (
            .O(N__41194),
            .I(N__41160));
    Sp12to4 I__9929 (
            .O(N__41191),
            .I(N__41156));
    LocalMux I__9928 (
            .O(N__41188),
            .I(N__41153));
    Span4Mux_h I__9927 (
            .O(N__41183),
            .I(N__41150));
    LocalMux I__9926 (
            .O(N__41178),
            .I(N__41147));
    LocalMux I__9925 (
            .O(N__41163),
            .I(N__41142));
    Sp12to4 I__9924 (
            .O(N__41160),
            .I(N__41142));
    InMux I__9923 (
            .O(N__41159),
            .I(N__41139));
    Span12Mux_v I__9922 (
            .O(N__41156),
            .I(N__41136));
    Span4Mux_v I__9921 (
            .O(N__41153),
            .I(N__41133));
    Span4Mux_h I__9920 (
            .O(N__41150),
            .I(N__41128));
    Span4Mux_h I__9919 (
            .O(N__41147),
            .I(N__41128));
    Span12Mux_s5_h I__9918 (
            .O(N__41142),
            .I(N__41123));
    LocalMux I__9917 (
            .O(N__41139),
            .I(N__41123));
    Odrv12 I__9916 (
            .O(N__41136),
            .I(\ALU.N_58_0 ));
    Odrv4 I__9915 (
            .O(N__41133),
            .I(\ALU.N_58_0 ));
    Odrv4 I__9914 (
            .O(N__41128),
            .I(\ALU.N_58_0 ));
    Odrv12 I__9913 (
            .O(N__41123),
            .I(\ALU.N_58_0 ));
    InMux I__9912 (
            .O(N__41114),
            .I(N__41109));
    CascadeMux I__9911 (
            .O(N__41113),
            .I(N__41104));
    InMux I__9910 (
            .O(N__41112),
            .I(N__41101));
    LocalMux I__9909 (
            .O(N__41109),
            .I(N__41098));
    CascadeMux I__9908 (
            .O(N__41108),
            .I(N__41095));
    InMux I__9907 (
            .O(N__41107),
            .I(N__41090));
    InMux I__9906 (
            .O(N__41104),
            .I(N__41090));
    LocalMux I__9905 (
            .O(N__41101),
            .I(N__41087));
    Span4Mux_v I__9904 (
            .O(N__41098),
            .I(N__41084));
    InMux I__9903 (
            .O(N__41095),
            .I(N__41081));
    LocalMux I__9902 (
            .O(N__41090),
            .I(N__41078));
    Span12Mux_s8_h I__9901 (
            .O(N__41087),
            .I(N__41075));
    Span4Mux_h I__9900 (
            .O(N__41084),
            .I(N__41072));
    LocalMux I__9899 (
            .O(N__41081),
            .I(testWordZ0Z_10));
    Odrv4 I__9898 (
            .O(N__41078),
            .I(testWordZ0Z_10));
    Odrv12 I__9897 (
            .O(N__41075),
            .I(testWordZ0Z_10));
    Odrv4 I__9896 (
            .O(N__41072),
            .I(testWordZ0Z_10));
    CEMux I__9895 (
            .O(N__41063),
            .I(N__41027));
    CEMux I__9894 (
            .O(N__41062),
            .I(N__41027));
    CEMux I__9893 (
            .O(N__41061),
            .I(N__41027));
    CEMux I__9892 (
            .O(N__41060),
            .I(N__41027));
    CEMux I__9891 (
            .O(N__41059),
            .I(N__41027));
    CEMux I__9890 (
            .O(N__41058),
            .I(N__41027));
    CEMux I__9889 (
            .O(N__41057),
            .I(N__41027));
    CEMux I__9888 (
            .O(N__41056),
            .I(N__41027));
    CEMux I__9887 (
            .O(N__41055),
            .I(N__41027));
    CEMux I__9886 (
            .O(N__41054),
            .I(N__41027));
    CEMux I__9885 (
            .O(N__41053),
            .I(N__41027));
    CEMux I__9884 (
            .O(N__41052),
            .I(N__41027));
    GlobalMux I__9883 (
            .O(N__41027),
            .I(N__41024));
    gio2CtrlBuf I__9882 (
            .O(N__41024),
            .I(testState_i_g_2));
    InMux I__9881 (
            .O(N__41021),
            .I(N__41018));
    LocalMux I__9880 (
            .O(N__41018),
            .I(N__41015));
    Odrv12 I__9879 (
            .O(N__41015),
            .I(\ALU.un9_addsub_cry_0_c_RNI2UZ0Z096 ));
    InMux I__9878 (
            .O(N__41012),
            .I(N__41009));
    LocalMux I__9877 (
            .O(N__41009),
            .I(N__41006));
    Span12Mux_h I__9876 (
            .O(N__41006),
            .I(N__41003));
    Odrv12 I__9875 (
            .O(N__41003),
            .I(\ALU.un2_addsub_cry_0_c_RNI5MA0EZ0 ));
    InMux I__9874 (
            .O(N__41000),
            .I(N__40995));
    InMux I__9873 (
            .O(N__40999),
            .I(N__40991));
    InMux I__9872 (
            .O(N__40998),
            .I(N__40988));
    LocalMux I__9871 (
            .O(N__40995),
            .I(N__40985));
    InMux I__9870 (
            .O(N__40994),
            .I(N__40982));
    LocalMux I__9869 (
            .O(N__40991),
            .I(N__40976));
    LocalMux I__9868 (
            .O(N__40988),
            .I(N__40969));
    Span4Mux_h I__9867 (
            .O(N__40985),
            .I(N__40969));
    LocalMux I__9866 (
            .O(N__40982),
            .I(N__40969));
    InMux I__9865 (
            .O(N__40981),
            .I(N__40966));
    InMux I__9864 (
            .O(N__40980),
            .I(N__40963));
    InMux I__9863 (
            .O(N__40979),
            .I(N__40960));
    Span4Mux_h I__9862 (
            .O(N__40976),
            .I(N__40956));
    Span4Mux_v I__9861 (
            .O(N__40969),
            .I(N__40951));
    LocalMux I__9860 (
            .O(N__40966),
            .I(N__40951));
    LocalMux I__9859 (
            .O(N__40963),
            .I(N__40946));
    LocalMux I__9858 (
            .O(N__40960),
            .I(N__40946));
    InMux I__9857 (
            .O(N__40959),
            .I(N__40943));
    Span4Mux_v I__9856 (
            .O(N__40956),
            .I(N__40940));
    Span4Mux_h I__9855 (
            .O(N__40951),
            .I(N__40937));
    Span4Mux_v I__9854 (
            .O(N__40946),
            .I(N__40932));
    LocalMux I__9853 (
            .O(N__40943),
            .I(N__40932));
    Odrv4 I__9852 (
            .O(N__40940),
            .I(\ALU.un9_addsub_cry_0_c_RNIEMTLKZ0 ));
    Odrv4 I__9851 (
            .O(N__40937),
            .I(\ALU.un9_addsub_cry_0_c_RNIEMTLKZ0 ));
    Odrv4 I__9850 (
            .O(N__40932),
            .I(\ALU.un9_addsub_cry_0_c_RNIEMTLKZ0 ));
    InMux I__9849 (
            .O(N__40925),
            .I(N__40922));
    LocalMux I__9848 (
            .O(N__40922),
            .I(N__40919));
    Odrv4 I__9847 (
            .O(N__40919),
            .I(\ALU.un9_addsub_cry_1_c_RNI6TDZ0Z17 ));
    InMux I__9846 (
            .O(N__40916),
            .I(N__40913));
    LocalMux I__9845 (
            .O(N__40913),
            .I(N__40910));
    Span4Mux_v I__9844 (
            .O(N__40910),
            .I(N__40907));
    Sp12to4 I__9843 (
            .O(N__40907),
            .I(N__40904));
    Odrv12 I__9842 (
            .O(N__40904),
            .I(\ALU.un2_addsub_cry_1_c_RNI966GEZ0 ));
    InMux I__9841 (
            .O(N__40901),
            .I(N__40898));
    LocalMux I__9840 (
            .O(N__40898),
            .I(N__40895));
    Odrv4 I__9839 (
            .O(N__40895),
            .I(\ALU.un9_addsub_cry_2_c_RNIA3LGZ0Z7 ));
    InMux I__9838 (
            .O(N__40892),
            .I(N__40889));
    LocalMux I__9837 (
            .O(N__40889),
            .I(N__40886));
    Span4Mux_h I__9836 (
            .O(N__40886),
            .I(N__40883));
    Span4Mux_h I__9835 (
            .O(N__40883),
            .I(N__40880));
    Odrv4 I__9834 (
            .O(N__40880),
            .I(\ALU.un2_addsub_cry_2_c_RNI5IV5FZ0 ));
    InMux I__9833 (
            .O(N__40877),
            .I(N__40874));
    LocalMux I__9832 (
            .O(N__40874),
            .I(N__40871));
    Span4Mux_v I__9831 (
            .O(N__40871),
            .I(N__40868));
    Span4Mux_h I__9830 (
            .O(N__40868),
            .I(N__40865));
    Odrv4 I__9829 (
            .O(N__40865),
            .I(\ALU.un2_addsub_cry_3_c_RNIOGGJGZ0 ));
    InMux I__9828 (
            .O(N__40862),
            .I(N__40859));
    LocalMux I__9827 (
            .O(N__40859),
            .I(N__40856));
    Odrv4 I__9826 (
            .O(N__40856),
            .I(\ALU.un9_addsub_cry_3_c_RNI525RZ0Z7 ));
    InMux I__9825 (
            .O(N__40853),
            .I(N__40850));
    LocalMux I__9824 (
            .O(N__40850),
            .I(N__40844));
    InMux I__9823 (
            .O(N__40849),
            .I(N__40841));
    InMux I__9822 (
            .O(N__40848),
            .I(N__40836));
    InMux I__9821 (
            .O(N__40847),
            .I(N__40836));
    Span4Mux_h I__9820 (
            .O(N__40844),
            .I(N__40833));
    LocalMux I__9819 (
            .O(N__40841),
            .I(N__40830));
    LocalMux I__9818 (
            .O(N__40836),
            .I(N__40827));
    Span4Mux_h I__9817 (
            .O(N__40833),
            .I(N__40823));
    Span4Mux_h I__9816 (
            .O(N__40830),
            .I(N__40820));
    Span4Mux_h I__9815 (
            .O(N__40827),
            .I(N__40817));
    InMux I__9814 (
            .O(N__40826),
            .I(N__40814));
    Odrv4 I__9813 (
            .O(N__40823),
            .I(\ALU.N_180_0 ));
    Odrv4 I__9812 (
            .O(N__40820),
            .I(\ALU.N_180_0 ));
    Odrv4 I__9811 (
            .O(N__40817),
            .I(\ALU.N_180_0 ));
    LocalMux I__9810 (
            .O(N__40814),
            .I(\ALU.N_180_0 ));
    CascadeMux I__9809 (
            .O(N__40805),
            .I(N__40802));
    InMux I__9808 (
            .O(N__40802),
            .I(N__40799));
    LocalMux I__9807 (
            .O(N__40799),
            .I(N__40796));
    Span4Mux_v I__9806 (
            .O(N__40796),
            .I(N__40793));
    Sp12to4 I__9805 (
            .O(N__40793),
            .I(N__40790));
    Odrv12 I__9804 (
            .O(N__40790),
            .I(\ALU.d_RNIFKNTEZ0Z_12 ));
    InMux I__9803 (
            .O(N__40787),
            .I(N__40784));
    LocalMux I__9802 (
            .O(N__40784),
            .I(N__40781));
    Span4Mux_h I__9801 (
            .O(N__40781),
            .I(N__40778));
    Odrv4 I__9800 (
            .O(N__40778),
            .I(\ALU.un9_addsub_cry_11_c_RNI10BQKZ0 ));
    InMux I__9799 (
            .O(N__40775),
            .I(\ALU.un9_addsub_cry_11 ));
    CascadeMux I__9798 (
            .O(N__40772),
            .I(N__40769));
    InMux I__9797 (
            .O(N__40769),
            .I(N__40760));
    InMux I__9796 (
            .O(N__40768),
            .I(N__40753));
    InMux I__9795 (
            .O(N__40767),
            .I(N__40753));
    InMux I__9794 (
            .O(N__40766),
            .I(N__40753));
    InMux I__9793 (
            .O(N__40765),
            .I(N__40748));
    CascadeMux I__9792 (
            .O(N__40764),
            .I(N__40743));
    InMux I__9791 (
            .O(N__40763),
            .I(N__40740));
    LocalMux I__9790 (
            .O(N__40760),
            .I(N__40737));
    LocalMux I__9789 (
            .O(N__40753),
            .I(N__40734));
    InMux I__9788 (
            .O(N__40752),
            .I(N__40729));
    InMux I__9787 (
            .O(N__40751),
            .I(N__40729));
    LocalMux I__9786 (
            .O(N__40748),
            .I(N__40726));
    InMux I__9785 (
            .O(N__40747),
            .I(N__40723));
    InMux I__9784 (
            .O(N__40746),
            .I(N__40718));
    InMux I__9783 (
            .O(N__40743),
            .I(N__40718));
    LocalMux I__9782 (
            .O(N__40740),
            .I(N__40715));
    Span4Mux_s3_h I__9781 (
            .O(N__40737),
            .I(N__40712));
    Span4Mux_v I__9780 (
            .O(N__40734),
            .I(N__40708));
    LocalMux I__9779 (
            .O(N__40729),
            .I(N__40701));
    Span4Mux_h I__9778 (
            .O(N__40726),
            .I(N__40701));
    LocalMux I__9777 (
            .O(N__40723),
            .I(N__40701));
    LocalMux I__9776 (
            .O(N__40718),
            .I(N__40696));
    Span4Mux_v I__9775 (
            .O(N__40715),
            .I(N__40696));
    Span4Mux_h I__9774 (
            .O(N__40712),
            .I(N__40693));
    InMux I__9773 (
            .O(N__40711),
            .I(N__40690));
    Span4Mux_h I__9772 (
            .O(N__40708),
            .I(N__40685));
    Span4Mux_v I__9771 (
            .O(N__40701),
            .I(N__40685));
    Span4Mux_h I__9770 (
            .O(N__40696),
            .I(N__40682));
    Span4Mux_h I__9769 (
            .O(N__40693),
            .I(N__40679));
    LocalMux I__9768 (
            .O(N__40690),
            .I(N__40674));
    Span4Mux_h I__9767 (
            .O(N__40685),
            .I(N__40674));
    Span4Mux_h I__9766 (
            .O(N__40682),
            .I(N__40671));
    Odrv4 I__9765 (
            .O(N__40679),
            .I(\ALU.aluOut_13 ));
    Odrv4 I__9764 (
            .O(N__40674),
            .I(\ALU.aluOut_13 ));
    Odrv4 I__9763 (
            .O(N__40671),
            .I(\ALU.aluOut_13 ));
    CascadeMux I__9762 (
            .O(N__40664),
            .I(N__40661));
    InMux I__9761 (
            .O(N__40661),
            .I(N__40658));
    LocalMux I__9760 (
            .O(N__40658),
            .I(N__40655));
    Span4Mux_v I__9759 (
            .O(N__40655),
            .I(N__40652));
    Odrv4 I__9758 (
            .O(N__40652),
            .I(\ALU.N_177_0_i ));
    InMux I__9757 (
            .O(N__40649),
            .I(N__40646));
    LocalMux I__9756 (
            .O(N__40646),
            .I(N__40643));
    Span4Mux_h I__9755 (
            .O(N__40643),
            .I(N__40640));
    Odrv4 I__9754 (
            .O(N__40640),
            .I(\ALU.un9_addsub_cry_12_c_RNIBB5QZ0Z9 ));
    InMux I__9753 (
            .O(N__40637),
            .I(\ALU.un9_addsub_cry_12 ));
    InMux I__9752 (
            .O(N__40634),
            .I(N__40631));
    LocalMux I__9751 (
            .O(N__40631),
            .I(N__40628));
    Span4Mux_h I__9750 (
            .O(N__40628),
            .I(N__40623));
    InMux I__9749 (
            .O(N__40627),
            .I(N__40620));
    InMux I__9748 (
            .O(N__40626),
            .I(N__40611));
    Span4Mux_v I__9747 (
            .O(N__40623),
            .I(N__40606));
    LocalMux I__9746 (
            .O(N__40620),
            .I(N__40606));
    InMux I__9745 (
            .O(N__40619),
            .I(N__40601));
    InMux I__9744 (
            .O(N__40618),
            .I(N__40601));
    InMux I__9743 (
            .O(N__40617),
            .I(N__40596));
    InMux I__9742 (
            .O(N__40616),
            .I(N__40593));
    InMux I__9741 (
            .O(N__40615),
            .I(N__40590));
    InMux I__9740 (
            .O(N__40614),
            .I(N__40587));
    LocalMux I__9739 (
            .O(N__40611),
            .I(N__40584));
    Span4Mux_h I__9738 (
            .O(N__40606),
            .I(N__40579));
    LocalMux I__9737 (
            .O(N__40601),
            .I(N__40579));
    InMux I__9736 (
            .O(N__40600),
            .I(N__40574));
    InMux I__9735 (
            .O(N__40599),
            .I(N__40574));
    LocalMux I__9734 (
            .O(N__40596),
            .I(\ALU.aluOut_14 ));
    LocalMux I__9733 (
            .O(N__40593),
            .I(\ALU.aluOut_14 ));
    LocalMux I__9732 (
            .O(N__40590),
            .I(\ALU.aluOut_14 ));
    LocalMux I__9731 (
            .O(N__40587),
            .I(\ALU.aluOut_14 ));
    Odrv4 I__9730 (
            .O(N__40584),
            .I(\ALU.aluOut_14 ));
    Odrv4 I__9729 (
            .O(N__40579),
            .I(\ALU.aluOut_14 ));
    LocalMux I__9728 (
            .O(N__40574),
            .I(\ALU.aluOut_14 ));
    CascadeMux I__9727 (
            .O(N__40559),
            .I(N__40556));
    InMux I__9726 (
            .O(N__40556),
            .I(N__40553));
    LocalMux I__9725 (
            .O(N__40553),
            .I(N__40550));
    Span4Mux_v I__9724 (
            .O(N__40550),
            .I(N__40547));
    Span4Mux_h I__9723 (
            .O(N__40547),
            .I(N__40544));
    Span4Mux_h I__9722 (
            .O(N__40544),
            .I(N__40541));
    Odrv4 I__9721 (
            .O(N__40541),
            .I(\ALU.N_171_0_i ));
    InMux I__9720 (
            .O(N__40538),
            .I(N__40535));
    LocalMux I__9719 (
            .O(N__40535),
            .I(N__40532));
    Span4Mux_h I__9718 (
            .O(N__40532),
            .I(N__40529));
    Odrv4 I__9717 (
            .O(N__40529),
            .I(\ALU.un9_addsub_cry_13_c_RNI4JGFZ0Z9 ));
    InMux I__9716 (
            .O(N__40526),
            .I(\ALU.un9_addsub_cry_13 ));
    InMux I__9715 (
            .O(N__40523),
            .I(N__40520));
    LocalMux I__9714 (
            .O(N__40520),
            .I(N__40517));
    Span4Mux_v I__9713 (
            .O(N__40517),
            .I(N__40514));
    Sp12to4 I__9712 (
            .O(N__40514),
            .I(N__40511));
    Odrv12 I__9711 (
            .O(N__40511),
            .I(\ALU.un9_addsub_axb_15 ));
    CascadeMux I__9710 (
            .O(N__40508),
            .I(N__40505));
    InMux I__9709 (
            .O(N__40505),
            .I(N__40502));
    LocalMux I__9708 (
            .O(N__40502),
            .I(N__40499));
    Span4Mux_v I__9707 (
            .O(N__40499),
            .I(N__40496));
    Sp12to4 I__9706 (
            .O(N__40496),
            .I(N__40493));
    Odrv12 I__9705 (
            .O(N__40493),
            .I(\ALU.un2_addsub_cry_14_c_RNINOKZ0Z69 ));
    InMux I__9704 (
            .O(N__40490),
            .I(\ALU.un9_addsub_cry_14 ));
    InMux I__9703 (
            .O(N__40487),
            .I(N__40484));
    LocalMux I__9702 (
            .O(N__40484),
            .I(\ALU.un9_addsub_cry_14_c_RNIS374JZ0 ));
    InMux I__9701 (
            .O(N__40481),
            .I(N__40478));
    LocalMux I__9700 (
            .O(N__40478),
            .I(N__40475));
    Span4Mux_v I__9699 (
            .O(N__40475),
            .I(N__40472));
    Span4Mux_h I__9698 (
            .O(N__40472),
            .I(N__40469));
    Odrv4 I__9697 (
            .O(N__40469),
            .I(\ALU.c_RNIA9V4LZ0Z_15 ));
    InMux I__9696 (
            .O(N__40466),
            .I(N__40463));
    LocalMux I__9695 (
            .O(N__40463),
            .I(N__40460));
    Span12Mux_v I__9694 (
            .O(N__40460),
            .I(N__40457));
    Odrv12 I__9693 (
            .O(N__40457),
            .I(\ALU.d_RNI9DPVUZ0Z_6 ));
    CascadeMux I__9692 (
            .O(N__40454),
            .I(\ALU.rshift_3_cascade_ ));
    InMux I__9691 (
            .O(N__40451),
            .I(N__40448));
    LocalMux I__9690 (
            .O(N__40448),
            .I(N__40445));
    Span12Mux_s9_v I__9689 (
            .O(N__40445),
            .I(N__40442));
    Span12Mux_h I__9688 (
            .O(N__40442),
            .I(N__40439));
    Odrv12 I__9687 (
            .O(N__40439),
            .I(\ALU.N_293_0 ));
    CascadeMux I__9686 (
            .O(N__40436),
            .I(\ALU.d_RNI3V2CP1Z0Z_3_cascade_ ));
    CascadeMux I__9685 (
            .O(N__40433),
            .I(N__40420));
    InMux I__9684 (
            .O(N__40432),
            .I(N__40414));
    InMux I__9683 (
            .O(N__40431),
            .I(N__40414));
    InMux I__9682 (
            .O(N__40430),
            .I(N__40411));
    InMux I__9681 (
            .O(N__40429),
            .I(N__40406));
    InMux I__9680 (
            .O(N__40428),
            .I(N__40403));
    InMux I__9679 (
            .O(N__40427),
            .I(N__40398));
    InMux I__9678 (
            .O(N__40426),
            .I(N__40395));
    InMux I__9677 (
            .O(N__40425),
            .I(N__40392));
    InMux I__9676 (
            .O(N__40424),
            .I(N__40385));
    InMux I__9675 (
            .O(N__40423),
            .I(N__40380));
    InMux I__9674 (
            .O(N__40420),
            .I(N__40380));
    InMux I__9673 (
            .O(N__40419),
            .I(N__40377));
    LocalMux I__9672 (
            .O(N__40414),
            .I(N__40372));
    LocalMux I__9671 (
            .O(N__40411),
            .I(N__40372));
    InMux I__9670 (
            .O(N__40410),
            .I(N__40369));
    CascadeMux I__9669 (
            .O(N__40409),
            .I(N__40363));
    LocalMux I__9668 (
            .O(N__40406),
            .I(N__40357));
    LocalMux I__9667 (
            .O(N__40403),
            .I(N__40357));
    InMux I__9666 (
            .O(N__40402),
            .I(N__40354));
    InMux I__9665 (
            .O(N__40401),
            .I(N__40351));
    LocalMux I__9664 (
            .O(N__40398),
            .I(N__40348));
    LocalMux I__9663 (
            .O(N__40395),
            .I(N__40343));
    LocalMux I__9662 (
            .O(N__40392),
            .I(N__40343));
    InMux I__9661 (
            .O(N__40391),
            .I(N__40340));
    InMux I__9660 (
            .O(N__40390),
            .I(N__40337));
    InMux I__9659 (
            .O(N__40389),
            .I(N__40332));
    InMux I__9658 (
            .O(N__40388),
            .I(N__40332));
    LocalMux I__9657 (
            .O(N__40385),
            .I(N__40329));
    LocalMux I__9656 (
            .O(N__40380),
            .I(N__40326));
    LocalMux I__9655 (
            .O(N__40377),
            .I(N__40319));
    Span4Mux_v I__9654 (
            .O(N__40372),
            .I(N__40319));
    LocalMux I__9653 (
            .O(N__40369),
            .I(N__40319));
    InMux I__9652 (
            .O(N__40368),
            .I(N__40316));
    InMux I__9651 (
            .O(N__40367),
            .I(N__40311));
    InMux I__9650 (
            .O(N__40366),
            .I(N__40311));
    InMux I__9649 (
            .O(N__40363),
            .I(N__40306));
    InMux I__9648 (
            .O(N__40362),
            .I(N__40306));
    Span12Mux_h I__9647 (
            .O(N__40357),
            .I(N__40301));
    LocalMux I__9646 (
            .O(N__40354),
            .I(N__40301));
    LocalMux I__9645 (
            .O(N__40351),
            .I(N__40298));
    Span4Mux_v I__9644 (
            .O(N__40348),
            .I(N__40293));
    Span4Mux_v I__9643 (
            .O(N__40343),
            .I(N__40293));
    LocalMux I__9642 (
            .O(N__40340),
            .I(N__40288));
    LocalMux I__9641 (
            .O(N__40337),
            .I(N__40283));
    LocalMux I__9640 (
            .O(N__40332),
            .I(N__40283));
    Span4Mux_v I__9639 (
            .O(N__40329),
            .I(N__40278));
    Span4Mux_h I__9638 (
            .O(N__40326),
            .I(N__40278));
    Span4Mux_v I__9637 (
            .O(N__40319),
            .I(N__40271));
    LocalMux I__9636 (
            .O(N__40316),
            .I(N__40271));
    LocalMux I__9635 (
            .O(N__40311),
            .I(N__40266));
    LocalMux I__9634 (
            .O(N__40306),
            .I(N__40266));
    Span12Mux_v I__9633 (
            .O(N__40301),
            .I(N__40263));
    Span12Mux_v I__9632 (
            .O(N__40298),
            .I(N__40258));
    Sp12to4 I__9631 (
            .O(N__40293),
            .I(N__40258));
    InMux I__9630 (
            .O(N__40292),
            .I(N__40253));
    InMux I__9629 (
            .O(N__40291),
            .I(N__40253));
    Span12Mux_h I__9628 (
            .O(N__40288),
            .I(N__40246));
    Span12Mux_s5_h I__9627 (
            .O(N__40283),
            .I(N__40246));
    Sp12to4 I__9626 (
            .O(N__40278),
            .I(N__40246));
    InMux I__9625 (
            .O(N__40277),
            .I(N__40241));
    InMux I__9624 (
            .O(N__40276),
            .I(N__40241));
    Span4Mux_v I__9623 (
            .O(N__40271),
            .I(N__40236));
    Span4Mux_v I__9622 (
            .O(N__40266),
            .I(N__40236));
    Odrv12 I__9621 (
            .O(N__40263),
            .I(\ALU.aluOut_5 ));
    Odrv12 I__9620 (
            .O(N__40258),
            .I(\ALU.aluOut_5 ));
    LocalMux I__9619 (
            .O(N__40253),
            .I(\ALU.aluOut_5 ));
    Odrv12 I__9618 (
            .O(N__40246),
            .I(\ALU.aluOut_5 ));
    LocalMux I__9617 (
            .O(N__40241),
            .I(\ALU.aluOut_5 ));
    Odrv4 I__9616 (
            .O(N__40236),
            .I(\ALU.aluOut_5 ));
    CascadeMux I__9615 (
            .O(N__40223),
            .I(N__40220));
    InMux I__9614 (
            .O(N__40220),
            .I(N__40217));
    LocalMux I__9613 (
            .O(N__40217),
            .I(N__40214));
    Span4Mux_h I__9612 (
            .O(N__40214),
            .I(N__40211));
    Span4Mux_v I__9611 (
            .O(N__40211),
            .I(N__40208));
    Span4Mux_v I__9610 (
            .O(N__40208),
            .I(N__40205));
    Span4Mux_h I__9609 (
            .O(N__40205),
            .I(N__40202));
    Span4Mux_h I__9608 (
            .O(N__40202),
            .I(N__40199));
    Odrv4 I__9607 (
            .O(N__40199),
            .I(\ALU.N_225_0_i ));
    InMux I__9606 (
            .O(N__40196),
            .I(\ALU.un9_addsub_cry_4 ));
    CascadeMux I__9605 (
            .O(N__40193),
            .I(N__40190));
    InMux I__9604 (
            .O(N__40190),
            .I(N__40187));
    LocalMux I__9603 (
            .O(N__40187),
            .I(N__40184));
    Span4Mux_h I__9602 (
            .O(N__40184),
            .I(N__40181));
    Span4Mux_h I__9601 (
            .O(N__40181),
            .I(N__40178));
    Odrv4 I__9600 (
            .O(N__40178),
            .I(\ALU.N_219_0_i ));
    InMux I__9599 (
            .O(N__40175),
            .I(\ALU.un9_addsub_cry_5 ));
    CascadeMux I__9598 (
            .O(N__40172),
            .I(N__40169));
    InMux I__9597 (
            .O(N__40169),
            .I(N__40166));
    LocalMux I__9596 (
            .O(N__40166),
            .I(N__40163));
    Span4Mux_h I__9595 (
            .O(N__40163),
            .I(N__40160));
    Span4Mux_v I__9594 (
            .O(N__40160),
            .I(N__40157));
    Span4Mux_v I__9593 (
            .O(N__40157),
            .I(N__40154));
    Span4Mux_h I__9592 (
            .O(N__40154),
            .I(N__40151));
    Span4Mux_h I__9591 (
            .O(N__40151),
            .I(N__40148));
    Odrv4 I__9590 (
            .O(N__40148),
            .I(\ALU.N_213_0_i ));
    InMux I__9589 (
            .O(N__40145),
            .I(N__40142));
    LocalMux I__9588 (
            .O(N__40142),
            .I(N__40139));
    Span4Mux_h I__9587 (
            .O(N__40139),
            .I(N__40136));
    Span4Mux_h I__9586 (
            .O(N__40136),
            .I(N__40133));
    Span4Mux_v I__9585 (
            .O(N__40133),
            .I(N__40130));
    Span4Mux_v I__9584 (
            .O(N__40130),
            .I(N__40127));
    Odrv4 I__9583 (
            .O(N__40127),
            .I(\ALU.un9_addsub_cry_6_c_RNI2EFHZ0Z8 ));
    InMux I__9582 (
            .O(N__40124),
            .I(\ALU.un9_addsub_cry_6 ));
    InMux I__9581 (
            .O(N__40121),
            .I(N__40116));
    CascadeMux I__9580 (
            .O(N__40120),
            .I(N__40113));
    InMux I__9579 (
            .O(N__40119),
            .I(N__40108));
    LocalMux I__9578 (
            .O(N__40116),
            .I(N__40104));
    InMux I__9577 (
            .O(N__40113),
            .I(N__40099));
    CascadeMux I__9576 (
            .O(N__40112),
            .I(N__40095));
    InMux I__9575 (
            .O(N__40111),
            .I(N__40090));
    LocalMux I__9574 (
            .O(N__40108),
            .I(N__40087));
    CascadeMux I__9573 (
            .O(N__40107),
            .I(N__40076));
    Span4Mux_v I__9572 (
            .O(N__40104),
            .I(N__40072));
    InMux I__9571 (
            .O(N__40103),
            .I(N__40066));
    InMux I__9570 (
            .O(N__40102),
            .I(N__40063));
    LocalMux I__9569 (
            .O(N__40099),
            .I(N__40060));
    InMux I__9568 (
            .O(N__40098),
            .I(N__40057));
    InMux I__9567 (
            .O(N__40095),
            .I(N__40053));
    InMux I__9566 (
            .O(N__40094),
            .I(N__40050));
    InMux I__9565 (
            .O(N__40093),
            .I(N__40047));
    LocalMux I__9564 (
            .O(N__40090),
            .I(N__40040));
    Span4Mux_v I__9563 (
            .O(N__40087),
            .I(N__40037));
    InMux I__9562 (
            .O(N__40086),
            .I(N__40032));
    InMux I__9561 (
            .O(N__40085),
            .I(N__40032));
    InMux I__9560 (
            .O(N__40084),
            .I(N__40029));
    InMux I__9559 (
            .O(N__40083),
            .I(N__40022));
    InMux I__9558 (
            .O(N__40082),
            .I(N__40022));
    InMux I__9557 (
            .O(N__40081),
            .I(N__40022));
    InMux I__9556 (
            .O(N__40080),
            .I(N__40015));
    InMux I__9555 (
            .O(N__40079),
            .I(N__40015));
    InMux I__9554 (
            .O(N__40076),
            .I(N__40015));
    InMux I__9553 (
            .O(N__40075),
            .I(N__40012));
    Span4Mux_h I__9552 (
            .O(N__40072),
            .I(N__40009));
    InMux I__9551 (
            .O(N__40071),
            .I(N__40006));
    InMux I__9550 (
            .O(N__40070),
            .I(N__40001));
    InMux I__9549 (
            .O(N__40069),
            .I(N__40001));
    LocalMux I__9548 (
            .O(N__40066),
            .I(N__39996));
    LocalMux I__9547 (
            .O(N__40063),
            .I(N__39996));
    Span4Mux_v I__9546 (
            .O(N__40060),
            .I(N__39993));
    LocalMux I__9545 (
            .O(N__40057),
            .I(N__39990));
    InMux I__9544 (
            .O(N__40056),
            .I(N__39987));
    LocalMux I__9543 (
            .O(N__40053),
            .I(N__39984));
    LocalMux I__9542 (
            .O(N__40050),
            .I(N__39979));
    LocalMux I__9541 (
            .O(N__40047),
            .I(N__39979));
    InMux I__9540 (
            .O(N__40046),
            .I(N__39976));
    InMux I__9539 (
            .O(N__40045),
            .I(N__39971));
    InMux I__9538 (
            .O(N__40044),
            .I(N__39971));
    InMux I__9537 (
            .O(N__40043),
            .I(N__39968));
    Span4Mux_v I__9536 (
            .O(N__40040),
            .I(N__39963));
    Span4Mux_h I__9535 (
            .O(N__40037),
            .I(N__39963));
    LocalMux I__9534 (
            .O(N__40032),
            .I(N__39960));
    LocalMux I__9533 (
            .O(N__40029),
            .I(N__39953));
    LocalMux I__9532 (
            .O(N__40022),
            .I(N__39953));
    LocalMux I__9531 (
            .O(N__40015),
            .I(N__39953));
    LocalMux I__9530 (
            .O(N__40012),
            .I(N__39950));
    Span4Mux_h I__9529 (
            .O(N__40009),
            .I(N__39943));
    LocalMux I__9528 (
            .O(N__40006),
            .I(N__39943));
    LocalMux I__9527 (
            .O(N__40001),
            .I(N__39943));
    Span4Mux_v I__9526 (
            .O(N__39996),
            .I(N__39940));
    Span4Mux_h I__9525 (
            .O(N__39993),
            .I(N__39933));
    Span4Mux_v I__9524 (
            .O(N__39990),
            .I(N__39933));
    LocalMux I__9523 (
            .O(N__39987),
            .I(N__39933));
    Span4Mux_s1_h I__9522 (
            .O(N__39984),
            .I(N__39928));
    Span4Mux_v I__9521 (
            .O(N__39979),
            .I(N__39928));
    LocalMux I__9520 (
            .O(N__39976),
            .I(N__39923));
    LocalMux I__9519 (
            .O(N__39971),
            .I(N__39923));
    LocalMux I__9518 (
            .O(N__39968),
            .I(N__39920));
    Span4Mux_v I__9517 (
            .O(N__39963),
            .I(N__39913));
    Span4Mux_v I__9516 (
            .O(N__39960),
            .I(N__39913));
    Span4Mux_v I__9515 (
            .O(N__39953),
            .I(N__39913));
    Span4Mux_v I__9514 (
            .O(N__39950),
            .I(N__39904));
    Span4Mux_v I__9513 (
            .O(N__39943),
            .I(N__39904));
    Span4Mux_h I__9512 (
            .O(N__39940),
            .I(N__39904));
    Span4Mux_v I__9511 (
            .O(N__39933),
            .I(N__39904));
    Span4Mux_h I__9510 (
            .O(N__39928),
            .I(N__39899));
    Span4Mux_v I__9509 (
            .O(N__39923),
            .I(N__39899));
    Odrv4 I__9508 (
            .O(N__39920),
            .I(\ALU.aluOut_8 ));
    Odrv4 I__9507 (
            .O(N__39913),
            .I(\ALU.aluOut_8 ));
    Odrv4 I__9506 (
            .O(N__39904),
            .I(\ALU.aluOut_8 ));
    Odrv4 I__9505 (
            .O(N__39899),
            .I(\ALU.aluOut_8 ));
    CascadeMux I__9504 (
            .O(N__39890),
            .I(N__39887));
    InMux I__9503 (
            .O(N__39887),
            .I(N__39884));
    LocalMux I__9502 (
            .O(N__39884),
            .I(N__39881));
    Span12Mux_h I__9501 (
            .O(N__39881),
            .I(N__39878));
    Odrv12 I__9500 (
            .O(N__39878),
            .I(\ALU.N_201_0_i ));
    InMux I__9499 (
            .O(N__39875),
            .I(N__39872));
    LocalMux I__9498 (
            .O(N__39872),
            .I(N__39869));
    Span4Mux_v I__9497 (
            .O(N__39869),
            .I(N__39866));
    Odrv4 I__9496 (
            .O(N__39866),
            .I(\ALU.un9_addsub_cry_7_c_RNIU7FZ0Z18 ));
    InMux I__9495 (
            .O(N__39863),
            .I(bfn_13_8_0_));
    InMux I__9494 (
            .O(N__39860),
            .I(N__39856));
    InMux I__9493 (
            .O(N__39859),
            .I(N__39844));
    LocalMux I__9492 (
            .O(N__39856),
            .I(N__39841));
    InMux I__9491 (
            .O(N__39855),
            .I(N__39838));
    CascadeMux I__9490 (
            .O(N__39854),
            .I(N__39833));
    InMux I__9489 (
            .O(N__39853),
            .I(N__39829));
    CascadeMux I__9488 (
            .O(N__39852),
            .I(N__39826));
    InMux I__9487 (
            .O(N__39851),
            .I(N__39822));
    InMux I__9486 (
            .O(N__39850),
            .I(N__39818));
    InMux I__9485 (
            .O(N__39849),
            .I(N__39815));
    InMux I__9484 (
            .O(N__39848),
            .I(N__39809));
    InMux I__9483 (
            .O(N__39847),
            .I(N__39809));
    LocalMux I__9482 (
            .O(N__39844),
            .I(N__39804));
    Span4Mux_h I__9481 (
            .O(N__39841),
            .I(N__39799));
    LocalMux I__9480 (
            .O(N__39838),
            .I(N__39799));
    CascadeMux I__9479 (
            .O(N__39837),
            .I(N__39796));
    InMux I__9478 (
            .O(N__39836),
            .I(N__39792));
    InMux I__9477 (
            .O(N__39833),
            .I(N__39789));
    InMux I__9476 (
            .O(N__39832),
            .I(N__39786));
    LocalMux I__9475 (
            .O(N__39829),
            .I(N__39783));
    InMux I__9474 (
            .O(N__39826),
            .I(N__39780));
    InMux I__9473 (
            .O(N__39825),
            .I(N__39777));
    LocalMux I__9472 (
            .O(N__39822),
            .I(N__39774));
    InMux I__9471 (
            .O(N__39821),
            .I(N__39771));
    LocalMux I__9470 (
            .O(N__39818),
            .I(N__39768));
    LocalMux I__9469 (
            .O(N__39815),
            .I(N__39765));
    InMux I__9468 (
            .O(N__39814),
            .I(N__39762));
    LocalMux I__9467 (
            .O(N__39809),
            .I(N__39759));
    InMux I__9466 (
            .O(N__39808),
            .I(N__39756));
    InMux I__9465 (
            .O(N__39807),
            .I(N__39753));
    Span4Mux_h I__9464 (
            .O(N__39804),
            .I(N__39748));
    Span4Mux_h I__9463 (
            .O(N__39799),
            .I(N__39745));
    InMux I__9462 (
            .O(N__39796),
            .I(N__39740));
    InMux I__9461 (
            .O(N__39795),
            .I(N__39740));
    LocalMux I__9460 (
            .O(N__39792),
            .I(N__39737));
    LocalMux I__9459 (
            .O(N__39789),
            .I(N__39734));
    LocalMux I__9458 (
            .O(N__39786),
            .I(N__39731));
    Span4Mux_v I__9457 (
            .O(N__39783),
            .I(N__39728));
    LocalMux I__9456 (
            .O(N__39780),
            .I(N__39725));
    LocalMux I__9455 (
            .O(N__39777),
            .I(N__39722));
    Span4Mux_v I__9454 (
            .O(N__39774),
            .I(N__39717));
    LocalMux I__9453 (
            .O(N__39771),
            .I(N__39717));
    Span4Mux_v I__9452 (
            .O(N__39768),
            .I(N__39712));
    Span4Mux_v I__9451 (
            .O(N__39765),
            .I(N__39712));
    LocalMux I__9450 (
            .O(N__39762),
            .I(N__39709));
    Span4Mux_v I__9449 (
            .O(N__39759),
            .I(N__39704));
    LocalMux I__9448 (
            .O(N__39756),
            .I(N__39704));
    LocalMux I__9447 (
            .O(N__39753),
            .I(N__39701));
    InMux I__9446 (
            .O(N__39752),
            .I(N__39698));
    InMux I__9445 (
            .O(N__39751),
            .I(N__39695));
    Span4Mux_h I__9444 (
            .O(N__39748),
            .I(N__39692));
    Span4Mux_v I__9443 (
            .O(N__39745),
            .I(N__39689));
    LocalMux I__9442 (
            .O(N__39740),
            .I(N__39686));
    Span4Mux_v I__9441 (
            .O(N__39737),
            .I(N__39681));
    Span4Mux_h I__9440 (
            .O(N__39734),
            .I(N__39681));
    Span4Mux_v I__9439 (
            .O(N__39731),
            .I(N__39676));
    Span4Mux_h I__9438 (
            .O(N__39728),
            .I(N__39676));
    Span4Mux_v I__9437 (
            .O(N__39725),
            .I(N__39665));
    Span4Mux_v I__9436 (
            .O(N__39722),
            .I(N__39665));
    Span4Mux_v I__9435 (
            .O(N__39717),
            .I(N__39665));
    Span4Mux_h I__9434 (
            .O(N__39712),
            .I(N__39665));
    Span4Mux_h I__9433 (
            .O(N__39709),
            .I(N__39665));
    Span4Mux_v I__9432 (
            .O(N__39704),
            .I(N__39656));
    Span4Mux_s3_h I__9431 (
            .O(N__39701),
            .I(N__39656));
    LocalMux I__9430 (
            .O(N__39698),
            .I(N__39656));
    LocalMux I__9429 (
            .O(N__39695),
            .I(N__39656));
    Odrv4 I__9428 (
            .O(N__39692),
            .I(\ALU.aluOut_9 ));
    Odrv4 I__9427 (
            .O(N__39689),
            .I(\ALU.aluOut_9 ));
    Odrv12 I__9426 (
            .O(N__39686),
            .I(\ALU.aluOut_9 ));
    Odrv4 I__9425 (
            .O(N__39681),
            .I(\ALU.aluOut_9 ));
    Odrv4 I__9424 (
            .O(N__39676),
            .I(\ALU.aluOut_9 ));
    Odrv4 I__9423 (
            .O(N__39665),
            .I(\ALU.aluOut_9 ));
    Odrv4 I__9422 (
            .O(N__39656),
            .I(\ALU.aluOut_9 ));
    CascadeMux I__9421 (
            .O(N__39641),
            .I(N__39638));
    InMux I__9420 (
            .O(N__39638),
            .I(N__39635));
    LocalMux I__9419 (
            .O(N__39635),
            .I(N__39632));
    Span4Mux_v I__9418 (
            .O(N__39632),
            .I(N__39629));
    Sp12to4 I__9417 (
            .O(N__39629),
            .I(N__39626));
    Odrv12 I__9416 (
            .O(N__39626),
            .I(\ALU.N_207_0_i ));
    InMux I__9415 (
            .O(N__39623),
            .I(N__39620));
    LocalMux I__9414 (
            .O(N__39620),
            .I(N__39617));
    Span4Mux_v I__9413 (
            .O(N__39617),
            .I(N__39614));
    Odrv4 I__9412 (
            .O(N__39614),
            .I(\ALU.un9_addsub_cry_8_c_RNIPV1SZ0Z8 ));
    InMux I__9411 (
            .O(N__39611),
            .I(\ALU.un9_addsub_cry_8 ));
    CascadeMux I__9410 (
            .O(N__39608),
            .I(N__39602));
    CascadeMux I__9409 (
            .O(N__39607),
            .I(N__39596));
    CascadeMux I__9408 (
            .O(N__39606),
            .I(N__39590));
    InMux I__9407 (
            .O(N__39605),
            .I(N__39587));
    InMux I__9406 (
            .O(N__39602),
            .I(N__39579));
    InMux I__9405 (
            .O(N__39601),
            .I(N__39579));
    InMux I__9404 (
            .O(N__39600),
            .I(N__39579));
    InMux I__9403 (
            .O(N__39599),
            .I(N__39572));
    InMux I__9402 (
            .O(N__39596),
            .I(N__39572));
    InMux I__9401 (
            .O(N__39595),
            .I(N__39572));
    InMux I__9400 (
            .O(N__39594),
            .I(N__39566));
    InMux I__9399 (
            .O(N__39593),
            .I(N__39566));
    InMux I__9398 (
            .O(N__39590),
            .I(N__39563));
    LocalMux I__9397 (
            .O(N__39587),
            .I(N__39560));
    InMux I__9396 (
            .O(N__39586),
            .I(N__39557));
    LocalMux I__9395 (
            .O(N__39579),
            .I(N__39554));
    LocalMux I__9394 (
            .O(N__39572),
            .I(N__39551));
    InMux I__9393 (
            .O(N__39571),
            .I(N__39548));
    LocalMux I__9392 (
            .O(N__39566),
            .I(N__39545));
    LocalMux I__9391 (
            .O(N__39563),
            .I(N__39540));
    Span4Mux_h I__9390 (
            .O(N__39560),
            .I(N__39540));
    LocalMux I__9389 (
            .O(N__39557),
            .I(N__39537));
    Span4Mux_v I__9388 (
            .O(N__39554),
            .I(N__39532));
    Span4Mux_s1_h I__9387 (
            .O(N__39551),
            .I(N__39532));
    LocalMux I__9386 (
            .O(N__39548),
            .I(N__39528));
    Span4Mux_h I__9385 (
            .O(N__39545),
            .I(N__39525));
    Span4Mux_h I__9384 (
            .O(N__39540),
            .I(N__39518));
    Span4Mux_v I__9383 (
            .O(N__39537),
            .I(N__39518));
    Span4Mux_h I__9382 (
            .O(N__39532),
            .I(N__39518));
    InMux I__9381 (
            .O(N__39531),
            .I(N__39515));
    Odrv12 I__9380 (
            .O(N__39528),
            .I(\ALU.N_192_0 ));
    Odrv4 I__9379 (
            .O(N__39525),
            .I(\ALU.N_192_0 ));
    Odrv4 I__9378 (
            .O(N__39518),
            .I(\ALU.N_192_0 ));
    LocalMux I__9377 (
            .O(N__39515),
            .I(\ALU.N_192_0 ));
    CascadeMux I__9376 (
            .O(N__39506),
            .I(N__39503));
    InMux I__9375 (
            .O(N__39503),
            .I(N__39500));
    LocalMux I__9374 (
            .O(N__39500),
            .I(N__39497));
    Sp12to4 I__9373 (
            .O(N__39497),
            .I(N__39494));
    Span12Mux_h I__9372 (
            .O(N__39494),
            .I(N__39491));
    Odrv12 I__9371 (
            .O(N__39491),
            .I(\ALU.a_RNIV2S0FZ0Z_10 ));
    InMux I__9370 (
            .O(N__39488),
            .I(N__39485));
    LocalMux I__9369 (
            .O(N__39485),
            .I(N__39482));
    Odrv12 I__9368 (
            .O(N__39482),
            .I(\ALU.un9_addsub_cry_9_c_RNI22U6KZ0 ));
    InMux I__9367 (
            .O(N__39479),
            .I(\ALU.un9_addsub_cry_9 ));
    InMux I__9366 (
            .O(N__39476),
            .I(N__39473));
    LocalMux I__9365 (
            .O(N__39473),
            .I(N__39468));
    InMux I__9364 (
            .O(N__39472),
            .I(N__39464));
    InMux I__9363 (
            .O(N__39471),
            .I(N__39460));
    Span4Mux_v I__9362 (
            .O(N__39468),
            .I(N__39457));
    InMux I__9361 (
            .O(N__39467),
            .I(N__39454));
    LocalMux I__9360 (
            .O(N__39464),
            .I(N__39449));
    InMux I__9359 (
            .O(N__39463),
            .I(N__39444));
    LocalMux I__9358 (
            .O(N__39460),
            .I(N__39441));
    Sp12to4 I__9357 (
            .O(N__39457),
            .I(N__39435));
    LocalMux I__9356 (
            .O(N__39454),
            .I(N__39435));
    InMux I__9355 (
            .O(N__39453),
            .I(N__39430));
    InMux I__9354 (
            .O(N__39452),
            .I(N__39430));
    Span4Mux_v I__9353 (
            .O(N__39449),
            .I(N__39427));
    InMux I__9352 (
            .O(N__39448),
            .I(N__39422));
    InMux I__9351 (
            .O(N__39447),
            .I(N__39422));
    LocalMux I__9350 (
            .O(N__39444),
            .I(N__39419));
    Span4Mux_v I__9349 (
            .O(N__39441),
            .I(N__39416));
    InMux I__9348 (
            .O(N__39440),
            .I(N__39413));
    Odrv12 I__9347 (
            .O(N__39435),
            .I(\ALU.N_186_0 ));
    LocalMux I__9346 (
            .O(N__39430),
            .I(\ALU.N_186_0 ));
    Odrv4 I__9345 (
            .O(N__39427),
            .I(\ALU.N_186_0 ));
    LocalMux I__9344 (
            .O(N__39422),
            .I(\ALU.N_186_0 ));
    Odrv4 I__9343 (
            .O(N__39419),
            .I(\ALU.N_186_0 ));
    Odrv4 I__9342 (
            .O(N__39416),
            .I(\ALU.N_186_0 ));
    LocalMux I__9341 (
            .O(N__39413),
            .I(\ALU.N_186_0 ));
    CascadeMux I__9340 (
            .O(N__39398),
            .I(N__39391));
    InMux I__9339 (
            .O(N__39397),
            .I(N__39379));
    CascadeMux I__9338 (
            .O(N__39396),
            .I(N__39376));
    InMux I__9337 (
            .O(N__39395),
            .I(N__39372));
    InMux I__9336 (
            .O(N__39394),
            .I(N__39369));
    InMux I__9335 (
            .O(N__39391),
            .I(N__39365));
    InMux I__9334 (
            .O(N__39390),
            .I(N__39362));
    InMux I__9333 (
            .O(N__39389),
            .I(N__39359));
    InMux I__9332 (
            .O(N__39388),
            .I(N__39356));
    InMux I__9331 (
            .O(N__39387),
            .I(N__39351));
    InMux I__9330 (
            .O(N__39386),
            .I(N__39351));
    InMux I__9329 (
            .O(N__39385),
            .I(N__39348));
    InMux I__9328 (
            .O(N__39384),
            .I(N__39345));
    CascadeMux I__9327 (
            .O(N__39383),
            .I(N__39342));
    InMux I__9326 (
            .O(N__39382),
            .I(N__39338));
    LocalMux I__9325 (
            .O(N__39379),
            .I(N__39335));
    InMux I__9324 (
            .O(N__39376),
            .I(N__39331));
    InMux I__9323 (
            .O(N__39375),
            .I(N__39328));
    LocalMux I__9322 (
            .O(N__39372),
            .I(N__39323));
    LocalMux I__9321 (
            .O(N__39369),
            .I(N__39323));
    InMux I__9320 (
            .O(N__39368),
            .I(N__39319));
    LocalMux I__9319 (
            .O(N__39365),
            .I(N__39316));
    LocalMux I__9318 (
            .O(N__39362),
            .I(N__39313));
    LocalMux I__9317 (
            .O(N__39359),
            .I(N__39308));
    LocalMux I__9316 (
            .O(N__39356),
            .I(N__39308));
    LocalMux I__9315 (
            .O(N__39351),
            .I(N__39301));
    LocalMux I__9314 (
            .O(N__39348),
            .I(N__39301));
    LocalMux I__9313 (
            .O(N__39345),
            .I(N__39301));
    InMux I__9312 (
            .O(N__39342),
            .I(N__39296));
    InMux I__9311 (
            .O(N__39341),
            .I(N__39296));
    LocalMux I__9310 (
            .O(N__39338),
            .I(N__39293));
    Span4Mux_v I__9309 (
            .O(N__39335),
            .I(N__39290));
    InMux I__9308 (
            .O(N__39334),
            .I(N__39287));
    LocalMux I__9307 (
            .O(N__39331),
            .I(N__39279));
    LocalMux I__9306 (
            .O(N__39328),
            .I(N__39279));
    Span4Mux_v I__9305 (
            .O(N__39323),
            .I(N__39279));
    InMux I__9304 (
            .O(N__39322),
            .I(N__39276));
    LocalMux I__9303 (
            .O(N__39319),
            .I(N__39273));
    Span4Mux_v I__9302 (
            .O(N__39316),
            .I(N__39270));
    Span4Mux_v I__9301 (
            .O(N__39313),
            .I(N__39267));
    Span4Mux_h I__9300 (
            .O(N__39308),
            .I(N__39260));
    Span4Mux_v I__9299 (
            .O(N__39301),
            .I(N__39260));
    LocalMux I__9298 (
            .O(N__39296),
            .I(N__39260));
    Span4Mux_v I__9297 (
            .O(N__39293),
            .I(N__39253));
    Span4Mux_h I__9296 (
            .O(N__39290),
            .I(N__39253));
    LocalMux I__9295 (
            .O(N__39287),
            .I(N__39253));
    InMux I__9294 (
            .O(N__39286),
            .I(N__39250));
    Span4Mux_v I__9293 (
            .O(N__39279),
            .I(N__39247));
    LocalMux I__9292 (
            .O(N__39276),
            .I(N__39244));
    Span4Mux_v I__9291 (
            .O(N__39273),
            .I(N__39241));
    Span4Mux_h I__9290 (
            .O(N__39270),
            .I(N__39232));
    Span4Mux_v I__9289 (
            .O(N__39267),
            .I(N__39232));
    Span4Mux_v I__9288 (
            .O(N__39260),
            .I(N__39232));
    Span4Mux_v I__9287 (
            .O(N__39253),
            .I(N__39232));
    LocalMux I__9286 (
            .O(N__39250),
            .I(N__39229));
    Span4Mux_s3_h I__9285 (
            .O(N__39247),
            .I(N__39224));
    Span4Mux_v I__9284 (
            .O(N__39244),
            .I(N__39224));
    Sp12to4 I__9283 (
            .O(N__39241),
            .I(N__39219));
    Sp12to4 I__9282 (
            .O(N__39232),
            .I(N__39219));
    Odrv12 I__9281 (
            .O(N__39229),
            .I(\ALU.aluOut_11 ));
    Odrv4 I__9280 (
            .O(N__39224),
            .I(\ALU.aluOut_11 ));
    Odrv12 I__9279 (
            .O(N__39219),
            .I(\ALU.aluOut_11 ));
    InMux I__9278 (
            .O(N__39212),
            .I(N__39209));
    LocalMux I__9277 (
            .O(N__39209),
            .I(N__39206));
    Odrv4 I__9276 (
            .O(N__39206),
            .I(\ALU.un9_addsub_cry_10_c_RNI9C0KZ0Z9 ));
    InMux I__9275 (
            .O(N__39203),
            .I(\ALU.un9_addsub_cry_10 ));
    InMux I__9274 (
            .O(N__39200),
            .I(N__39196));
    InMux I__9273 (
            .O(N__39199),
            .I(N__39193));
    LocalMux I__9272 (
            .O(N__39196),
            .I(N__39188));
    LocalMux I__9271 (
            .O(N__39193),
            .I(N__39188));
    Odrv12 I__9270 (
            .O(N__39188),
            .I(\ALU.N_361 ));
    InMux I__9269 (
            .O(N__39185),
            .I(N__39182));
    LocalMux I__9268 (
            .O(N__39182),
            .I(N__39177));
    InMux I__9267 (
            .O(N__39181),
            .I(N__39174));
    InMux I__9266 (
            .O(N__39180),
            .I(N__39171));
    Span4Mux_h I__9265 (
            .O(N__39177),
            .I(N__39168));
    LocalMux I__9264 (
            .O(N__39174),
            .I(N__39165));
    LocalMux I__9263 (
            .O(N__39171),
            .I(N__39162));
    Span4Mux_h I__9262 (
            .O(N__39168),
            .I(N__39157));
    Span4Mux_h I__9261 (
            .O(N__39165),
            .I(N__39157));
    Odrv4 I__9260 (
            .O(N__39162),
            .I(\ALU.N_244 ));
    Odrv4 I__9259 (
            .O(N__39157),
            .I(\ALU.N_244 ));
    InMux I__9258 (
            .O(N__39152),
            .I(N__39134));
    InMux I__9257 (
            .O(N__39151),
            .I(N__39134));
    InMux I__9256 (
            .O(N__39150),
            .I(N__39129));
    InMux I__9255 (
            .O(N__39149),
            .I(N__39129));
    InMux I__9254 (
            .O(N__39148),
            .I(N__39122));
    InMux I__9253 (
            .O(N__39147),
            .I(N__39122));
    InMux I__9252 (
            .O(N__39146),
            .I(N__39122));
    InMux I__9251 (
            .O(N__39145),
            .I(N__39117));
    InMux I__9250 (
            .O(N__39144),
            .I(N__39117));
    InMux I__9249 (
            .O(N__39143),
            .I(N__39112));
    InMux I__9248 (
            .O(N__39142),
            .I(N__39112));
    InMux I__9247 (
            .O(N__39141),
            .I(N__39109));
    CascadeMux I__9246 (
            .O(N__39140),
            .I(N__39106));
    CascadeMux I__9245 (
            .O(N__39139),
            .I(N__39102));
    LocalMux I__9244 (
            .O(N__39134),
            .I(N__39099));
    LocalMux I__9243 (
            .O(N__39129),
            .I(N__39088));
    LocalMux I__9242 (
            .O(N__39122),
            .I(N__39088));
    LocalMux I__9241 (
            .O(N__39117),
            .I(N__39088));
    LocalMux I__9240 (
            .O(N__39112),
            .I(N__39088));
    LocalMux I__9239 (
            .O(N__39109),
            .I(N__39088));
    InMux I__9238 (
            .O(N__39106),
            .I(N__39085));
    InMux I__9237 (
            .O(N__39105),
            .I(N__39071));
    InMux I__9236 (
            .O(N__39102),
            .I(N__39071));
    Span4Mux_v I__9235 (
            .O(N__39099),
            .I(N__39062));
    Span4Mux_v I__9234 (
            .O(N__39088),
            .I(N__39062));
    LocalMux I__9233 (
            .O(N__39085),
            .I(N__39062));
    CascadeMux I__9232 (
            .O(N__39084),
            .I(N__39058));
    CascadeMux I__9231 (
            .O(N__39083),
            .I(N__39055));
    CascadeMux I__9230 (
            .O(N__39082),
            .I(N__39050));
    CascadeMux I__9229 (
            .O(N__39081),
            .I(N__39047));
    CascadeMux I__9228 (
            .O(N__39080),
            .I(N__39041));
    CascadeMux I__9227 (
            .O(N__39079),
            .I(N__39038));
    CascadeMux I__9226 (
            .O(N__39078),
            .I(N__39033));
    CascadeMux I__9225 (
            .O(N__39077),
            .I(N__39030));
    InMux I__9224 (
            .O(N__39076),
            .I(N__39026));
    LocalMux I__9223 (
            .O(N__39071),
            .I(N__39023));
    InMux I__9222 (
            .O(N__39070),
            .I(N__39019));
    CascadeMux I__9221 (
            .O(N__39069),
            .I(N__39007));
    Span4Mux_h I__9220 (
            .O(N__39062),
            .I(N__39002));
    InMux I__9219 (
            .O(N__39061),
            .I(N__38995));
    InMux I__9218 (
            .O(N__39058),
            .I(N__38995));
    InMux I__9217 (
            .O(N__39055),
            .I(N__38995));
    InMux I__9216 (
            .O(N__39054),
            .I(N__38986));
    InMux I__9215 (
            .O(N__39053),
            .I(N__38986));
    InMux I__9214 (
            .O(N__39050),
            .I(N__38986));
    InMux I__9213 (
            .O(N__39047),
            .I(N__38986));
    InMux I__9212 (
            .O(N__39046),
            .I(N__38975));
    InMux I__9211 (
            .O(N__39045),
            .I(N__38975));
    InMux I__9210 (
            .O(N__39044),
            .I(N__38975));
    InMux I__9209 (
            .O(N__39041),
            .I(N__38975));
    InMux I__9208 (
            .O(N__39038),
            .I(N__38975));
    InMux I__9207 (
            .O(N__39037),
            .I(N__38962));
    InMux I__9206 (
            .O(N__39036),
            .I(N__38955));
    InMux I__9205 (
            .O(N__39033),
            .I(N__38955));
    InMux I__9204 (
            .O(N__39030),
            .I(N__38955));
    InMux I__9203 (
            .O(N__39029),
            .I(N__38952));
    LocalMux I__9202 (
            .O(N__39026),
            .I(N__38949));
    Span4Mux_h I__9201 (
            .O(N__39023),
            .I(N__38946));
    InMux I__9200 (
            .O(N__39022),
            .I(N__38943));
    LocalMux I__9199 (
            .O(N__39019),
            .I(N__38940));
    InMux I__9198 (
            .O(N__39018),
            .I(N__38933));
    InMux I__9197 (
            .O(N__39017),
            .I(N__38933));
    InMux I__9196 (
            .O(N__39016),
            .I(N__38933));
    InMux I__9195 (
            .O(N__39015),
            .I(N__38930));
    InMux I__9194 (
            .O(N__39014),
            .I(N__38927));
    InMux I__9193 (
            .O(N__39013),
            .I(N__38924));
    InMux I__9192 (
            .O(N__39012),
            .I(N__38919));
    InMux I__9191 (
            .O(N__39011),
            .I(N__38912));
    InMux I__9190 (
            .O(N__39010),
            .I(N__38912));
    InMux I__9189 (
            .O(N__39007),
            .I(N__38912));
    InMux I__9188 (
            .O(N__39006),
            .I(N__38907));
    InMux I__9187 (
            .O(N__39005),
            .I(N__38907));
    Span4Mux_v I__9186 (
            .O(N__39002),
            .I(N__38902));
    LocalMux I__9185 (
            .O(N__38995),
            .I(N__38902));
    LocalMux I__9184 (
            .O(N__38986),
            .I(N__38897));
    LocalMux I__9183 (
            .O(N__38975),
            .I(N__38897));
    InMux I__9182 (
            .O(N__38974),
            .I(N__38892));
    InMux I__9181 (
            .O(N__38973),
            .I(N__38892));
    CascadeMux I__9180 (
            .O(N__38972),
            .I(N__38889));
    CascadeMux I__9179 (
            .O(N__38971),
            .I(N__38884));
    CascadeMux I__9178 (
            .O(N__38970),
            .I(N__38881));
    CascadeMux I__9177 (
            .O(N__38969),
            .I(N__38878));
    CascadeMux I__9176 (
            .O(N__38968),
            .I(N__38875));
    InMux I__9175 (
            .O(N__38967),
            .I(N__38868));
    InMux I__9174 (
            .O(N__38966),
            .I(N__38868));
    InMux I__9173 (
            .O(N__38965),
            .I(N__38868));
    LocalMux I__9172 (
            .O(N__38962),
            .I(N__38865));
    LocalMux I__9171 (
            .O(N__38955),
            .I(N__38860));
    LocalMux I__9170 (
            .O(N__38952),
            .I(N__38860));
    Span4Mux_h I__9169 (
            .O(N__38949),
            .I(N__38855));
    Span4Mux_v I__9168 (
            .O(N__38946),
            .I(N__38855));
    LocalMux I__9167 (
            .O(N__38943),
            .I(N__38850));
    Span4Mux_v I__9166 (
            .O(N__38940),
            .I(N__38850));
    LocalMux I__9165 (
            .O(N__38933),
            .I(N__38847));
    LocalMux I__9164 (
            .O(N__38930),
            .I(N__38840));
    LocalMux I__9163 (
            .O(N__38927),
            .I(N__38840));
    LocalMux I__9162 (
            .O(N__38924),
            .I(N__38840));
    InMux I__9161 (
            .O(N__38923),
            .I(N__38835));
    InMux I__9160 (
            .O(N__38922),
            .I(N__38835));
    LocalMux I__9159 (
            .O(N__38919),
            .I(N__38822));
    LocalMux I__9158 (
            .O(N__38912),
            .I(N__38822));
    LocalMux I__9157 (
            .O(N__38907),
            .I(N__38822));
    Span4Mux_s2_v I__9156 (
            .O(N__38902),
            .I(N__38822));
    Span4Mux_h I__9155 (
            .O(N__38897),
            .I(N__38822));
    LocalMux I__9154 (
            .O(N__38892),
            .I(N__38822));
    InMux I__9153 (
            .O(N__38889),
            .I(N__38819));
    InMux I__9152 (
            .O(N__38888),
            .I(N__38814));
    InMux I__9151 (
            .O(N__38887),
            .I(N__38814));
    InMux I__9150 (
            .O(N__38884),
            .I(N__38807));
    InMux I__9149 (
            .O(N__38881),
            .I(N__38807));
    InMux I__9148 (
            .O(N__38878),
            .I(N__38807));
    InMux I__9147 (
            .O(N__38875),
            .I(N__38804));
    LocalMux I__9146 (
            .O(N__38868),
            .I(N__38801));
    Span4Mux_v I__9145 (
            .O(N__38865),
            .I(N__38794));
    Span4Mux_h I__9144 (
            .O(N__38860),
            .I(N__38794));
    Span4Mux_v I__9143 (
            .O(N__38855),
            .I(N__38794));
    Span4Mux_h I__9142 (
            .O(N__38850),
            .I(N__38785));
    Span4Mux_v I__9141 (
            .O(N__38847),
            .I(N__38785));
    Span4Mux_v I__9140 (
            .O(N__38840),
            .I(N__38785));
    LocalMux I__9139 (
            .O(N__38835),
            .I(N__38785));
    Span4Mux_h I__9138 (
            .O(N__38822),
            .I(N__38782));
    LocalMux I__9137 (
            .O(N__38819),
            .I(aluParams_1));
    LocalMux I__9136 (
            .O(N__38814),
            .I(aluParams_1));
    LocalMux I__9135 (
            .O(N__38807),
            .I(aluParams_1));
    LocalMux I__9134 (
            .O(N__38804),
            .I(aluParams_1));
    Odrv4 I__9133 (
            .O(N__38801),
            .I(aluParams_1));
    Odrv4 I__9132 (
            .O(N__38794),
            .I(aluParams_1));
    Odrv4 I__9131 (
            .O(N__38785),
            .I(aluParams_1));
    Odrv4 I__9130 (
            .O(N__38782),
            .I(aluParams_1));
    InMux I__9129 (
            .O(N__38765),
            .I(N__38762));
    LocalMux I__9128 (
            .O(N__38762),
            .I(N__38759));
    Span4Mux_v I__9127 (
            .O(N__38759),
            .I(N__38756));
    Span4Mux_h I__9126 (
            .O(N__38756),
            .I(N__38752));
    InMux I__9125 (
            .O(N__38755),
            .I(N__38749));
    Odrv4 I__9124 (
            .O(N__38752),
            .I(\ALU.N_588 ));
    LocalMux I__9123 (
            .O(N__38749),
            .I(\ALU.N_588 ));
    InMux I__9122 (
            .O(N__38744),
            .I(N__38740));
    InMux I__9121 (
            .O(N__38743),
            .I(N__38736));
    LocalMux I__9120 (
            .O(N__38740),
            .I(N__38719));
    CascadeMux I__9119 (
            .O(N__38739),
            .I(N__38716));
    LocalMux I__9118 (
            .O(N__38736),
            .I(N__38710));
    InMux I__9117 (
            .O(N__38735),
            .I(N__38707));
    CascadeMux I__9116 (
            .O(N__38734),
            .I(N__38704));
    InMux I__9115 (
            .O(N__38733),
            .I(N__38701));
    InMux I__9114 (
            .O(N__38732),
            .I(N__38698));
    InMux I__9113 (
            .O(N__38731),
            .I(N__38693));
    InMux I__9112 (
            .O(N__38730),
            .I(N__38690));
    CascadeMux I__9111 (
            .O(N__38729),
            .I(N__38686));
    InMux I__9110 (
            .O(N__38728),
            .I(N__38682));
    CascadeMux I__9109 (
            .O(N__38727),
            .I(N__38679));
    InMux I__9108 (
            .O(N__38726),
            .I(N__38673));
    InMux I__9107 (
            .O(N__38725),
            .I(N__38668));
    InMux I__9106 (
            .O(N__38724),
            .I(N__38668));
    InMux I__9105 (
            .O(N__38723),
            .I(N__38663));
    InMux I__9104 (
            .O(N__38722),
            .I(N__38663));
    Span4Mux_v I__9103 (
            .O(N__38719),
            .I(N__38660));
    InMux I__9102 (
            .O(N__38716),
            .I(N__38657));
    CascadeMux I__9101 (
            .O(N__38715),
            .I(N__38654));
    CascadeMux I__9100 (
            .O(N__38714),
            .I(N__38649));
    InMux I__9099 (
            .O(N__38713),
            .I(N__38643));
    Span4Mux_h I__9098 (
            .O(N__38710),
            .I(N__38640));
    LocalMux I__9097 (
            .O(N__38707),
            .I(N__38637));
    InMux I__9096 (
            .O(N__38704),
            .I(N__38634));
    LocalMux I__9095 (
            .O(N__38701),
            .I(N__38631));
    LocalMux I__9094 (
            .O(N__38698),
            .I(N__38628));
    InMux I__9093 (
            .O(N__38697),
            .I(N__38623));
    InMux I__9092 (
            .O(N__38696),
            .I(N__38623));
    LocalMux I__9091 (
            .O(N__38693),
            .I(N__38620));
    LocalMux I__9090 (
            .O(N__38690),
            .I(N__38617));
    InMux I__9089 (
            .O(N__38689),
            .I(N__38610));
    InMux I__9088 (
            .O(N__38686),
            .I(N__38610));
    InMux I__9087 (
            .O(N__38685),
            .I(N__38610));
    LocalMux I__9086 (
            .O(N__38682),
            .I(N__38607));
    InMux I__9085 (
            .O(N__38679),
            .I(N__38604));
    CascadeMux I__9084 (
            .O(N__38678),
            .I(N__38600));
    CascadeMux I__9083 (
            .O(N__38677),
            .I(N__38597));
    CascadeMux I__9082 (
            .O(N__38676),
            .I(N__38594));
    LocalMux I__9081 (
            .O(N__38673),
            .I(N__38584));
    LocalMux I__9080 (
            .O(N__38668),
            .I(N__38584));
    LocalMux I__9079 (
            .O(N__38663),
            .I(N__38584));
    Sp12to4 I__9078 (
            .O(N__38660),
            .I(N__38579));
    LocalMux I__9077 (
            .O(N__38657),
            .I(N__38579));
    InMux I__9076 (
            .O(N__38654),
            .I(N__38576));
    InMux I__9075 (
            .O(N__38653),
            .I(N__38571));
    InMux I__9074 (
            .O(N__38652),
            .I(N__38571));
    InMux I__9073 (
            .O(N__38649),
            .I(N__38566));
    InMux I__9072 (
            .O(N__38648),
            .I(N__38566));
    InMux I__9071 (
            .O(N__38647),
            .I(N__38561));
    InMux I__9070 (
            .O(N__38646),
            .I(N__38561));
    LocalMux I__9069 (
            .O(N__38643),
            .I(N__38556));
    Span4Mux_v I__9068 (
            .O(N__38640),
            .I(N__38553));
    Span4Mux_v I__9067 (
            .O(N__38637),
            .I(N__38548));
    LocalMux I__9066 (
            .O(N__38634),
            .I(N__38548));
    Span4Mux_s3_h I__9065 (
            .O(N__38631),
            .I(N__38541));
    Span4Mux_v I__9064 (
            .O(N__38628),
            .I(N__38541));
    LocalMux I__9063 (
            .O(N__38623),
            .I(N__38541));
    Span4Mux_h I__9062 (
            .O(N__38620),
            .I(N__38529));
    Span4Mux_h I__9061 (
            .O(N__38617),
            .I(N__38529));
    LocalMux I__9060 (
            .O(N__38610),
            .I(N__38529));
    Span4Mux_h I__9059 (
            .O(N__38607),
            .I(N__38529));
    LocalMux I__9058 (
            .O(N__38604),
            .I(N__38529));
    CascadeMux I__9057 (
            .O(N__38603),
            .I(N__38525));
    InMux I__9056 (
            .O(N__38600),
            .I(N__38522));
    InMux I__9055 (
            .O(N__38597),
            .I(N__38517));
    InMux I__9054 (
            .O(N__38594),
            .I(N__38517));
    InMux I__9053 (
            .O(N__38593),
            .I(N__38514));
    InMux I__9052 (
            .O(N__38592),
            .I(N__38509));
    InMux I__9051 (
            .O(N__38591),
            .I(N__38509));
    Sp12to4 I__9050 (
            .O(N__38584),
            .I(N__38504));
    Span12Mux_h I__9049 (
            .O(N__38579),
            .I(N__38504));
    LocalMux I__9048 (
            .O(N__38576),
            .I(N__38495));
    LocalMux I__9047 (
            .O(N__38571),
            .I(N__38495));
    LocalMux I__9046 (
            .O(N__38566),
            .I(N__38495));
    LocalMux I__9045 (
            .O(N__38561),
            .I(N__38495));
    InMux I__9044 (
            .O(N__38560),
            .I(N__38490));
    InMux I__9043 (
            .O(N__38559),
            .I(N__38490));
    Span4Mux_h I__9042 (
            .O(N__38556),
            .I(N__38485));
    Span4Mux_v I__9041 (
            .O(N__38553),
            .I(N__38485));
    Span4Mux_h I__9040 (
            .O(N__38548),
            .I(N__38480));
    Span4Mux_h I__9039 (
            .O(N__38541),
            .I(N__38480));
    InMux I__9038 (
            .O(N__38540),
            .I(N__38477));
    Span4Mux_v I__9037 (
            .O(N__38529),
            .I(N__38474));
    InMux I__9036 (
            .O(N__38528),
            .I(N__38469));
    InMux I__9035 (
            .O(N__38525),
            .I(N__38469));
    LocalMux I__9034 (
            .O(N__38522),
            .I(aluParams_2));
    LocalMux I__9033 (
            .O(N__38517),
            .I(aluParams_2));
    LocalMux I__9032 (
            .O(N__38514),
            .I(aluParams_2));
    LocalMux I__9031 (
            .O(N__38509),
            .I(aluParams_2));
    Odrv12 I__9030 (
            .O(N__38504),
            .I(aluParams_2));
    Odrv12 I__9029 (
            .O(N__38495),
            .I(aluParams_2));
    LocalMux I__9028 (
            .O(N__38490),
            .I(aluParams_2));
    Odrv4 I__9027 (
            .O(N__38485),
            .I(aluParams_2));
    Odrv4 I__9026 (
            .O(N__38480),
            .I(aluParams_2));
    LocalMux I__9025 (
            .O(N__38477),
            .I(aluParams_2));
    Odrv4 I__9024 (
            .O(N__38474),
            .I(aluParams_2));
    LocalMux I__9023 (
            .O(N__38469),
            .I(aluParams_2));
    InMux I__9022 (
            .O(N__38444),
            .I(N__38441));
    LocalMux I__9021 (
            .O(N__38441),
            .I(N__38438));
    Span4Mux_v I__9020 (
            .O(N__38438),
            .I(N__38433));
    InMux I__9019 (
            .O(N__38437),
            .I(N__38428));
    InMux I__9018 (
            .O(N__38436),
            .I(N__38425));
    Sp12to4 I__9017 (
            .O(N__38433),
            .I(N__38422));
    InMux I__9016 (
            .O(N__38432),
            .I(N__38417));
    InMux I__9015 (
            .O(N__38431),
            .I(N__38417));
    LocalMux I__9014 (
            .O(N__38428),
            .I(N__38414));
    LocalMux I__9013 (
            .O(N__38425),
            .I(\ALU.N_590 ));
    Odrv12 I__9012 (
            .O(N__38422),
            .I(\ALU.N_590 ));
    LocalMux I__9011 (
            .O(N__38417),
            .I(\ALU.N_590 ));
    Odrv4 I__9010 (
            .O(N__38414),
            .I(\ALU.N_590 ));
    InMux I__9009 (
            .O(N__38405),
            .I(N__38402));
    LocalMux I__9008 (
            .O(N__38402),
            .I(N__38398));
    CascadeMux I__9007 (
            .O(N__38401),
            .I(N__38395));
    Span4Mux_v I__9006 (
            .O(N__38398),
            .I(N__38392));
    InMux I__9005 (
            .O(N__38395),
            .I(N__38388));
    Span4Mux_h I__9004 (
            .O(N__38392),
            .I(N__38385));
    InMux I__9003 (
            .O(N__38391),
            .I(N__38382));
    LocalMux I__9002 (
            .O(N__38388),
            .I(\ALU.eZ0Z_9 ));
    Odrv4 I__9001 (
            .O(N__38385),
            .I(\ALU.eZ0Z_9 ));
    LocalMux I__9000 (
            .O(N__38382),
            .I(\ALU.eZ0Z_9 ));
    InMux I__8999 (
            .O(N__38375),
            .I(N__38372));
    LocalMux I__8998 (
            .O(N__38372),
            .I(N__38368));
    InMux I__8997 (
            .O(N__38371),
            .I(N__38365));
    Span4Mux_v I__8996 (
            .O(N__38368),
            .I(N__38361));
    LocalMux I__8995 (
            .O(N__38365),
            .I(N__38358));
    InMux I__8994 (
            .O(N__38364),
            .I(N__38355));
    Span4Mux_h I__8993 (
            .O(N__38361),
            .I(N__38350));
    Span4Mux_v I__8992 (
            .O(N__38358),
            .I(N__38350));
    LocalMux I__8991 (
            .O(N__38355),
            .I(\ALU.aZ0Z_9 ));
    Odrv4 I__8990 (
            .O(N__38350),
            .I(\ALU.aZ0Z_9 ));
    InMux I__8989 (
            .O(N__38345),
            .I(N__38342));
    LocalMux I__8988 (
            .O(N__38342),
            .I(\ALU.e_RNIR49HZ0Z_9 ));
    CascadeMux I__8987 (
            .O(N__38339),
            .I(N__38333));
    InMux I__8986 (
            .O(N__38338),
            .I(N__38326));
    CascadeMux I__8985 (
            .O(N__38337),
            .I(N__38319));
    CascadeMux I__8984 (
            .O(N__38336),
            .I(N__38312));
    InMux I__8983 (
            .O(N__38333),
            .I(N__38303));
    InMux I__8982 (
            .O(N__38332),
            .I(N__38300));
    InMux I__8981 (
            .O(N__38331),
            .I(N__38292));
    InMux I__8980 (
            .O(N__38330),
            .I(N__38292));
    InMux I__8979 (
            .O(N__38329),
            .I(N__38292));
    LocalMux I__8978 (
            .O(N__38326),
            .I(N__38288));
    InMux I__8977 (
            .O(N__38325),
            .I(N__38285));
    InMux I__8976 (
            .O(N__38324),
            .I(N__38282));
    InMux I__8975 (
            .O(N__38323),
            .I(N__38275));
    InMux I__8974 (
            .O(N__38322),
            .I(N__38275));
    InMux I__8973 (
            .O(N__38319),
            .I(N__38275));
    InMux I__8972 (
            .O(N__38318),
            .I(N__38269));
    InMux I__8971 (
            .O(N__38317),
            .I(N__38264));
    InMux I__8970 (
            .O(N__38316),
            .I(N__38264));
    InMux I__8969 (
            .O(N__38315),
            .I(N__38257));
    InMux I__8968 (
            .O(N__38312),
            .I(N__38257));
    InMux I__8967 (
            .O(N__38311),
            .I(N__38257));
    InMux I__8966 (
            .O(N__38310),
            .I(N__38250));
    InMux I__8965 (
            .O(N__38309),
            .I(N__38250));
    InMux I__8964 (
            .O(N__38308),
            .I(N__38250));
    InMux I__8963 (
            .O(N__38307),
            .I(N__38242));
    InMux I__8962 (
            .O(N__38306),
            .I(N__38242));
    LocalMux I__8961 (
            .O(N__38303),
            .I(N__38239));
    LocalMux I__8960 (
            .O(N__38300),
            .I(N__38236));
    InMux I__8959 (
            .O(N__38299),
            .I(N__38233));
    LocalMux I__8958 (
            .O(N__38292),
            .I(N__38230));
    InMux I__8957 (
            .O(N__38291),
            .I(N__38227));
    Span4Mux_h I__8956 (
            .O(N__38288),
            .I(N__38222));
    LocalMux I__8955 (
            .O(N__38285),
            .I(N__38219));
    LocalMux I__8954 (
            .O(N__38282),
            .I(N__38214));
    LocalMux I__8953 (
            .O(N__38275),
            .I(N__38214));
    InMux I__8952 (
            .O(N__38274),
            .I(N__38210));
    CascadeMux I__8951 (
            .O(N__38273),
            .I(N__38207));
    InMux I__8950 (
            .O(N__38272),
            .I(N__38204));
    LocalMux I__8949 (
            .O(N__38269),
            .I(N__38199));
    LocalMux I__8948 (
            .O(N__38264),
            .I(N__38199));
    LocalMux I__8947 (
            .O(N__38257),
            .I(N__38196));
    LocalMux I__8946 (
            .O(N__38250),
            .I(N__38193));
    InMux I__8945 (
            .O(N__38249),
            .I(N__38183));
    InMux I__8944 (
            .O(N__38248),
            .I(N__38183));
    InMux I__8943 (
            .O(N__38247),
            .I(N__38183));
    LocalMux I__8942 (
            .O(N__38242),
            .I(N__38180));
    Span4Mux_v I__8941 (
            .O(N__38239),
            .I(N__38173));
    Span4Mux_v I__8940 (
            .O(N__38236),
            .I(N__38170));
    LocalMux I__8939 (
            .O(N__38233),
            .I(N__38163));
    Span4Mux_v I__8938 (
            .O(N__38230),
            .I(N__38163));
    LocalMux I__8937 (
            .O(N__38227),
            .I(N__38163));
    InMux I__8936 (
            .O(N__38226),
            .I(N__38158));
    InMux I__8935 (
            .O(N__38225),
            .I(N__38158));
    Span4Mux_v I__8934 (
            .O(N__38222),
            .I(N__38153));
    Span4Mux_h I__8933 (
            .O(N__38219),
            .I(N__38153));
    Span4Mux_h I__8932 (
            .O(N__38214),
            .I(N__38150));
    InMux I__8931 (
            .O(N__38213),
            .I(N__38147));
    LocalMux I__8930 (
            .O(N__38210),
            .I(N__38144));
    InMux I__8929 (
            .O(N__38207),
            .I(N__38141));
    LocalMux I__8928 (
            .O(N__38204),
            .I(N__38138));
    Span4Mux_v I__8927 (
            .O(N__38199),
            .I(N__38131));
    Span4Mux_v I__8926 (
            .O(N__38196),
            .I(N__38131));
    Span4Mux_s1_h I__8925 (
            .O(N__38193),
            .I(N__38131));
    InMux I__8924 (
            .O(N__38192),
            .I(N__38126));
    InMux I__8923 (
            .O(N__38191),
            .I(N__38126));
    InMux I__8922 (
            .O(N__38190),
            .I(N__38123));
    LocalMux I__8921 (
            .O(N__38183),
            .I(N__38120));
    Span12Mux_s4_v I__8920 (
            .O(N__38180),
            .I(N__38117));
    InMux I__8919 (
            .O(N__38179),
            .I(N__38114));
    InMux I__8918 (
            .O(N__38178),
            .I(N__38111));
    InMux I__8917 (
            .O(N__38177),
            .I(N__38108));
    InMux I__8916 (
            .O(N__38176),
            .I(N__38105));
    Span4Mux_s2_h I__8915 (
            .O(N__38173),
            .I(N__38100));
    Span4Mux_v I__8914 (
            .O(N__38170),
            .I(N__38100));
    Span4Mux_v I__8913 (
            .O(N__38163),
            .I(N__38095));
    LocalMux I__8912 (
            .O(N__38158),
            .I(N__38095));
    Span4Mux_h I__8911 (
            .O(N__38153),
            .I(N__38092));
    Span4Mux_v I__8910 (
            .O(N__38150),
            .I(N__38085));
    LocalMux I__8909 (
            .O(N__38147),
            .I(N__38085));
    Span4Mux_v I__8908 (
            .O(N__38144),
            .I(N__38085));
    LocalMux I__8907 (
            .O(N__38141),
            .I(N__38076));
    Span4Mux_h I__8906 (
            .O(N__38138),
            .I(N__38076));
    Span4Mux_h I__8905 (
            .O(N__38131),
            .I(N__38076));
    LocalMux I__8904 (
            .O(N__38126),
            .I(N__38076));
    LocalMux I__8903 (
            .O(N__38123),
            .I(\ALU.N_252_0 ));
    Odrv12 I__8902 (
            .O(N__38120),
            .I(\ALU.N_252_0 ));
    Odrv12 I__8901 (
            .O(N__38117),
            .I(\ALU.N_252_0 ));
    LocalMux I__8900 (
            .O(N__38114),
            .I(\ALU.N_252_0 ));
    LocalMux I__8899 (
            .O(N__38111),
            .I(\ALU.N_252_0 ));
    LocalMux I__8898 (
            .O(N__38108),
            .I(\ALU.N_252_0 ));
    LocalMux I__8897 (
            .O(N__38105),
            .I(\ALU.N_252_0 ));
    Odrv4 I__8896 (
            .O(N__38100),
            .I(\ALU.N_252_0 ));
    Odrv4 I__8895 (
            .O(N__38095),
            .I(\ALU.N_252_0 ));
    Odrv4 I__8894 (
            .O(N__38092),
            .I(\ALU.N_252_0 ));
    Odrv4 I__8893 (
            .O(N__38085),
            .I(\ALU.N_252_0 ));
    Odrv4 I__8892 (
            .O(N__38076),
            .I(\ALU.N_252_0 ));
    CascadeMux I__8891 (
            .O(N__38051),
            .I(N__38048));
    InMux I__8890 (
            .O(N__38048),
            .I(N__38042));
    CascadeMux I__8889 (
            .O(N__38047),
            .I(N__38038));
    CascadeMux I__8888 (
            .O(N__38046),
            .I(N__38030));
    CascadeMux I__8887 (
            .O(N__38045),
            .I(N__38019));
    LocalMux I__8886 (
            .O(N__38042),
            .I(N__38016));
    InMux I__8885 (
            .O(N__38041),
            .I(N__38013));
    InMux I__8884 (
            .O(N__38038),
            .I(N__38006));
    InMux I__8883 (
            .O(N__38037),
            .I(N__38006));
    InMux I__8882 (
            .O(N__38036),
            .I(N__38006));
    InMux I__8881 (
            .O(N__38035),
            .I(N__38003));
    InMux I__8880 (
            .O(N__38034),
            .I(N__37998));
    InMux I__8879 (
            .O(N__38033),
            .I(N__37987));
    InMux I__8878 (
            .O(N__38030),
            .I(N__37987));
    InMux I__8877 (
            .O(N__38029),
            .I(N__37987));
    InMux I__8876 (
            .O(N__38028),
            .I(N__37982));
    InMux I__8875 (
            .O(N__38027),
            .I(N__37976));
    InMux I__8874 (
            .O(N__38026),
            .I(N__37976));
    InMux I__8873 (
            .O(N__38025),
            .I(N__37969));
    InMux I__8872 (
            .O(N__38024),
            .I(N__37969));
    InMux I__8871 (
            .O(N__38023),
            .I(N__37969));
    InMux I__8870 (
            .O(N__38022),
            .I(N__37963));
    InMux I__8869 (
            .O(N__38019),
            .I(N__37963));
    Span4Mux_h I__8868 (
            .O(N__38016),
            .I(N__37956));
    LocalMux I__8867 (
            .O(N__38013),
            .I(N__37956));
    LocalMux I__8866 (
            .O(N__38006),
            .I(N__37953));
    LocalMux I__8865 (
            .O(N__38003),
            .I(N__37950));
    InMux I__8864 (
            .O(N__38002),
            .I(N__37947));
    InMux I__8863 (
            .O(N__38001),
            .I(N__37944));
    LocalMux I__8862 (
            .O(N__37998),
            .I(N__37941));
    InMux I__8861 (
            .O(N__37997),
            .I(N__37938));
    InMux I__8860 (
            .O(N__37996),
            .I(N__37926));
    InMux I__8859 (
            .O(N__37995),
            .I(N__37926));
    InMux I__8858 (
            .O(N__37994),
            .I(N__37926));
    LocalMux I__8857 (
            .O(N__37987),
            .I(N__37923));
    InMux I__8856 (
            .O(N__37986),
            .I(N__37918));
    InMux I__8855 (
            .O(N__37985),
            .I(N__37918));
    LocalMux I__8854 (
            .O(N__37982),
            .I(N__37915));
    InMux I__8853 (
            .O(N__37981),
            .I(N__37912));
    LocalMux I__8852 (
            .O(N__37976),
            .I(N__37907));
    LocalMux I__8851 (
            .O(N__37969),
            .I(N__37907));
    InMux I__8850 (
            .O(N__37968),
            .I(N__37904));
    LocalMux I__8849 (
            .O(N__37963),
            .I(N__37901));
    InMux I__8848 (
            .O(N__37962),
            .I(N__37898));
    InMux I__8847 (
            .O(N__37961),
            .I(N__37895));
    Span4Mux_v I__8846 (
            .O(N__37956),
            .I(N__37891));
    Span4Mux_v I__8845 (
            .O(N__37953),
            .I(N__37888));
    Span4Mux_v I__8844 (
            .O(N__37950),
            .I(N__37883));
    LocalMux I__8843 (
            .O(N__37947),
            .I(N__37883));
    LocalMux I__8842 (
            .O(N__37944),
            .I(N__37876));
    Span4Mux_h I__8841 (
            .O(N__37941),
            .I(N__37876));
    LocalMux I__8840 (
            .O(N__37938),
            .I(N__37876));
    InMux I__8839 (
            .O(N__37937),
            .I(N__37867));
    InMux I__8838 (
            .O(N__37936),
            .I(N__37867));
    InMux I__8837 (
            .O(N__37935),
            .I(N__37867));
    InMux I__8836 (
            .O(N__37934),
            .I(N__37867));
    InMux I__8835 (
            .O(N__37933),
            .I(N__37864));
    LocalMux I__8834 (
            .O(N__37926),
            .I(N__37861));
    Span4Mux_v I__8833 (
            .O(N__37923),
            .I(N__37856));
    LocalMux I__8832 (
            .O(N__37918),
            .I(N__37856));
    Span4Mux_v I__8831 (
            .O(N__37915),
            .I(N__37847));
    LocalMux I__8830 (
            .O(N__37912),
            .I(N__37847));
    Span4Mux_h I__8829 (
            .O(N__37907),
            .I(N__37847));
    LocalMux I__8828 (
            .O(N__37904),
            .I(N__37847));
    Span12Mux_s3_v I__8827 (
            .O(N__37901),
            .I(N__37840));
    LocalMux I__8826 (
            .O(N__37898),
            .I(N__37840));
    LocalMux I__8825 (
            .O(N__37895),
            .I(N__37840));
    InMux I__8824 (
            .O(N__37894),
            .I(N__37837));
    Span4Mux_h I__8823 (
            .O(N__37891),
            .I(N__37834));
    Span4Mux_h I__8822 (
            .O(N__37888),
            .I(N__37827));
    Span4Mux_v I__8821 (
            .O(N__37883),
            .I(N__37827));
    Span4Mux_v I__8820 (
            .O(N__37876),
            .I(N__37827));
    LocalMux I__8819 (
            .O(N__37867),
            .I(N__37824));
    LocalMux I__8818 (
            .O(N__37864),
            .I(N__37819));
    Span4Mux_v I__8817 (
            .O(N__37861),
            .I(N__37819));
    Span4Mux_v I__8816 (
            .O(N__37856),
            .I(N__37816));
    Span4Mux_v I__8815 (
            .O(N__37847),
            .I(N__37813));
    Odrv12 I__8814 (
            .O(N__37840),
            .I(\ALU.aluOut_0 ));
    LocalMux I__8813 (
            .O(N__37837),
            .I(\ALU.aluOut_0 ));
    Odrv4 I__8812 (
            .O(N__37834),
            .I(\ALU.aluOut_0 ));
    Odrv4 I__8811 (
            .O(N__37827),
            .I(\ALU.aluOut_0 ));
    Odrv12 I__8810 (
            .O(N__37824),
            .I(\ALU.aluOut_0 ));
    Odrv4 I__8809 (
            .O(N__37819),
            .I(\ALU.aluOut_0 ));
    Odrv4 I__8808 (
            .O(N__37816),
            .I(\ALU.aluOut_0 ));
    Odrv4 I__8807 (
            .O(N__37813),
            .I(\ALU.aluOut_0 ));
    InMux I__8806 (
            .O(N__37796),
            .I(N__37793));
    LocalMux I__8805 (
            .O(N__37793),
            .I(N__37790));
    Odrv4 I__8804 (
            .O(N__37790),
            .I(\ALU.a0_b_2 ));
    InMux I__8803 (
            .O(N__37787),
            .I(N__37783));
    CascadeMux I__8802 (
            .O(N__37786),
            .I(N__37780));
    LocalMux I__8801 (
            .O(N__37783),
            .I(N__37777));
    InMux I__8800 (
            .O(N__37780),
            .I(N__37774));
    Span4Mux_v I__8799 (
            .O(N__37777),
            .I(N__37770));
    LocalMux I__8798 (
            .O(N__37774),
            .I(N__37764));
    InMux I__8797 (
            .O(N__37773),
            .I(N__37754));
    Span4Mux_h I__8796 (
            .O(N__37770),
            .I(N__37751));
    InMux I__8795 (
            .O(N__37769),
            .I(N__37746));
    InMux I__8794 (
            .O(N__37768),
            .I(N__37746));
    CascadeMux I__8793 (
            .O(N__37767),
            .I(N__37743));
    Span4Mux_h I__8792 (
            .O(N__37764),
            .I(N__37738));
    InMux I__8791 (
            .O(N__37763),
            .I(N__37733));
    InMux I__8790 (
            .O(N__37762),
            .I(N__37733));
    InMux I__8789 (
            .O(N__37761),
            .I(N__37725));
    InMux I__8788 (
            .O(N__37760),
            .I(N__37725));
    InMux I__8787 (
            .O(N__37759),
            .I(N__37722));
    CascadeMux I__8786 (
            .O(N__37758),
            .I(N__37719));
    InMux I__8785 (
            .O(N__37757),
            .I(N__37712));
    LocalMux I__8784 (
            .O(N__37754),
            .I(N__37709));
    Span4Mux_h I__8783 (
            .O(N__37751),
            .I(N__37704));
    LocalMux I__8782 (
            .O(N__37746),
            .I(N__37704));
    InMux I__8781 (
            .O(N__37743),
            .I(N__37699));
    InMux I__8780 (
            .O(N__37742),
            .I(N__37696));
    InMux I__8779 (
            .O(N__37741),
            .I(N__37693));
    Span4Mux_v I__8778 (
            .O(N__37738),
            .I(N__37688));
    LocalMux I__8777 (
            .O(N__37733),
            .I(N__37688));
    InMux I__8776 (
            .O(N__37732),
            .I(N__37683));
    InMux I__8775 (
            .O(N__37731),
            .I(N__37683));
    InMux I__8774 (
            .O(N__37730),
            .I(N__37680));
    LocalMux I__8773 (
            .O(N__37725),
            .I(N__37675));
    LocalMux I__8772 (
            .O(N__37722),
            .I(N__37675));
    InMux I__8771 (
            .O(N__37719),
            .I(N__37672));
    InMux I__8770 (
            .O(N__37718),
            .I(N__37669));
    InMux I__8769 (
            .O(N__37717),
            .I(N__37664));
    InMux I__8768 (
            .O(N__37716),
            .I(N__37664));
    InMux I__8767 (
            .O(N__37715),
            .I(N__37661));
    LocalMux I__8766 (
            .O(N__37712),
            .I(N__37648));
    Span4Mux_h I__8765 (
            .O(N__37709),
            .I(N__37641));
    Span4Mux_v I__8764 (
            .O(N__37704),
            .I(N__37641));
    InMux I__8763 (
            .O(N__37703),
            .I(N__37636));
    InMux I__8762 (
            .O(N__37702),
            .I(N__37636));
    LocalMux I__8761 (
            .O(N__37699),
            .I(N__37633));
    LocalMux I__8760 (
            .O(N__37696),
            .I(N__37628));
    LocalMux I__8759 (
            .O(N__37693),
            .I(N__37628));
    Span4Mux_h I__8758 (
            .O(N__37688),
            .I(N__37623));
    LocalMux I__8757 (
            .O(N__37683),
            .I(N__37620));
    LocalMux I__8756 (
            .O(N__37680),
            .I(N__37617));
    Span4Mux_v I__8755 (
            .O(N__37675),
            .I(N__37614));
    LocalMux I__8754 (
            .O(N__37672),
            .I(N__37611));
    LocalMux I__8753 (
            .O(N__37669),
            .I(N__37608));
    LocalMux I__8752 (
            .O(N__37664),
            .I(N__37603));
    LocalMux I__8751 (
            .O(N__37661),
            .I(N__37603));
    InMux I__8750 (
            .O(N__37660),
            .I(N__37596));
    InMux I__8749 (
            .O(N__37659),
            .I(N__37596));
    InMux I__8748 (
            .O(N__37658),
            .I(N__37596));
    InMux I__8747 (
            .O(N__37657),
            .I(N__37593));
    InMux I__8746 (
            .O(N__37656),
            .I(N__37586));
    InMux I__8745 (
            .O(N__37655),
            .I(N__37586));
    InMux I__8744 (
            .O(N__37654),
            .I(N__37586));
    InMux I__8743 (
            .O(N__37653),
            .I(N__37583));
    InMux I__8742 (
            .O(N__37652),
            .I(N__37578));
    InMux I__8741 (
            .O(N__37651),
            .I(N__37578));
    Span4Mux_h I__8740 (
            .O(N__37648),
            .I(N__37575));
    InMux I__8739 (
            .O(N__37647),
            .I(N__37570));
    InMux I__8738 (
            .O(N__37646),
            .I(N__37570));
    Span4Mux_v I__8737 (
            .O(N__37641),
            .I(N__37567));
    LocalMux I__8736 (
            .O(N__37636),
            .I(N__37560));
    Span4Mux_v I__8735 (
            .O(N__37633),
            .I(N__37560));
    Span4Mux_v I__8734 (
            .O(N__37628),
            .I(N__37560));
    InMux I__8733 (
            .O(N__37627),
            .I(N__37555));
    InMux I__8732 (
            .O(N__37626),
            .I(N__37555));
    Span4Mux_h I__8731 (
            .O(N__37623),
            .I(N__37538));
    Span4Mux_s3_h I__8730 (
            .O(N__37620),
            .I(N__37538));
    Span4Mux_v I__8729 (
            .O(N__37617),
            .I(N__37538));
    Span4Mux_v I__8728 (
            .O(N__37614),
            .I(N__37538));
    Span4Mux_s3_h I__8727 (
            .O(N__37611),
            .I(N__37538));
    Span4Mux_v I__8726 (
            .O(N__37608),
            .I(N__37538));
    Span4Mux_v I__8725 (
            .O(N__37603),
            .I(N__37538));
    LocalMux I__8724 (
            .O(N__37596),
            .I(N__37538));
    LocalMux I__8723 (
            .O(N__37593),
            .I(N__37533));
    LocalMux I__8722 (
            .O(N__37586),
            .I(N__37533));
    LocalMux I__8721 (
            .O(N__37583),
            .I(\ALU.N_249_0_i ));
    LocalMux I__8720 (
            .O(N__37578),
            .I(\ALU.N_249_0_i ));
    Odrv4 I__8719 (
            .O(N__37575),
            .I(\ALU.N_249_0_i ));
    LocalMux I__8718 (
            .O(N__37570),
            .I(\ALU.N_249_0_i ));
    Odrv4 I__8717 (
            .O(N__37567),
            .I(\ALU.N_249_0_i ));
    Odrv4 I__8716 (
            .O(N__37560),
            .I(\ALU.N_249_0_i ));
    LocalMux I__8715 (
            .O(N__37555),
            .I(\ALU.N_249_0_i ));
    Odrv4 I__8714 (
            .O(N__37538),
            .I(\ALU.N_249_0_i ));
    Odrv12 I__8713 (
            .O(N__37533),
            .I(\ALU.N_249_0_i ));
    InMux I__8712 (
            .O(N__37514),
            .I(N__37510));
    InMux I__8711 (
            .O(N__37513),
            .I(N__37507));
    LocalMux I__8710 (
            .O(N__37510),
            .I(N__37504));
    LocalMux I__8709 (
            .O(N__37507),
            .I(N__37497));
    Span4Mux_v I__8708 (
            .O(N__37504),
            .I(N__37494));
    InMux I__8707 (
            .O(N__37503),
            .I(N__37491));
    CascadeMux I__8706 (
            .O(N__37502),
            .I(N__37481));
    CascadeMux I__8705 (
            .O(N__37501),
            .I(N__37476));
    InMux I__8704 (
            .O(N__37500),
            .I(N__37473));
    Span4Mux_v I__8703 (
            .O(N__37497),
            .I(N__37468));
    Span4Mux_s2_h I__8702 (
            .O(N__37494),
            .I(N__37463));
    LocalMux I__8701 (
            .O(N__37491),
            .I(N__37463));
    InMux I__8700 (
            .O(N__37490),
            .I(N__37456));
    InMux I__8699 (
            .O(N__37489),
            .I(N__37456));
    InMux I__8698 (
            .O(N__37488),
            .I(N__37456));
    InMux I__8697 (
            .O(N__37487),
            .I(N__37451));
    InMux I__8696 (
            .O(N__37486),
            .I(N__37451));
    InMux I__8695 (
            .O(N__37485),
            .I(N__37448));
    InMux I__8694 (
            .O(N__37484),
            .I(N__37444));
    InMux I__8693 (
            .O(N__37481),
            .I(N__37439));
    InMux I__8692 (
            .O(N__37480),
            .I(N__37439));
    InMux I__8691 (
            .O(N__37479),
            .I(N__37436));
    InMux I__8690 (
            .O(N__37476),
            .I(N__37433));
    LocalMux I__8689 (
            .O(N__37473),
            .I(N__37430));
    InMux I__8688 (
            .O(N__37472),
            .I(N__37420));
    InMux I__8687 (
            .O(N__37471),
            .I(N__37420));
    Span4Mux_s2_h I__8686 (
            .O(N__37468),
            .I(N__37406));
    Span4Mux_v I__8685 (
            .O(N__37463),
            .I(N__37406));
    LocalMux I__8684 (
            .O(N__37456),
            .I(N__37406));
    LocalMux I__8683 (
            .O(N__37451),
            .I(N__37406));
    LocalMux I__8682 (
            .O(N__37448),
            .I(N__37406));
    InMux I__8681 (
            .O(N__37447),
            .I(N__37403));
    LocalMux I__8680 (
            .O(N__37444),
            .I(N__37400));
    LocalMux I__8679 (
            .O(N__37439),
            .I(N__37397));
    LocalMux I__8678 (
            .O(N__37436),
            .I(N__37392));
    LocalMux I__8677 (
            .O(N__37433),
            .I(N__37392));
    Span4Mux_v I__8676 (
            .O(N__37430),
            .I(N__37388));
    InMux I__8675 (
            .O(N__37429),
            .I(N__37383));
    InMux I__8674 (
            .O(N__37428),
            .I(N__37383));
    InMux I__8673 (
            .O(N__37427),
            .I(N__37380));
    InMux I__8672 (
            .O(N__37426),
            .I(N__37377));
    CascadeMux I__8671 (
            .O(N__37425),
            .I(N__37373));
    LocalMux I__8670 (
            .O(N__37420),
            .I(N__37368));
    InMux I__8669 (
            .O(N__37419),
            .I(N__37365));
    InMux I__8668 (
            .O(N__37418),
            .I(N__37362));
    InMux I__8667 (
            .O(N__37417),
            .I(N__37359));
    Span4Mux_v I__8666 (
            .O(N__37406),
            .I(N__37356));
    LocalMux I__8665 (
            .O(N__37403),
            .I(N__37353));
    Span4Mux_s2_h I__8664 (
            .O(N__37400),
            .I(N__37350));
    Span4Mux_v I__8663 (
            .O(N__37397),
            .I(N__37342));
    Span4Mux_v I__8662 (
            .O(N__37392),
            .I(N__37342));
    InMux I__8661 (
            .O(N__37391),
            .I(N__37339));
    Span4Mux_v I__8660 (
            .O(N__37388),
            .I(N__37334));
    LocalMux I__8659 (
            .O(N__37383),
            .I(N__37334));
    LocalMux I__8658 (
            .O(N__37380),
            .I(N__37329));
    LocalMux I__8657 (
            .O(N__37377),
            .I(N__37329));
    InMux I__8656 (
            .O(N__37376),
            .I(N__37326));
    InMux I__8655 (
            .O(N__37373),
            .I(N__37319));
    InMux I__8654 (
            .O(N__37372),
            .I(N__37319));
    InMux I__8653 (
            .O(N__37371),
            .I(N__37319));
    Span4Mux_h I__8652 (
            .O(N__37368),
            .I(N__37313));
    LocalMux I__8651 (
            .O(N__37365),
            .I(N__37313));
    LocalMux I__8650 (
            .O(N__37362),
            .I(N__37302));
    LocalMux I__8649 (
            .O(N__37359),
            .I(N__37302));
    Span4Mux_s2_h I__8648 (
            .O(N__37356),
            .I(N__37302));
    Span4Mux_v I__8647 (
            .O(N__37353),
            .I(N__37302));
    Span4Mux_v I__8646 (
            .O(N__37350),
            .I(N__37302));
    InMux I__8645 (
            .O(N__37349),
            .I(N__37295));
    InMux I__8644 (
            .O(N__37348),
            .I(N__37295));
    InMux I__8643 (
            .O(N__37347),
            .I(N__37295));
    Span4Mux_h I__8642 (
            .O(N__37342),
            .I(N__37290));
    LocalMux I__8641 (
            .O(N__37339),
            .I(N__37290));
    Span4Mux_h I__8640 (
            .O(N__37334),
            .I(N__37287));
    Span4Mux_v I__8639 (
            .O(N__37329),
            .I(N__37280));
    LocalMux I__8638 (
            .O(N__37326),
            .I(N__37280));
    LocalMux I__8637 (
            .O(N__37319),
            .I(N__37280));
    InMux I__8636 (
            .O(N__37318),
            .I(N__37277));
    Span4Mux_v I__8635 (
            .O(N__37313),
            .I(N__37272));
    Span4Mux_h I__8634 (
            .O(N__37302),
            .I(N__37272));
    LocalMux I__8633 (
            .O(N__37295),
            .I(\ALU.aluOut_1 ));
    Odrv4 I__8632 (
            .O(N__37290),
            .I(\ALU.aluOut_1 ));
    Odrv4 I__8631 (
            .O(N__37287),
            .I(\ALU.aluOut_1 ));
    Odrv4 I__8630 (
            .O(N__37280),
            .I(\ALU.aluOut_1 ));
    LocalMux I__8629 (
            .O(N__37277),
            .I(\ALU.aluOut_1 ));
    Odrv4 I__8628 (
            .O(N__37272),
            .I(\ALU.aluOut_1 ));
    InMux I__8627 (
            .O(N__37259),
            .I(\ALU.un9_addsub_cry_0 ));
    InMux I__8626 (
            .O(N__37256),
            .I(N__37251));
    InMux I__8625 (
            .O(N__37255),
            .I(N__37246));
    InMux I__8624 (
            .O(N__37254),
            .I(N__37246));
    LocalMux I__8623 (
            .O(N__37251),
            .I(N__37241));
    LocalMux I__8622 (
            .O(N__37246),
            .I(N__37238));
    InMux I__8621 (
            .O(N__37245),
            .I(N__37228));
    InMux I__8620 (
            .O(N__37244),
            .I(N__37225));
    Span4Mux_v I__8619 (
            .O(N__37241),
            .I(N__37222));
    Span4Mux_v I__8618 (
            .O(N__37238),
            .I(N__37219));
    CascadeMux I__8617 (
            .O(N__37237),
            .I(N__37215));
    InMux I__8616 (
            .O(N__37236),
            .I(N__37211));
    InMux I__8615 (
            .O(N__37235),
            .I(N__37206));
    InMux I__8614 (
            .O(N__37234),
            .I(N__37206));
    CascadeMux I__8613 (
            .O(N__37233),
            .I(N__37196));
    InMux I__8612 (
            .O(N__37232),
            .I(N__37191));
    InMux I__8611 (
            .O(N__37231),
            .I(N__37188));
    LocalMux I__8610 (
            .O(N__37228),
            .I(N__37183));
    LocalMux I__8609 (
            .O(N__37225),
            .I(N__37183));
    Span4Mux_v I__8608 (
            .O(N__37222),
            .I(N__37180));
    Span4Mux_v I__8607 (
            .O(N__37219),
            .I(N__37177));
    InMux I__8606 (
            .O(N__37218),
            .I(N__37174));
    InMux I__8605 (
            .O(N__37215),
            .I(N__37169));
    InMux I__8604 (
            .O(N__37214),
            .I(N__37169));
    LocalMux I__8603 (
            .O(N__37211),
            .I(N__37164));
    LocalMux I__8602 (
            .O(N__37206),
            .I(N__37164));
    InMux I__8601 (
            .O(N__37205),
            .I(N__37159));
    InMux I__8600 (
            .O(N__37204),
            .I(N__37159));
    CascadeMux I__8599 (
            .O(N__37203),
            .I(N__37153));
    InMux I__8598 (
            .O(N__37202),
            .I(N__37146));
    InMux I__8597 (
            .O(N__37201),
            .I(N__37146));
    InMux I__8596 (
            .O(N__37200),
            .I(N__37146));
    InMux I__8595 (
            .O(N__37199),
            .I(N__37142));
    InMux I__8594 (
            .O(N__37196),
            .I(N__37139));
    InMux I__8593 (
            .O(N__37195),
            .I(N__37136));
    InMux I__8592 (
            .O(N__37194),
            .I(N__37133));
    LocalMux I__8591 (
            .O(N__37191),
            .I(N__37130));
    LocalMux I__8590 (
            .O(N__37188),
            .I(N__37125));
    Span4Mux_h I__8589 (
            .O(N__37183),
            .I(N__37125));
    Span4Mux_h I__8588 (
            .O(N__37180),
            .I(N__37122));
    Span4Mux_h I__8587 (
            .O(N__37177),
            .I(N__37119));
    LocalMux I__8586 (
            .O(N__37174),
            .I(N__37105));
    LocalMux I__8585 (
            .O(N__37169),
            .I(N__37105));
    Span4Mux_v I__8584 (
            .O(N__37164),
            .I(N__37105));
    LocalMux I__8583 (
            .O(N__37159),
            .I(N__37105));
    CascadeMux I__8582 (
            .O(N__37158),
            .I(N__37102));
    CascadeMux I__8581 (
            .O(N__37157),
            .I(N__37099));
    CascadeMux I__8580 (
            .O(N__37156),
            .I(N__37095));
    InMux I__8579 (
            .O(N__37153),
            .I(N__37091));
    LocalMux I__8578 (
            .O(N__37146),
            .I(N__37088));
    InMux I__8577 (
            .O(N__37145),
            .I(N__37085));
    LocalMux I__8576 (
            .O(N__37142),
            .I(N__37080));
    LocalMux I__8575 (
            .O(N__37139),
            .I(N__37080));
    LocalMux I__8574 (
            .O(N__37136),
            .I(N__37077));
    LocalMux I__8573 (
            .O(N__37133),
            .I(N__37074));
    Span4Mux_h I__8572 (
            .O(N__37130),
            .I(N__37069));
    Span4Mux_v I__8571 (
            .O(N__37125),
            .I(N__37069));
    Span4Mux_v I__8570 (
            .O(N__37122),
            .I(N__37064));
    Span4Mux_h I__8569 (
            .O(N__37119),
            .I(N__37064));
    InMux I__8568 (
            .O(N__37118),
            .I(N__37059));
    InMux I__8567 (
            .O(N__37117),
            .I(N__37059));
    InMux I__8566 (
            .O(N__37116),
            .I(N__37052));
    InMux I__8565 (
            .O(N__37115),
            .I(N__37052));
    InMux I__8564 (
            .O(N__37114),
            .I(N__37052));
    Span4Mux_h I__8563 (
            .O(N__37105),
            .I(N__37049));
    InMux I__8562 (
            .O(N__37102),
            .I(N__37044));
    InMux I__8561 (
            .O(N__37099),
            .I(N__37044));
    InMux I__8560 (
            .O(N__37098),
            .I(N__37037));
    InMux I__8559 (
            .O(N__37095),
            .I(N__37037));
    InMux I__8558 (
            .O(N__37094),
            .I(N__37037));
    LocalMux I__8557 (
            .O(N__37091),
            .I(N__37030));
    Span12Mux_s7_v I__8556 (
            .O(N__37088),
            .I(N__37030));
    LocalMux I__8555 (
            .O(N__37085),
            .I(N__37030));
    Span4Mux_s1_h I__8554 (
            .O(N__37080),
            .I(N__37021));
    Span4Mux_v I__8553 (
            .O(N__37077),
            .I(N__37021));
    Span4Mux_v I__8552 (
            .O(N__37074),
            .I(N__37021));
    Span4Mux_v I__8551 (
            .O(N__37069),
            .I(N__37021));
    Odrv4 I__8550 (
            .O(N__37064),
            .I(\ALU.N_240_0 ));
    LocalMux I__8549 (
            .O(N__37059),
            .I(\ALU.N_240_0 ));
    LocalMux I__8548 (
            .O(N__37052),
            .I(\ALU.N_240_0 ));
    Odrv4 I__8547 (
            .O(N__37049),
            .I(\ALU.N_240_0 ));
    LocalMux I__8546 (
            .O(N__37044),
            .I(\ALU.N_240_0 ));
    LocalMux I__8545 (
            .O(N__37037),
            .I(\ALU.N_240_0 ));
    Odrv12 I__8544 (
            .O(N__37030),
            .I(\ALU.N_240_0 ));
    Odrv4 I__8543 (
            .O(N__37021),
            .I(\ALU.N_240_0 ));
    CascadeMux I__8542 (
            .O(N__37004),
            .I(N__36990));
    CascadeMux I__8541 (
            .O(N__37003),
            .I(N__36986));
    CascadeMux I__8540 (
            .O(N__37002),
            .I(N__36976));
    CascadeMux I__8539 (
            .O(N__37001),
            .I(N__36973));
    CascadeMux I__8538 (
            .O(N__37000),
            .I(N__36970));
    CascadeMux I__8537 (
            .O(N__36999),
            .I(N__36967));
    CascadeMux I__8536 (
            .O(N__36998),
            .I(N__36959));
    CascadeMux I__8535 (
            .O(N__36997),
            .I(N__36954));
    InMux I__8534 (
            .O(N__36996),
            .I(N__36949));
    InMux I__8533 (
            .O(N__36995),
            .I(N__36946));
    InMux I__8532 (
            .O(N__36994),
            .I(N__36941));
    InMux I__8531 (
            .O(N__36993),
            .I(N__36933));
    InMux I__8530 (
            .O(N__36990),
            .I(N__36930));
    InMux I__8529 (
            .O(N__36989),
            .I(N__36925));
    InMux I__8528 (
            .O(N__36986),
            .I(N__36925));
    InMux I__8527 (
            .O(N__36985),
            .I(N__36922));
    InMux I__8526 (
            .O(N__36984),
            .I(N__36915));
    InMux I__8525 (
            .O(N__36983),
            .I(N__36915));
    InMux I__8524 (
            .O(N__36982),
            .I(N__36915));
    InMux I__8523 (
            .O(N__36981),
            .I(N__36912));
    InMux I__8522 (
            .O(N__36980),
            .I(N__36905));
    InMux I__8521 (
            .O(N__36979),
            .I(N__36905));
    InMux I__8520 (
            .O(N__36976),
            .I(N__36905));
    InMux I__8519 (
            .O(N__36973),
            .I(N__36902));
    InMux I__8518 (
            .O(N__36970),
            .I(N__36897));
    InMux I__8517 (
            .O(N__36967),
            .I(N__36897));
    InMux I__8516 (
            .O(N__36966),
            .I(N__36890));
    InMux I__8515 (
            .O(N__36965),
            .I(N__36890));
    InMux I__8514 (
            .O(N__36964),
            .I(N__36890));
    InMux I__8513 (
            .O(N__36963),
            .I(N__36887));
    InMux I__8512 (
            .O(N__36962),
            .I(N__36884));
    InMux I__8511 (
            .O(N__36959),
            .I(N__36879));
    InMux I__8510 (
            .O(N__36958),
            .I(N__36879));
    InMux I__8509 (
            .O(N__36957),
            .I(N__36875));
    InMux I__8508 (
            .O(N__36954),
            .I(N__36868));
    InMux I__8507 (
            .O(N__36953),
            .I(N__36868));
    InMux I__8506 (
            .O(N__36952),
            .I(N__36868));
    LocalMux I__8505 (
            .O(N__36949),
            .I(N__36865));
    LocalMux I__8504 (
            .O(N__36946),
            .I(N__36862));
    CascadeMux I__8503 (
            .O(N__36945),
            .I(N__36858));
    CascadeMux I__8502 (
            .O(N__36944),
            .I(N__36855));
    LocalMux I__8501 (
            .O(N__36941),
            .I(N__36852));
    InMux I__8500 (
            .O(N__36940),
            .I(N__36845));
    InMux I__8499 (
            .O(N__36939),
            .I(N__36845));
    InMux I__8498 (
            .O(N__36938),
            .I(N__36845));
    InMux I__8497 (
            .O(N__36937),
            .I(N__36839));
    InMux I__8496 (
            .O(N__36936),
            .I(N__36839));
    LocalMux I__8495 (
            .O(N__36933),
            .I(N__36836));
    LocalMux I__8494 (
            .O(N__36930),
            .I(N__36833));
    LocalMux I__8493 (
            .O(N__36925),
            .I(N__36828));
    LocalMux I__8492 (
            .O(N__36922),
            .I(N__36828));
    LocalMux I__8491 (
            .O(N__36915),
            .I(N__36825));
    LocalMux I__8490 (
            .O(N__36912),
            .I(N__36820));
    LocalMux I__8489 (
            .O(N__36905),
            .I(N__36820));
    LocalMux I__8488 (
            .O(N__36902),
            .I(N__36817));
    LocalMux I__8487 (
            .O(N__36897),
            .I(N__36814));
    LocalMux I__8486 (
            .O(N__36890),
            .I(N__36804));
    LocalMux I__8485 (
            .O(N__36887),
            .I(N__36804));
    LocalMux I__8484 (
            .O(N__36884),
            .I(N__36804));
    LocalMux I__8483 (
            .O(N__36879),
            .I(N__36804));
    InMux I__8482 (
            .O(N__36878),
            .I(N__36801));
    LocalMux I__8481 (
            .O(N__36875),
            .I(N__36796));
    LocalMux I__8480 (
            .O(N__36868),
            .I(N__36796));
    Span4Mux_v I__8479 (
            .O(N__36865),
            .I(N__36791));
    Span4Mux_v I__8478 (
            .O(N__36862),
            .I(N__36791));
    InMux I__8477 (
            .O(N__36861),
            .I(N__36784));
    InMux I__8476 (
            .O(N__36858),
            .I(N__36784));
    InMux I__8475 (
            .O(N__36855),
            .I(N__36784));
    Span4Mux_s2_h I__8474 (
            .O(N__36852),
            .I(N__36779));
    LocalMux I__8473 (
            .O(N__36845),
            .I(N__36779));
    InMux I__8472 (
            .O(N__36844),
            .I(N__36776));
    LocalMux I__8471 (
            .O(N__36839),
            .I(N__36773));
    Span4Mux_h I__8470 (
            .O(N__36836),
            .I(N__36770));
    Span4Mux_v I__8469 (
            .O(N__36833),
            .I(N__36765));
    Span4Mux_v I__8468 (
            .O(N__36828),
            .I(N__36765));
    Span4Mux_h I__8467 (
            .O(N__36825),
            .I(N__36760));
    Span4Mux_v I__8466 (
            .O(N__36820),
            .I(N__36760));
    Span4Mux_h I__8465 (
            .O(N__36817),
            .I(N__36757));
    Span4Mux_v I__8464 (
            .O(N__36814),
            .I(N__36754));
    InMux I__8463 (
            .O(N__36813),
            .I(N__36751));
    Span4Mux_v I__8462 (
            .O(N__36804),
            .I(N__36748));
    LocalMux I__8461 (
            .O(N__36801),
            .I(N__36741));
    Span4Mux_v I__8460 (
            .O(N__36796),
            .I(N__36741));
    Span4Mux_h I__8459 (
            .O(N__36791),
            .I(N__36741));
    LocalMux I__8458 (
            .O(N__36784),
            .I(N__36734));
    Span4Mux_h I__8457 (
            .O(N__36779),
            .I(N__36734));
    LocalMux I__8456 (
            .O(N__36776),
            .I(N__36734));
    Span12Mux_s3_v I__8455 (
            .O(N__36773),
            .I(N__36731));
    Span4Mux_v I__8454 (
            .O(N__36770),
            .I(N__36728));
    Span4Mux_h I__8453 (
            .O(N__36765),
            .I(N__36725));
    Span4Mux_h I__8452 (
            .O(N__36760),
            .I(N__36722));
    Span4Mux_v I__8451 (
            .O(N__36757),
            .I(N__36709));
    Span4Mux_h I__8450 (
            .O(N__36754),
            .I(N__36709));
    LocalMux I__8449 (
            .O(N__36751),
            .I(N__36709));
    Span4Mux_h I__8448 (
            .O(N__36748),
            .I(N__36709));
    Span4Mux_v I__8447 (
            .O(N__36741),
            .I(N__36709));
    Span4Mux_v I__8446 (
            .O(N__36734),
            .I(N__36709));
    Odrv12 I__8445 (
            .O(N__36731),
            .I(\ALU.aluOut_2 ));
    Odrv4 I__8444 (
            .O(N__36728),
            .I(\ALU.aluOut_2 ));
    Odrv4 I__8443 (
            .O(N__36725),
            .I(\ALU.aluOut_2 ));
    Odrv4 I__8442 (
            .O(N__36722),
            .I(\ALU.aluOut_2 ));
    Odrv4 I__8441 (
            .O(N__36709),
            .I(\ALU.aluOut_2 ));
    InMux I__8440 (
            .O(N__36698),
            .I(\ALU.un9_addsub_cry_1 ));
    CascadeMux I__8439 (
            .O(N__36695),
            .I(N__36692));
    InMux I__8438 (
            .O(N__36692),
            .I(N__36689));
    LocalMux I__8437 (
            .O(N__36689),
            .I(N__36686));
    Span12Mux_h I__8436 (
            .O(N__36686),
            .I(N__36683));
    Odrv12 I__8435 (
            .O(N__36683),
            .I(\ALU.N_237_0_i ));
    InMux I__8434 (
            .O(N__36680),
            .I(\ALU.un9_addsub_cry_2 ));
    CascadeMux I__8433 (
            .O(N__36677),
            .I(N__36674));
    InMux I__8432 (
            .O(N__36674),
            .I(N__36671));
    LocalMux I__8431 (
            .O(N__36671),
            .I(N__36668));
    Odrv12 I__8430 (
            .O(N__36668),
            .I(\ALU.N_231_0_i ));
    InMux I__8429 (
            .O(N__36665),
            .I(\ALU.un9_addsub_cry_3 ));
    CascadeMux I__8428 (
            .O(N__36662),
            .I(N__36659));
    InMux I__8427 (
            .O(N__36659),
            .I(N__36656));
    LocalMux I__8426 (
            .O(N__36656),
            .I(N__36653));
    Span4Mux_h I__8425 (
            .O(N__36653),
            .I(N__36650));
    Odrv4 I__8424 (
            .O(N__36650),
            .I(\ALU.madd_axb_0_l_ofx ));
    CascadeMux I__8423 (
            .O(N__36647),
            .I(\ALU.mult_1_cascade_ ));
    InMux I__8422 (
            .O(N__36644),
            .I(N__36641));
    LocalMux I__8421 (
            .O(N__36641),
            .I(N__36638));
    Span4Mux_v I__8420 (
            .O(N__36638),
            .I(N__36635));
    Span4Mux_h I__8419 (
            .O(N__36635),
            .I(N__36632));
    Span4Mux_v I__8418 (
            .O(N__36632),
            .I(N__36629));
    Odrv4 I__8417 (
            .O(N__36629),
            .I(\ALU.a_15_m5_1 ));
    CascadeMux I__8416 (
            .O(N__36626),
            .I(\ALU.d_RNIEICQ63Z0Z_1_cascade_ ));
    InMux I__8415 (
            .O(N__36623),
            .I(N__36617));
    InMux I__8414 (
            .O(N__36622),
            .I(N__36617));
    LocalMux I__8413 (
            .O(N__36617),
            .I(\ALU.bZ0Z_1 ));
    InMux I__8412 (
            .O(N__36614),
            .I(N__36610));
    InMux I__8411 (
            .O(N__36613),
            .I(N__36607));
    LocalMux I__8410 (
            .O(N__36610),
            .I(N__36602));
    LocalMux I__8409 (
            .O(N__36607),
            .I(N__36599));
    InMux I__8408 (
            .O(N__36606),
            .I(N__36596));
    InMux I__8407 (
            .O(N__36605),
            .I(N__36593));
    Span4Mux_h I__8406 (
            .O(N__36602),
            .I(N__36587));
    Span4Mux_h I__8405 (
            .O(N__36599),
            .I(N__36584));
    LocalMux I__8404 (
            .O(N__36596),
            .I(N__36581));
    LocalMux I__8403 (
            .O(N__36593),
            .I(N__36578));
    InMux I__8402 (
            .O(N__36592),
            .I(N__36575));
    InMux I__8401 (
            .O(N__36591),
            .I(N__36572));
    InMux I__8400 (
            .O(N__36590),
            .I(N__36569));
    Odrv4 I__8399 (
            .O(N__36587),
            .I(\ALU.d_RNIEICQ63Z0Z_1 ));
    Odrv4 I__8398 (
            .O(N__36584),
            .I(\ALU.d_RNIEICQ63Z0Z_1 ));
    Odrv4 I__8397 (
            .O(N__36581),
            .I(\ALU.d_RNIEICQ63Z0Z_1 ));
    Odrv12 I__8396 (
            .O(N__36578),
            .I(\ALU.d_RNIEICQ63Z0Z_1 ));
    LocalMux I__8395 (
            .O(N__36575),
            .I(\ALU.d_RNIEICQ63Z0Z_1 ));
    LocalMux I__8394 (
            .O(N__36572),
            .I(\ALU.d_RNIEICQ63Z0Z_1 ));
    LocalMux I__8393 (
            .O(N__36569),
            .I(\ALU.d_RNIEICQ63Z0Z_1 ));
    InMux I__8392 (
            .O(N__36554),
            .I(N__36548));
    InMux I__8391 (
            .O(N__36553),
            .I(N__36548));
    LocalMux I__8390 (
            .O(N__36548),
            .I(N__36545));
    Odrv4 I__8389 (
            .O(N__36545),
            .I(\ALU.dZ0Z_1 ));
    InMux I__8388 (
            .O(N__36542),
            .I(N__36539));
    LocalMux I__8387 (
            .O(N__36539),
            .I(N__36536));
    Span4Mux_h I__8386 (
            .O(N__36536),
            .I(N__36532));
    InMux I__8385 (
            .O(N__36535),
            .I(N__36529));
    Span4Mux_h I__8384 (
            .O(N__36532),
            .I(N__36526));
    LocalMux I__8383 (
            .O(N__36529),
            .I(N__36523));
    Odrv4 I__8382 (
            .O(N__36526),
            .I(\ALU.hZ0Z_4 ));
    Odrv12 I__8381 (
            .O(N__36523),
            .I(\ALU.hZ0Z_4 ));
    InMux I__8380 (
            .O(N__36518),
            .I(N__36514));
    InMux I__8379 (
            .O(N__36517),
            .I(N__36511));
    LocalMux I__8378 (
            .O(N__36514),
            .I(\FTDI.un3_TX_0_i ));
    LocalMux I__8377 (
            .O(N__36511),
            .I(\FTDI.un3_TX_0_i ));
    InMux I__8376 (
            .O(N__36506),
            .I(N__36503));
    LocalMux I__8375 (
            .O(N__36503),
            .I(\FTDI.un3_TX_axb_3 ));
    InMux I__8374 (
            .O(N__36500),
            .I(N__36497));
    LocalMux I__8373 (
            .O(N__36497),
            .I(N__36494));
    Span4Mux_s2_v I__8372 (
            .O(N__36494),
            .I(N__36491));
    Odrv4 I__8371 (
            .O(N__36491),
            .I(\FTDI.TXshiftZ0Z_0 ));
    InMux I__8370 (
            .O(N__36488),
            .I(\FTDI.un3_TX_cry_3 ));
    IoInMux I__8369 (
            .O(N__36485),
            .I(N__36482));
    LocalMux I__8368 (
            .O(N__36482),
            .I(N__36479));
    Span4Mux_s1_v I__8367 (
            .O(N__36479),
            .I(N__36476));
    Span4Mux_h I__8366 (
            .O(N__36476),
            .I(N__36473));
    Span4Mux_h I__8365 (
            .O(N__36473),
            .I(N__36470));
    Odrv4 I__8364 (
            .O(N__36470),
            .I(FTDI_TX_0_i));
    InMux I__8363 (
            .O(N__36467),
            .I(N__36461));
    InMux I__8362 (
            .O(N__36466),
            .I(N__36461));
    LocalMux I__8361 (
            .O(N__36461),
            .I(\ALU.fZ0Z_1 ));
    InMux I__8360 (
            .O(N__36458),
            .I(N__36455));
    LocalMux I__8359 (
            .O(N__36455),
            .I(N__36452));
    Span4Mux_h I__8358 (
            .O(N__36452),
            .I(N__36448));
    InMux I__8357 (
            .O(N__36451),
            .I(N__36445));
    Odrv4 I__8356 (
            .O(N__36448),
            .I(\ALU.fZ0Z_2 ));
    LocalMux I__8355 (
            .O(N__36445),
            .I(\ALU.fZ0Z_2 ));
    CascadeMux I__8354 (
            .O(N__36440),
            .I(N__36437));
    InMux I__8353 (
            .O(N__36437),
            .I(N__36434));
    LocalMux I__8352 (
            .O(N__36434),
            .I(N__36430));
    InMux I__8351 (
            .O(N__36433),
            .I(N__36427));
    Span4Mux_h I__8350 (
            .O(N__36430),
            .I(N__36424));
    LocalMux I__8349 (
            .O(N__36427),
            .I(\ALU.fZ0Z_5 ));
    Odrv4 I__8348 (
            .O(N__36424),
            .I(\ALU.fZ0Z_5 ));
    InMux I__8347 (
            .O(N__36419),
            .I(N__36416));
    LocalMux I__8346 (
            .O(N__36416),
            .I(N__36412));
    InMux I__8345 (
            .O(N__36415),
            .I(N__36409));
    Span4Mux_h I__8344 (
            .O(N__36412),
            .I(N__36406));
    LocalMux I__8343 (
            .O(N__36409),
            .I(N__36403));
    Span4Mux_h I__8342 (
            .O(N__36406),
            .I(N__36400));
    Odrv4 I__8341 (
            .O(N__36403),
            .I(\ALU.fZ0Z_6 ));
    Odrv4 I__8340 (
            .O(N__36400),
            .I(\ALU.fZ0Z_6 ));
    CascadeMux I__8339 (
            .O(N__36395),
            .I(N__36392));
    InMux I__8338 (
            .O(N__36392),
            .I(N__36386));
    InMux I__8337 (
            .O(N__36391),
            .I(N__36386));
    LocalMux I__8336 (
            .O(N__36386),
            .I(N__36383));
    Odrv4 I__8335 (
            .O(N__36383),
            .I(\ALU.fZ0Z_7 ));
    CEMux I__8334 (
            .O(N__36380),
            .I(N__36377));
    LocalMux I__8333 (
            .O(N__36377),
            .I(N__36373));
    CEMux I__8332 (
            .O(N__36376),
            .I(N__36370));
    Span4Mux_v I__8331 (
            .O(N__36373),
            .I(N__36367));
    LocalMux I__8330 (
            .O(N__36370),
            .I(N__36364));
    Span4Mux_v I__8329 (
            .O(N__36367),
            .I(N__36360));
    Span4Mux_v I__8328 (
            .O(N__36364),
            .I(N__36357));
    CEMux I__8327 (
            .O(N__36363),
            .I(N__36354));
    Span4Mux_h I__8326 (
            .O(N__36360),
            .I(N__36351));
    Span4Mux_v I__8325 (
            .O(N__36357),
            .I(N__36348));
    LocalMux I__8324 (
            .O(N__36354),
            .I(N__36345));
    Span4Mux_h I__8323 (
            .O(N__36351),
            .I(N__36342));
    Sp12to4 I__8322 (
            .O(N__36348),
            .I(N__36339));
    Span4Mux_h I__8321 (
            .O(N__36345),
            .I(N__36336));
    Odrv4 I__8320 (
            .O(N__36342),
            .I(\ALU.f_cnvZ0Z_0 ));
    Odrv12 I__8319 (
            .O(N__36339),
            .I(\ALU.f_cnvZ0Z_0 ));
    Odrv4 I__8318 (
            .O(N__36336),
            .I(\ALU.f_cnvZ0Z_0 ));
    InMux I__8317 (
            .O(N__36329),
            .I(N__36326));
    LocalMux I__8316 (
            .O(N__36326),
            .I(N__36322));
    CascadeMux I__8315 (
            .O(N__36325),
            .I(N__36319));
    Span4Mux_h I__8314 (
            .O(N__36322),
            .I(N__36316));
    InMux I__8313 (
            .O(N__36319),
            .I(N__36313));
    Span4Mux_v I__8312 (
            .O(N__36316),
            .I(N__36308));
    LocalMux I__8311 (
            .O(N__36313),
            .I(N__36308));
    Span4Mux_h I__8310 (
            .O(N__36308),
            .I(N__36305));
    Odrv4 I__8309 (
            .O(N__36305),
            .I(\ALU.N_1700_i ));
    CascadeMux I__8308 (
            .O(N__36302),
            .I(\ALU.d_RNIO75MAZ0Z_0_cascade_ ));
    CascadeMux I__8307 (
            .O(N__36299),
            .I(N__36296));
    InMux I__8306 (
            .O(N__36296),
            .I(N__36293));
    LocalMux I__8305 (
            .O(N__36293),
            .I(N__36290));
    Span4Mux_h I__8304 (
            .O(N__36290),
            .I(N__36287));
    Span4Mux_h I__8303 (
            .O(N__36287),
            .I(N__36283));
    InMux I__8302 (
            .O(N__36286),
            .I(N__36280));
    Odrv4 I__8301 (
            .O(N__36283),
            .I(\ALU.bZ0Z_0 ));
    LocalMux I__8300 (
            .O(N__36280),
            .I(\ALU.bZ0Z_0 ));
    InMux I__8299 (
            .O(N__36275),
            .I(N__36272));
    LocalMux I__8298 (
            .O(N__36272),
            .I(N__36269));
    Span4Mux_v I__8297 (
            .O(N__36269),
            .I(N__36265));
    InMux I__8296 (
            .O(N__36268),
            .I(N__36261));
    Span4Mux_h I__8295 (
            .O(N__36265),
            .I(N__36254));
    InMux I__8294 (
            .O(N__36264),
            .I(N__36251));
    LocalMux I__8293 (
            .O(N__36261),
            .I(N__36248));
    InMux I__8292 (
            .O(N__36260),
            .I(N__36245));
    InMux I__8291 (
            .O(N__36259),
            .I(N__36242));
    InMux I__8290 (
            .O(N__36258),
            .I(N__36239));
    InMux I__8289 (
            .O(N__36257),
            .I(N__36236));
    Span4Mux_v I__8288 (
            .O(N__36254),
            .I(N__36231));
    LocalMux I__8287 (
            .O(N__36251),
            .I(N__36231));
    Span4Mux_h I__8286 (
            .O(N__36248),
            .I(N__36228));
    LocalMux I__8285 (
            .O(N__36245),
            .I(N__36223));
    LocalMux I__8284 (
            .O(N__36242),
            .I(N__36223));
    LocalMux I__8283 (
            .O(N__36239),
            .I(N__36218));
    LocalMux I__8282 (
            .O(N__36236),
            .I(N__36218));
    Odrv4 I__8281 (
            .O(N__36231),
            .I(\ALU.a_15_ns_1_9 ));
    Odrv4 I__8280 (
            .O(N__36228),
            .I(\ALU.a_15_ns_1_9 ));
    Odrv4 I__8279 (
            .O(N__36223),
            .I(\ALU.a_15_ns_1_9 ));
    Odrv4 I__8278 (
            .O(N__36218),
            .I(\ALU.a_15_ns_1_9 ));
    CascadeMux I__8277 (
            .O(N__36209),
            .I(N__36206));
    InMux I__8276 (
            .O(N__36206),
            .I(N__36199));
    InMux I__8275 (
            .O(N__36205),
            .I(N__36196));
    InMux I__8274 (
            .O(N__36204),
            .I(N__36191));
    InMux I__8273 (
            .O(N__36203),
            .I(N__36188));
    CascadeMux I__8272 (
            .O(N__36202),
            .I(N__36185));
    LocalMux I__8271 (
            .O(N__36199),
            .I(N__36182));
    LocalMux I__8270 (
            .O(N__36196),
            .I(N__36179));
    InMux I__8269 (
            .O(N__36195),
            .I(N__36175));
    InMux I__8268 (
            .O(N__36194),
            .I(N__36172));
    LocalMux I__8267 (
            .O(N__36191),
            .I(N__36167));
    LocalMux I__8266 (
            .O(N__36188),
            .I(N__36167));
    InMux I__8265 (
            .O(N__36185),
            .I(N__36164));
    Span4Mux_v I__8264 (
            .O(N__36182),
            .I(N__36161));
    Span4Mux_v I__8263 (
            .O(N__36179),
            .I(N__36158));
    InMux I__8262 (
            .O(N__36178),
            .I(N__36155));
    LocalMux I__8261 (
            .O(N__36175),
            .I(N__36152));
    LocalMux I__8260 (
            .O(N__36172),
            .I(N__36147));
    Span4Mux_h I__8259 (
            .O(N__36167),
            .I(N__36147));
    LocalMux I__8258 (
            .O(N__36164),
            .I(N__36140));
    Span4Mux_h I__8257 (
            .O(N__36161),
            .I(N__36140));
    Span4Mux_v I__8256 (
            .O(N__36158),
            .I(N__36140));
    LocalMux I__8255 (
            .O(N__36155),
            .I(\ALU.mult_9 ));
    Odrv4 I__8254 (
            .O(N__36152),
            .I(\ALU.mult_9 ));
    Odrv4 I__8253 (
            .O(N__36147),
            .I(\ALU.mult_9 ));
    Odrv4 I__8252 (
            .O(N__36140),
            .I(\ALU.mult_9 ));
    InMux I__8251 (
            .O(N__36131),
            .I(N__36128));
    LocalMux I__8250 (
            .O(N__36128),
            .I(N__36125));
    Span4Mux_h I__8249 (
            .O(N__36125),
            .I(N__36120));
    InMux I__8248 (
            .O(N__36124),
            .I(N__36115));
    InMux I__8247 (
            .O(N__36123),
            .I(N__36115));
    Span4Mux_h I__8246 (
            .O(N__36120),
            .I(N__36112));
    LocalMux I__8245 (
            .O(N__36115),
            .I(N__36109));
    Odrv4 I__8244 (
            .O(N__36112),
            .I(\ALU.gZ0Z_9 ));
    Odrv12 I__8243 (
            .O(N__36109),
            .I(\ALU.gZ0Z_9 ));
    CEMux I__8242 (
            .O(N__36104),
            .I(N__36101));
    LocalMux I__8241 (
            .O(N__36101),
            .I(N__36097));
    CEMux I__8240 (
            .O(N__36100),
            .I(N__36094));
    Span4Mux_v I__8239 (
            .O(N__36097),
            .I(N__36090));
    LocalMux I__8238 (
            .O(N__36094),
            .I(N__36087));
    CEMux I__8237 (
            .O(N__36093),
            .I(N__36084));
    Span4Mux_v I__8236 (
            .O(N__36090),
            .I(N__36081));
    Span4Mux_v I__8235 (
            .O(N__36087),
            .I(N__36076));
    LocalMux I__8234 (
            .O(N__36084),
            .I(N__36076));
    Span4Mux_h I__8233 (
            .O(N__36081),
            .I(N__36073));
    Span4Mux_h I__8232 (
            .O(N__36076),
            .I(N__36070));
    Span4Mux_v I__8231 (
            .O(N__36073),
            .I(N__36066));
    Span4Mux_h I__8230 (
            .O(N__36070),
            .I(N__36063));
    CEMux I__8229 (
            .O(N__36069),
            .I(N__36060));
    Span4Mux_v I__8228 (
            .O(N__36066),
            .I(N__36057));
    Sp12to4 I__8227 (
            .O(N__36063),
            .I(N__36054));
    LocalMux I__8226 (
            .O(N__36060),
            .I(N__36051));
    Sp12to4 I__8225 (
            .O(N__36057),
            .I(N__36046));
    Span12Mux_v I__8224 (
            .O(N__36054),
            .I(N__36046));
    Span4Mux_v I__8223 (
            .O(N__36051),
            .I(N__36043));
    Odrv12 I__8222 (
            .O(N__36046),
            .I(\ALU.g_cnvZ0Z_0 ));
    Odrv4 I__8221 (
            .O(N__36043),
            .I(\ALU.g_cnvZ0Z_0 ));
    InMux I__8220 (
            .O(N__36038),
            .I(N__36035));
    LocalMux I__8219 (
            .O(N__36035),
            .I(N__36032));
    Span4Mux_h I__8218 (
            .O(N__36032),
            .I(N__36028));
    InMux I__8217 (
            .O(N__36031),
            .I(N__36025));
    Odrv4 I__8216 (
            .O(N__36028),
            .I(\ALU.eZ0Z_13 ));
    LocalMux I__8215 (
            .O(N__36025),
            .I(\ALU.eZ0Z_13 ));
    InMux I__8214 (
            .O(N__36020),
            .I(N__36016));
    InMux I__8213 (
            .O(N__36019),
            .I(N__36013));
    LocalMux I__8212 (
            .O(N__36016),
            .I(N__36010));
    LocalMux I__8211 (
            .O(N__36013),
            .I(\ALU.aZ0Z_13 ));
    Odrv4 I__8210 (
            .O(N__36010),
            .I(\ALU.aZ0Z_13 ));
    CascadeMux I__8209 (
            .O(N__36005),
            .I(N__36000));
    CascadeMux I__8208 (
            .O(N__36004),
            .I(N__35997));
    CascadeMux I__8207 (
            .O(N__36003),
            .I(N__35993));
    InMux I__8206 (
            .O(N__36000),
            .I(N__35990));
    InMux I__8205 (
            .O(N__35997),
            .I(N__35986));
    InMux I__8204 (
            .O(N__35996),
            .I(N__35982));
    InMux I__8203 (
            .O(N__35993),
            .I(N__35979));
    LocalMux I__8202 (
            .O(N__35990),
            .I(N__35976));
    InMux I__8201 (
            .O(N__35989),
            .I(N__35973));
    LocalMux I__8200 (
            .O(N__35986),
            .I(N__35970));
    CascadeMux I__8199 (
            .O(N__35985),
            .I(N__35967));
    LocalMux I__8198 (
            .O(N__35982),
            .I(N__35962));
    LocalMux I__8197 (
            .O(N__35979),
            .I(N__35959));
    Span4Mux_v I__8196 (
            .O(N__35976),
            .I(N__35954));
    LocalMux I__8195 (
            .O(N__35973),
            .I(N__35954));
    Span4Mux_v I__8194 (
            .O(N__35970),
            .I(N__35951));
    InMux I__8193 (
            .O(N__35967),
            .I(N__35948));
    CascadeMux I__8192 (
            .O(N__35966),
            .I(N__35945));
    CascadeMux I__8191 (
            .O(N__35965),
            .I(N__35942));
    Span4Mux_v I__8190 (
            .O(N__35962),
            .I(N__35937));
    Span4Mux_v I__8189 (
            .O(N__35959),
            .I(N__35937));
    Span4Mux_h I__8188 (
            .O(N__35954),
            .I(N__35934));
    Span4Mux_h I__8187 (
            .O(N__35951),
            .I(N__35931));
    LocalMux I__8186 (
            .O(N__35948),
            .I(N__35928));
    InMux I__8185 (
            .O(N__35945),
            .I(N__35923));
    InMux I__8184 (
            .O(N__35942),
            .I(N__35923));
    Odrv4 I__8183 (
            .O(N__35937),
            .I(aluOperand1_2_rep2));
    Odrv4 I__8182 (
            .O(N__35934),
            .I(aluOperand1_2_rep2));
    Odrv4 I__8181 (
            .O(N__35931),
            .I(aluOperand1_2_rep2));
    Odrv12 I__8180 (
            .O(N__35928),
            .I(aluOperand1_2_rep2));
    LocalMux I__8179 (
            .O(N__35923),
            .I(aluOperand1_2_rep2));
    InMux I__8178 (
            .O(N__35912),
            .I(N__35907));
    CascadeMux I__8177 (
            .O(N__35911),
            .I(N__35903));
    InMux I__8176 (
            .O(N__35910),
            .I(N__35900));
    LocalMux I__8175 (
            .O(N__35907),
            .I(N__35894));
    InMux I__8174 (
            .O(N__35906),
            .I(N__35889));
    InMux I__8173 (
            .O(N__35903),
            .I(N__35889));
    LocalMux I__8172 (
            .O(N__35900),
            .I(N__35886));
    InMux I__8171 (
            .O(N__35899),
            .I(N__35883));
    InMux I__8170 (
            .O(N__35898),
            .I(N__35880));
    InMux I__8169 (
            .O(N__35897),
            .I(N__35877));
    Span4Mux_h I__8168 (
            .O(N__35894),
            .I(N__35872));
    LocalMux I__8167 (
            .O(N__35889),
            .I(N__35863));
    Span4Mux_v I__8166 (
            .O(N__35886),
            .I(N__35863));
    LocalMux I__8165 (
            .O(N__35883),
            .I(N__35863));
    LocalMux I__8164 (
            .O(N__35880),
            .I(N__35860));
    LocalMux I__8163 (
            .O(N__35877),
            .I(N__35857));
    InMux I__8162 (
            .O(N__35876),
            .I(N__35854));
    CascadeMux I__8161 (
            .O(N__35875),
            .I(N__35849));
    Span4Mux_v I__8160 (
            .O(N__35872),
            .I(N__35846));
    InMux I__8159 (
            .O(N__35871),
            .I(N__35841));
    InMux I__8158 (
            .O(N__35870),
            .I(N__35841));
    Span4Mux_h I__8157 (
            .O(N__35863),
            .I(N__35838));
    Span4Mux_h I__8156 (
            .O(N__35860),
            .I(N__35833));
    Span4Mux_h I__8155 (
            .O(N__35857),
            .I(N__35833));
    LocalMux I__8154 (
            .O(N__35854),
            .I(N__35830));
    InMux I__8153 (
            .O(N__35853),
            .I(N__35823));
    InMux I__8152 (
            .O(N__35852),
            .I(N__35823));
    InMux I__8151 (
            .O(N__35849),
            .I(N__35823));
    Odrv4 I__8150 (
            .O(N__35846),
            .I(aluOperand1_1_rep1));
    LocalMux I__8149 (
            .O(N__35841),
            .I(aluOperand1_1_rep1));
    Odrv4 I__8148 (
            .O(N__35838),
            .I(aluOperand1_1_rep1));
    Odrv4 I__8147 (
            .O(N__35833),
            .I(aluOperand1_1_rep1));
    Odrv12 I__8146 (
            .O(N__35830),
            .I(aluOperand1_1_rep1));
    LocalMux I__8145 (
            .O(N__35823),
            .I(aluOperand1_1_rep1));
    InMux I__8144 (
            .O(N__35810),
            .I(N__35806));
    InMux I__8143 (
            .O(N__35809),
            .I(N__35803));
    LocalMux I__8142 (
            .O(N__35806),
            .I(\ALU.cZ0Z_13 ));
    LocalMux I__8141 (
            .O(N__35803),
            .I(\ALU.cZ0Z_13 ));
    CascadeMux I__8140 (
            .O(N__35798),
            .I(\ALU.dout_3_ns_1_13_cascade_ ));
    InMux I__8139 (
            .O(N__35795),
            .I(N__35791));
    InMux I__8138 (
            .O(N__35794),
            .I(N__35788));
    LocalMux I__8137 (
            .O(N__35791),
            .I(\ALU.gZ0Z_13 ));
    LocalMux I__8136 (
            .O(N__35788),
            .I(\ALU.gZ0Z_13 ));
    InMux I__8135 (
            .O(N__35783),
            .I(N__35776));
    InMux I__8134 (
            .O(N__35782),
            .I(N__35776));
    InMux I__8133 (
            .O(N__35781),
            .I(N__35773));
    LocalMux I__8132 (
            .O(N__35776),
            .I(N__35770));
    LocalMux I__8131 (
            .O(N__35773),
            .I(N__35767));
    Odrv4 I__8130 (
            .O(N__35770),
            .I(\ALU.bZ0Z_13 ));
    Odrv4 I__8129 (
            .O(N__35767),
            .I(\ALU.bZ0Z_13 ));
    InMux I__8128 (
            .O(N__35762),
            .I(N__35758));
    InMux I__8127 (
            .O(N__35761),
            .I(N__35755));
    LocalMux I__8126 (
            .O(N__35758),
            .I(N__35749));
    LocalMux I__8125 (
            .O(N__35755),
            .I(N__35745));
    CascadeMux I__8124 (
            .O(N__35754),
            .I(N__35742));
    CascadeMux I__8123 (
            .O(N__35753),
            .I(N__35739));
    InMux I__8122 (
            .O(N__35752),
            .I(N__35734));
    Span4Mux_h I__8121 (
            .O(N__35749),
            .I(N__35731));
    InMux I__8120 (
            .O(N__35748),
            .I(N__35728));
    Span4Mux_h I__8119 (
            .O(N__35745),
            .I(N__35725));
    InMux I__8118 (
            .O(N__35742),
            .I(N__35720));
    InMux I__8117 (
            .O(N__35739),
            .I(N__35720));
    CascadeMux I__8116 (
            .O(N__35738),
            .I(N__35717));
    InMux I__8115 (
            .O(N__35737),
            .I(N__35714));
    LocalMux I__8114 (
            .O(N__35734),
            .I(N__35710));
    Span4Mux_v I__8113 (
            .O(N__35731),
            .I(N__35703));
    LocalMux I__8112 (
            .O(N__35728),
            .I(N__35700));
    Span4Mux_v I__8111 (
            .O(N__35725),
            .I(N__35695));
    LocalMux I__8110 (
            .O(N__35720),
            .I(N__35692));
    InMux I__8109 (
            .O(N__35717),
            .I(N__35689));
    LocalMux I__8108 (
            .O(N__35714),
            .I(N__35686));
    InMux I__8107 (
            .O(N__35713),
            .I(N__35683));
    Span4Mux_h I__8106 (
            .O(N__35710),
            .I(N__35680));
    InMux I__8105 (
            .O(N__35709),
            .I(N__35677));
    InMux I__8104 (
            .O(N__35708),
            .I(N__35672));
    InMux I__8103 (
            .O(N__35707),
            .I(N__35672));
    InMux I__8102 (
            .O(N__35706),
            .I(N__35668));
    Span4Mux_v I__8101 (
            .O(N__35703),
            .I(N__35663));
    Span4Mux_v I__8100 (
            .O(N__35700),
            .I(N__35663));
    InMux I__8099 (
            .O(N__35699),
            .I(N__35658));
    InMux I__8098 (
            .O(N__35698),
            .I(N__35658));
    Span4Mux_v I__8097 (
            .O(N__35695),
            .I(N__35653));
    Span4Mux_h I__8096 (
            .O(N__35692),
            .I(N__35653));
    LocalMux I__8095 (
            .O(N__35689),
            .I(N__35648));
    Span4Mux_v I__8094 (
            .O(N__35686),
            .I(N__35648));
    LocalMux I__8093 (
            .O(N__35683),
            .I(N__35645));
    Span4Mux_h I__8092 (
            .O(N__35680),
            .I(N__35638));
    LocalMux I__8091 (
            .O(N__35677),
            .I(N__35638));
    LocalMux I__8090 (
            .O(N__35672),
            .I(N__35638));
    InMux I__8089 (
            .O(N__35671),
            .I(N__35635));
    LocalMux I__8088 (
            .O(N__35668),
            .I(N__35632));
    Odrv4 I__8087 (
            .O(N__35663),
            .I(aluOperand1_1_rep2));
    LocalMux I__8086 (
            .O(N__35658),
            .I(aluOperand1_1_rep2));
    Odrv4 I__8085 (
            .O(N__35653),
            .I(aluOperand1_1_rep2));
    Odrv4 I__8084 (
            .O(N__35648),
            .I(aluOperand1_1_rep2));
    Odrv12 I__8083 (
            .O(N__35645),
            .I(aluOperand1_1_rep2));
    Odrv4 I__8082 (
            .O(N__35638),
            .I(aluOperand1_1_rep2));
    LocalMux I__8081 (
            .O(N__35635),
            .I(aluOperand1_1_rep2));
    Odrv4 I__8080 (
            .O(N__35632),
            .I(aluOperand1_1_rep2));
    CascadeMux I__8079 (
            .O(N__35615),
            .I(N__35611));
    CascadeMux I__8078 (
            .O(N__35614),
            .I(N__35608));
    InMux I__8077 (
            .O(N__35611),
            .I(N__35604));
    InMux I__8076 (
            .O(N__35608),
            .I(N__35599));
    InMux I__8075 (
            .O(N__35607),
            .I(N__35599));
    LocalMux I__8074 (
            .O(N__35604),
            .I(N__35596));
    LocalMux I__8073 (
            .O(N__35599),
            .I(N__35591));
    Span4Mux_v I__8072 (
            .O(N__35596),
            .I(N__35591));
    Odrv4 I__8071 (
            .O(N__35591),
            .I(\ALU.fZ0Z_13 ));
    InMux I__8070 (
            .O(N__35588),
            .I(N__35583));
    CascadeMux I__8069 (
            .O(N__35587),
            .I(N__35578));
    CascadeMux I__8068 (
            .O(N__35586),
            .I(N__35573));
    LocalMux I__8067 (
            .O(N__35583),
            .I(N__35570));
    CascadeMux I__8066 (
            .O(N__35582),
            .I(N__35567));
    CascadeMux I__8065 (
            .O(N__35581),
            .I(N__35564));
    InMux I__8064 (
            .O(N__35578),
            .I(N__35561));
    InMux I__8063 (
            .O(N__35577),
            .I(N__35558));
    InMux I__8062 (
            .O(N__35576),
            .I(N__35555));
    InMux I__8061 (
            .O(N__35573),
            .I(N__35551));
    Span4Mux_v I__8060 (
            .O(N__35570),
            .I(N__35548));
    InMux I__8059 (
            .O(N__35567),
            .I(N__35545));
    InMux I__8058 (
            .O(N__35564),
            .I(N__35542));
    LocalMux I__8057 (
            .O(N__35561),
            .I(N__35539));
    LocalMux I__8056 (
            .O(N__35558),
            .I(N__35536));
    LocalMux I__8055 (
            .O(N__35555),
            .I(N__35533));
    CascadeMux I__8054 (
            .O(N__35554),
            .I(N__35528));
    LocalMux I__8053 (
            .O(N__35551),
            .I(N__35525));
    Span4Mux_h I__8052 (
            .O(N__35548),
            .I(N__35522));
    LocalMux I__8051 (
            .O(N__35545),
            .I(N__35519));
    LocalMux I__8050 (
            .O(N__35542),
            .I(N__35516));
    Span4Mux_h I__8049 (
            .O(N__35539),
            .I(N__35513));
    Span4Mux_v I__8048 (
            .O(N__35536),
            .I(N__35510));
    Span4Mux_h I__8047 (
            .O(N__35533),
            .I(N__35507));
    InMux I__8046 (
            .O(N__35532),
            .I(N__35504));
    CascadeMux I__8045 (
            .O(N__35531),
            .I(N__35501));
    InMux I__8044 (
            .O(N__35528),
            .I(N__35498));
    Span4Mux_h I__8043 (
            .O(N__35525),
            .I(N__35495));
    Span4Mux_v I__8042 (
            .O(N__35522),
            .I(N__35488));
    Span4Mux_v I__8041 (
            .O(N__35519),
            .I(N__35488));
    Span4Mux_v I__8040 (
            .O(N__35516),
            .I(N__35488));
    Span4Mux_v I__8039 (
            .O(N__35513),
            .I(N__35483));
    Span4Mux_h I__8038 (
            .O(N__35510),
            .I(N__35483));
    Span4Mux_v I__8037 (
            .O(N__35507),
            .I(N__35478));
    LocalMux I__8036 (
            .O(N__35504),
            .I(N__35478));
    InMux I__8035 (
            .O(N__35501),
            .I(N__35475));
    LocalMux I__8034 (
            .O(N__35498),
            .I(aluOperand1_2));
    Odrv4 I__8033 (
            .O(N__35495),
            .I(aluOperand1_2));
    Odrv4 I__8032 (
            .O(N__35488),
            .I(aluOperand1_2));
    Odrv4 I__8031 (
            .O(N__35483),
            .I(aluOperand1_2));
    Odrv4 I__8030 (
            .O(N__35478),
            .I(aluOperand1_2));
    LocalMux I__8029 (
            .O(N__35475),
            .I(aluOperand1_2));
    InMux I__8028 (
            .O(N__35462),
            .I(N__35458));
    InMux I__8027 (
            .O(N__35461),
            .I(N__35455));
    LocalMux I__8026 (
            .O(N__35458),
            .I(N__35452));
    LocalMux I__8025 (
            .O(N__35455),
            .I(N__35447));
    Span4Mux_v I__8024 (
            .O(N__35452),
            .I(N__35447));
    Span4Mux_h I__8023 (
            .O(N__35447),
            .I(N__35443));
    InMux I__8022 (
            .O(N__35446),
            .I(N__35440));
    Odrv4 I__8021 (
            .O(N__35443),
            .I(\ALU.hZ0Z_13 ));
    LocalMux I__8020 (
            .O(N__35440),
            .I(\ALU.hZ0Z_13 ));
    InMux I__8019 (
            .O(N__35435),
            .I(N__35431));
    InMux I__8018 (
            .O(N__35434),
            .I(N__35428));
    LocalMux I__8017 (
            .O(N__35431),
            .I(N__35425));
    LocalMux I__8016 (
            .O(N__35428),
            .I(N__35421));
    Span4Mux_v I__8015 (
            .O(N__35425),
            .I(N__35418));
    InMux I__8014 (
            .O(N__35424),
            .I(N__35415));
    Span4Mux_h I__8013 (
            .O(N__35421),
            .I(N__35410));
    Span4Mux_h I__8012 (
            .O(N__35418),
            .I(N__35410));
    LocalMux I__8011 (
            .O(N__35415),
            .I(\ALU.dZ0Z_13 ));
    Odrv4 I__8010 (
            .O(N__35410),
            .I(\ALU.dZ0Z_13 ));
    CascadeMux I__8009 (
            .O(N__35405),
            .I(\ALU.dout_6_ns_1_13_cascade_ ));
    InMux I__8008 (
            .O(N__35402),
            .I(N__35396));
    InMux I__8007 (
            .O(N__35401),
            .I(N__35396));
    LocalMux I__8006 (
            .O(N__35396),
            .I(N__35391));
    InMux I__8005 (
            .O(N__35395),
            .I(N__35386));
    InMux I__8004 (
            .O(N__35394),
            .I(N__35386));
    Span4Mux_v I__8003 (
            .O(N__35391),
            .I(N__35379));
    LocalMux I__8002 (
            .O(N__35386),
            .I(N__35379));
    CascadeMux I__8001 (
            .O(N__35385),
            .I(N__35371));
    CascadeMux I__8000 (
            .O(N__35384),
            .I(N__35368));
    Span4Mux_v I__7999 (
            .O(N__35379),
            .I(N__35362));
    InMux I__7998 (
            .O(N__35378),
            .I(N__35357));
    InMux I__7997 (
            .O(N__35377),
            .I(N__35357));
    InMux I__7996 (
            .O(N__35376),
            .I(N__35353));
    InMux I__7995 (
            .O(N__35375),
            .I(N__35347));
    InMux I__7994 (
            .O(N__35374),
            .I(N__35347));
    InMux I__7993 (
            .O(N__35371),
            .I(N__35344));
    InMux I__7992 (
            .O(N__35368),
            .I(N__35341));
    InMux I__7991 (
            .O(N__35367),
            .I(N__35338));
    InMux I__7990 (
            .O(N__35366),
            .I(N__35335));
    CascadeMux I__7989 (
            .O(N__35365),
            .I(N__35332));
    Span4Mux_h I__7988 (
            .O(N__35362),
            .I(N__35329));
    LocalMux I__7987 (
            .O(N__35357),
            .I(N__35326));
    InMux I__7986 (
            .O(N__35356),
            .I(N__35323));
    LocalMux I__7985 (
            .O(N__35353),
            .I(N__35320));
    InMux I__7984 (
            .O(N__35352),
            .I(N__35317));
    LocalMux I__7983 (
            .O(N__35347),
            .I(N__35314));
    LocalMux I__7982 (
            .O(N__35344),
            .I(N__35311));
    LocalMux I__7981 (
            .O(N__35341),
            .I(N__35308));
    LocalMux I__7980 (
            .O(N__35338),
            .I(N__35303));
    LocalMux I__7979 (
            .O(N__35335),
            .I(N__35303));
    InMux I__7978 (
            .O(N__35332),
            .I(N__35300));
    Span4Mux_h I__7977 (
            .O(N__35329),
            .I(N__35294));
    Span4Mux_h I__7976 (
            .O(N__35326),
            .I(N__35289));
    LocalMux I__7975 (
            .O(N__35323),
            .I(N__35289));
    Span4Mux_v I__7974 (
            .O(N__35320),
            .I(N__35280));
    LocalMux I__7973 (
            .O(N__35317),
            .I(N__35280));
    Span4Mux_v I__7972 (
            .O(N__35314),
            .I(N__35280));
    Span4Mux_v I__7971 (
            .O(N__35311),
            .I(N__35280));
    Span4Mux_v I__7970 (
            .O(N__35308),
            .I(N__35275));
    Span4Mux_v I__7969 (
            .O(N__35303),
            .I(N__35275));
    LocalMux I__7968 (
            .O(N__35300),
            .I(N__35272));
    InMux I__7967 (
            .O(N__35299),
            .I(N__35265));
    InMux I__7966 (
            .O(N__35298),
            .I(N__35265));
    InMux I__7965 (
            .O(N__35297),
            .I(N__35265));
    Odrv4 I__7964 (
            .O(N__35294),
            .I(aluOperand1_1));
    Odrv4 I__7963 (
            .O(N__35289),
            .I(aluOperand1_1));
    Odrv4 I__7962 (
            .O(N__35280),
            .I(aluOperand1_1));
    Odrv4 I__7961 (
            .O(N__35275),
            .I(aluOperand1_1));
    Odrv12 I__7960 (
            .O(N__35272),
            .I(aluOperand1_1));
    LocalMux I__7959 (
            .O(N__35265),
            .I(aluOperand1_1));
    InMux I__7958 (
            .O(N__35252),
            .I(N__35249));
    LocalMux I__7957 (
            .O(N__35249),
            .I(\ALU.N_712 ));
    CascadeMux I__7956 (
            .O(N__35246),
            .I(\ALU.N_760_cascade_ ));
    InMux I__7955 (
            .O(N__35243),
            .I(N__35236));
    InMux I__7954 (
            .O(N__35242),
            .I(N__35236));
    InMux I__7953 (
            .O(N__35241),
            .I(N__35233));
    LocalMux I__7952 (
            .O(N__35236),
            .I(N__35226));
    LocalMux I__7951 (
            .O(N__35233),
            .I(N__35217));
    InMux I__7950 (
            .O(N__35232),
            .I(N__35214));
    InMux I__7949 (
            .O(N__35231),
            .I(N__35211));
    InMux I__7948 (
            .O(N__35230),
            .I(N__35208));
    InMux I__7947 (
            .O(N__35229),
            .I(N__35203));
    Span4Mux_v I__7946 (
            .O(N__35226),
            .I(N__35199));
    InMux I__7945 (
            .O(N__35225),
            .I(N__35196));
    InMux I__7944 (
            .O(N__35224),
            .I(N__35193));
    InMux I__7943 (
            .O(N__35223),
            .I(N__35190));
    InMux I__7942 (
            .O(N__35222),
            .I(N__35187));
    InMux I__7941 (
            .O(N__35221),
            .I(N__35184));
    InMux I__7940 (
            .O(N__35220),
            .I(N__35180));
    Span4Mux_v I__7939 (
            .O(N__35217),
            .I(N__35175));
    LocalMux I__7938 (
            .O(N__35214),
            .I(N__35175));
    LocalMux I__7937 (
            .O(N__35211),
            .I(N__35170));
    LocalMux I__7936 (
            .O(N__35208),
            .I(N__35170));
    InMux I__7935 (
            .O(N__35207),
            .I(N__35167));
    InMux I__7934 (
            .O(N__35206),
            .I(N__35164));
    LocalMux I__7933 (
            .O(N__35203),
            .I(N__35161));
    InMux I__7932 (
            .O(N__35202),
            .I(N__35158));
    Span4Mux_v I__7931 (
            .O(N__35199),
            .I(N__35151));
    LocalMux I__7930 (
            .O(N__35196),
            .I(N__35151));
    LocalMux I__7929 (
            .O(N__35193),
            .I(N__35151));
    LocalMux I__7928 (
            .O(N__35190),
            .I(N__35148));
    LocalMux I__7927 (
            .O(N__35187),
            .I(N__35145));
    LocalMux I__7926 (
            .O(N__35184),
            .I(N__35142));
    InMux I__7925 (
            .O(N__35183),
            .I(N__35139));
    LocalMux I__7924 (
            .O(N__35180),
            .I(N__35136));
    Span4Mux_v I__7923 (
            .O(N__35175),
            .I(N__35125));
    Span4Mux_v I__7922 (
            .O(N__35170),
            .I(N__35125));
    LocalMux I__7921 (
            .O(N__35167),
            .I(N__35125));
    LocalMux I__7920 (
            .O(N__35164),
            .I(N__35125));
    Span4Mux_v I__7919 (
            .O(N__35161),
            .I(N__35122));
    LocalMux I__7918 (
            .O(N__35158),
            .I(N__35119));
    Span4Mux_h I__7917 (
            .O(N__35151),
            .I(N__35116));
    Span12Mux_v I__7916 (
            .O(N__35148),
            .I(N__35113));
    Span12Mux_v I__7915 (
            .O(N__35145),
            .I(N__35110));
    Span4Mux_h I__7914 (
            .O(N__35142),
            .I(N__35107));
    LocalMux I__7913 (
            .O(N__35139),
            .I(N__35102));
    Span4Mux_v I__7912 (
            .O(N__35136),
            .I(N__35102));
    InMux I__7911 (
            .O(N__35135),
            .I(N__35097));
    InMux I__7910 (
            .O(N__35134),
            .I(N__35097));
    Span4Mux_h I__7909 (
            .O(N__35125),
            .I(N__35094));
    Span4Mux_h I__7908 (
            .O(N__35122),
            .I(N__35087));
    Span4Mux_v I__7907 (
            .O(N__35119),
            .I(N__35087));
    Span4Mux_v I__7906 (
            .O(N__35116),
            .I(N__35087));
    Odrv12 I__7905 (
            .O(N__35113),
            .I(aluOperand1_0));
    Odrv12 I__7904 (
            .O(N__35110),
            .I(aluOperand1_0));
    Odrv4 I__7903 (
            .O(N__35107),
            .I(aluOperand1_0));
    Odrv4 I__7902 (
            .O(N__35102),
            .I(aluOperand1_0));
    LocalMux I__7901 (
            .O(N__35097),
            .I(aluOperand1_0));
    Odrv4 I__7900 (
            .O(N__35094),
            .I(aluOperand1_0));
    Odrv4 I__7899 (
            .O(N__35087),
            .I(aluOperand1_0));
    CascadeMux I__7898 (
            .O(N__35072),
            .I(\ALU.aluOut_13_cascade_ ));
    CascadeMux I__7897 (
            .O(N__35069),
            .I(N__35066));
    InMux I__7896 (
            .O(N__35066),
            .I(N__35062));
    InMux I__7895 (
            .O(N__35065),
            .I(N__35059));
    LocalMux I__7894 (
            .O(N__35062),
            .I(N__35054));
    LocalMux I__7893 (
            .O(N__35059),
            .I(N__35054));
    Odrv12 I__7892 (
            .O(N__35054),
            .I(\ALU.a13_b_0 ));
    InMux I__7891 (
            .O(N__35051),
            .I(N__35048));
    LocalMux I__7890 (
            .O(N__35048),
            .I(N__35045));
    Span4Mux_h I__7889 (
            .O(N__35045),
            .I(N__35041));
    InMux I__7888 (
            .O(N__35044),
            .I(N__35038));
    Odrv4 I__7887 (
            .O(N__35041),
            .I(\ALU.fZ0Z_0 ));
    LocalMux I__7886 (
            .O(N__35038),
            .I(\ALU.fZ0Z_0 ));
    InMux I__7885 (
            .O(N__35033),
            .I(N__35023));
    InMux I__7884 (
            .O(N__35032),
            .I(N__35020));
    InMux I__7883 (
            .O(N__35031),
            .I(N__35017));
    InMux I__7882 (
            .O(N__35030),
            .I(N__35014));
    InMux I__7881 (
            .O(N__35029),
            .I(N__35009));
    InMux I__7880 (
            .O(N__35028),
            .I(N__35006));
    InMux I__7879 (
            .O(N__35027),
            .I(N__35003));
    InMux I__7878 (
            .O(N__35026),
            .I(N__35000));
    LocalMux I__7877 (
            .O(N__35023),
            .I(N__34995));
    LocalMux I__7876 (
            .O(N__35020),
            .I(N__34995));
    LocalMux I__7875 (
            .O(N__35017),
            .I(N__34988));
    LocalMux I__7874 (
            .O(N__35014),
            .I(N__34988));
    InMux I__7873 (
            .O(N__35013),
            .I(N__34983));
    InMux I__7872 (
            .O(N__35012),
            .I(N__34983));
    LocalMux I__7871 (
            .O(N__35009),
            .I(N__34980));
    LocalMux I__7870 (
            .O(N__35006),
            .I(N__34977));
    LocalMux I__7869 (
            .O(N__35003),
            .I(N__34972));
    LocalMux I__7868 (
            .O(N__35000),
            .I(N__34972));
    Span4Mux_h I__7867 (
            .O(N__34995),
            .I(N__34969));
    InMux I__7866 (
            .O(N__34994),
            .I(N__34966));
    InMux I__7865 (
            .O(N__34993),
            .I(N__34963));
    Span4Mux_v I__7864 (
            .O(N__34988),
            .I(N__34960));
    LocalMux I__7863 (
            .O(N__34983),
            .I(N__34957));
    Span4Mux_h I__7862 (
            .O(N__34980),
            .I(N__34954));
    Span4Mux_h I__7861 (
            .O(N__34977),
            .I(N__34947));
    Span4Mux_h I__7860 (
            .O(N__34972),
            .I(N__34947));
    Span4Mux_v I__7859 (
            .O(N__34969),
            .I(N__34947));
    LocalMux I__7858 (
            .O(N__34966),
            .I(aluOperand2_1_rep1));
    LocalMux I__7857 (
            .O(N__34963),
            .I(aluOperand2_1_rep1));
    Odrv4 I__7856 (
            .O(N__34960),
            .I(aluOperand2_1_rep1));
    Odrv12 I__7855 (
            .O(N__34957),
            .I(aluOperand2_1_rep1));
    Odrv4 I__7854 (
            .O(N__34954),
            .I(aluOperand2_1_rep1));
    Odrv4 I__7853 (
            .O(N__34947),
            .I(aluOperand2_1_rep1));
    InMux I__7852 (
            .O(N__34934),
            .I(N__34930));
    InMux I__7851 (
            .O(N__34933),
            .I(N__34927));
    LocalMux I__7850 (
            .O(N__34930),
            .I(N__34924));
    LocalMux I__7849 (
            .O(N__34927),
            .I(N__34921));
    Span4Mux_h I__7848 (
            .O(N__34924),
            .I(N__34918));
    Span4Mux_h I__7847 (
            .O(N__34921),
            .I(N__34914));
    Span4Mux_h I__7846 (
            .O(N__34918),
            .I(N__34911));
    InMux I__7845 (
            .O(N__34917),
            .I(N__34908));
    Odrv4 I__7844 (
            .O(N__34914),
            .I(\ALU.cZ0Z_10 ));
    Odrv4 I__7843 (
            .O(N__34911),
            .I(\ALU.cZ0Z_10 ));
    LocalMux I__7842 (
            .O(N__34908),
            .I(\ALU.cZ0Z_10 ));
    InMux I__7841 (
            .O(N__34901),
            .I(N__34898));
    LocalMux I__7840 (
            .O(N__34898),
            .I(N__34895));
    Span4Mux_v I__7839 (
            .O(N__34895),
            .I(N__34892));
    Span4Mux_v I__7838 (
            .O(N__34892),
            .I(N__34888));
    InMux I__7837 (
            .O(N__34891),
            .I(N__34885));
    Span4Mux_h I__7836 (
            .O(N__34888),
            .I(N__34877));
    LocalMux I__7835 (
            .O(N__34885),
            .I(N__34877));
    InMux I__7834 (
            .O(N__34884),
            .I(N__34872));
    InMux I__7833 (
            .O(N__34883),
            .I(N__34872));
    InMux I__7832 (
            .O(N__34882),
            .I(N__34869));
    Span4Mux_v I__7831 (
            .O(N__34877),
            .I(N__34864));
    LocalMux I__7830 (
            .O(N__34872),
            .I(N__34859));
    LocalMux I__7829 (
            .O(N__34869),
            .I(N__34856));
    CascadeMux I__7828 (
            .O(N__34868),
            .I(N__34851));
    InMux I__7827 (
            .O(N__34867),
            .I(N__34848));
    Span4Mux_h I__7826 (
            .O(N__34864),
            .I(N__34845));
    InMux I__7825 (
            .O(N__34863),
            .I(N__34840));
    InMux I__7824 (
            .O(N__34862),
            .I(N__34840));
    Span4Mux_h I__7823 (
            .O(N__34859),
            .I(N__34837));
    Span4Mux_h I__7822 (
            .O(N__34856),
            .I(N__34834));
    InMux I__7821 (
            .O(N__34855),
            .I(N__34827));
    InMux I__7820 (
            .O(N__34854),
            .I(N__34827));
    InMux I__7819 (
            .O(N__34851),
            .I(N__34827));
    LocalMux I__7818 (
            .O(N__34848),
            .I(aluOperand2_fast_2));
    Odrv4 I__7817 (
            .O(N__34845),
            .I(aluOperand2_fast_2));
    LocalMux I__7816 (
            .O(N__34840),
            .I(aluOperand2_fast_2));
    Odrv4 I__7815 (
            .O(N__34837),
            .I(aluOperand2_fast_2));
    Odrv4 I__7814 (
            .O(N__34834),
            .I(aluOperand2_fast_2));
    LocalMux I__7813 (
            .O(N__34827),
            .I(aluOperand2_fast_2));
    InMux I__7812 (
            .O(N__34814),
            .I(N__34811));
    LocalMux I__7811 (
            .O(N__34811),
            .I(N__34808));
    Span4Mux_h I__7810 (
            .O(N__34808),
            .I(N__34805));
    Span4Mux_h I__7809 (
            .O(N__34805),
            .I(N__34802));
    Odrv4 I__7808 (
            .O(N__34802),
            .I(\ALU.g0_7_m4_1 ));
    InMux I__7807 (
            .O(N__34799),
            .I(N__34791));
    InMux I__7806 (
            .O(N__34798),
            .I(N__34788));
    InMux I__7805 (
            .O(N__34797),
            .I(N__34784));
    InMux I__7804 (
            .O(N__34796),
            .I(N__34777));
    InMux I__7803 (
            .O(N__34795),
            .I(N__34777));
    InMux I__7802 (
            .O(N__34794),
            .I(N__34777));
    LocalMux I__7801 (
            .O(N__34791),
            .I(N__34774));
    LocalMux I__7800 (
            .O(N__34788),
            .I(N__34771));
    CascadeMux I__7799 (
            .O(N__34787),
            .I(N__34766));
    LocalMux I__7798 (
            .O(N__34784),
            .I(N__34759));
    LocalMux I__7797 (
            .O(N__34777),
            .I(N__34759));
    Span4Mux_v I__7796 (
            .O(N__34774),
            .I(N__34756));
    Span4Mux_v I__7795 (
            .O(N__34771),
            .I(N__34753));
    InMux I__7794 (
            .O(N__34770),
            .I(N__34748));
    InMux I__7793 (
            .O(N__34769),
            .I(N__34748));
    InMux I__7792 (
            .O(N__34766),
            .I(N__34741));
    InMux I__7791 (
            .O(N__34765),
            .I(N__34741));
    InMux I__7790 (
            .O(N__34764),
            .I(N__34741));
    Span4Mux_v I__7789 (
            .O(N__34759),
            .I(N__34738));
    Sp12to4 I__7788 (
            .O(N__34756),
            .I(N__34735));
    Sp12to4 I__7787 (
            .O(N__34753),
            .I(N__34732));
    LocalMux I__7786 (
            .O(N__34748),
            .I(N_287_0));
    LocalMux I__7785 (
            .O(N__34741),
            .I(N_287_0));
    Odrv4 I__7784 (
            .O(N__34738),
            .I(N_287_0));
    Odrv12 I__7783 (
            .O(N__34735),
            .I(N_287_0));
    Odrv12 I__7782 (
            .O(N__34732),
            .I(N_287_0));
    CascadeMux I__7781 (
            .O(N__34721),
            .I(N__34717));
    CascadeMux I__7780 (
            .O(N__34720),
            .I(N__34711));
    InMux I__7779 (
            .O(N__34717),
            .I(N__34705));
    InMux I__7778 (
            .O(N__34716),
            .I(N__34698));
    InMux I__7777 (
            .O(N__34715),
            .I(N__34698));
    InMux I__7776 (
            .O(N__34714),
            .I(N__34698));
    InMux I__7775 (
            .O(N__34711),
            .I(N__34695));
    CEMux I__7774 (
            .O(N__34710),
            .I(N__34692));
    CascadeMux I__7773 (
            .O(N__34709),
            .I(N__34688));
    CascadeMux I__7772 (
            .O(N__34708),
            .I(N__34682));
    LocalMux I__7771 (
            .O(N__34705),
            .I(N__34678));
    LocalMux I__7770 (
            .O(N__34698),
            .I(N__34675));
    LocalMux I__7769 (
            .O(N__34695),
            .I(N__34672));
    LocalMux I__7768 (
            .O(N__34692),
            .I(N__34669));
    CEMux I__7767 (
            .O(N__34691),
            .I(N__34665));
    InMux I__7766 (
            .O(N__34688),
            .I(N__34662));
    InMux I__7765 (
            .O(N__34687),
            .I(N__34657));
    InMux I__7764 (
            .O(N__34686),
            .I(N__34657));
    InMux I__7763 (
            .O(N__34685),
            .I(N__34652));
    InMux I__7762 (
            .O(N__34682),
            .I(N__34652));
    InMux I__7761 (
            .O(N__34681),
            .I(N__34649));
    Span4Mux_h I__7760 (
            .O(N__34678),
            .I(N__34646));
    Span4Mux_v I__7759 (
            .O(N__34675),
            .I(N__34643));
    Span4Mux_h I__7758 (
            .O(N__34672),
            .I(N__34640));
    Span4Mux_s3_h I__7757 (
            .O(N__34669),
            .I(N__34637));
    InMux I__7756 (
            .O(N__34668),
            .I(N__34634));
    LocalMux I__7755 (
            .O(N__34665),
            .I(N__34631));
    LocalMux I__7754 (
            .O(N__34662),
            .I(N__34624));
    LocalMux I__7753 (
            .O(N__34657),
            .I(N__34624));
    LocalMux I__7752 (
            .O(N__34652),
            .I(N__34624));
    LocalMux I__7751 (
            .O(N__34649),
            .I(N__34621));
    Span4Mux_h I__7750 (
            .O(N__34646),
            .I(N__34618));
    Span4Mux_h I__7749 (
            .O(N__34643),
            .I(N__34613));
    Span4Mux_h I__7748 (
            .O(N__34640),
            .I(N__34610));
    Span4Mux_h I__7747 (
            .O(N__34637),
            .I(N__34605));
    LocalMux I__7746 (
            .O(N__34634),
            .I(N__34605));
    Span4Mux_v I__7745 (
            .O(N__34631),
            .I(N__34601));
    Span12Mux_h I__7744 (
            .O(N__34624),
            .I(N__34594));
    Sp12to4 I__7743 (
            .O(N__34621),
            .I(N__34594));
    Sp12to4 I__7742 (
            .O(N__34618),
            .I(N__34594));
    InMux I__7741 (
            .O(N__34617),
            .I(N__34589));
    InMux I__7740 (
            .O(N__34616),
            .I(N__34589));
    Span4Mux_h I__7739 (
            .O(N__34613),
            .I(N__34582));
    Span4Mux_v I__7738 (
            .O(N__34610),
            .I(N__34582));
    Span4Mux_s3_h I__7737 (
            .O(N__34605),
            .I(N__34582));
    InMux I__7736 (
            .O(N__34604),
            .I(N__34579));
    Odrv4 I__7735 (
            .O(N__34601),
            .I(G_566));
    Odrv12 I__7734 (
            .O(N__34594),
            .I(G_566));
    LocalMux I__7733 (
            .O(N__34589),
            .I(G_566));
    Odrv4 I__7732 (
            .O(N__34582),
            .I(G_566));
    LocalMux I__7731 (
            .O(N__34579),
            .I(G_566));
    CascadeMux I__7730 (
            .O(N__34568),
            .I(N__34563));
    InMux I__7729 (
            .O(N__34567),
            .I(N__34558));
    InMux I__7728 (
            .O(N__34566),
            .I(N__34558));
    InMux I__7727 (
            .O(N__34563),
            .I(N__34555));
    LocalMux I__7726 (
            .O(N__34558),
            .I(N__34552));
    LocalMux I__7725 (
            .O(N__34555),
            .I(N__34549));
    Span4Mux_v I__7724 (
            .O(N__34552),
            .I(N__34546));
    Span4Mux_v I__7723 (
            .O(N__34549),
            .I(N__34542));
    Sp12to4 I__7722 (
            .O(N__34546),
            .I(N__34539));
    CascadeMux I__7721 (
            .O(N__34545),
            .I(N__34536));
    Span4Mux_v I__7720 (
            .O(N__34542),
            .I(N__34533));
    Span12Mux_h I__7719 (
            .O(N__34539),
            .I(N__34530));
    InMux I__7718 (
            .O(N__34536),
            .I(N__34527));
    Sp12to4 I__7717 (
            .O(N__34533),
            .I(N__34524));
    Span12Mux_v I__7716 (
            .O(N__34530),
            .I(N__34521));
    LocalMux I__7715 (
            .O(N__34527),
            .I(testWordZ0Z_11));
    Odrv12 I__7714 (
            .O(N__34524),
            .I(testWordZ0Z_11));
    Odrv12 I__7713 (
            .O(N__34521),
            .I(testWordZ0Z_11));
    CascadeMux I__7712 (
            .O(N__34514),
            .I(N__34509));
    InMux I__7711 (
            .O(N__34513),
            .I(N__34505));
    InMux I__7710 (
            .O(N__34512),
            .I(N__34502));
    InMux I__7709 (
            .O(N__34509),
            .I(N__34497));
    InMux I__7708 (
            .O(N__34508),
            .I(N__34497));
    LocalMux I__7707 (
            .O(N__34505),
            .I(N__34489));
    LocalMux I__7706 (
            .O(N__34502),
            .I(N__34489));
    LocalMux I__7705 (
            .O(N__34497),
            .I(N__34485));
    InMux I__7704 (
            .O(N__34496),
            .I(N__34482));
    InMux I__7703 (
            .O(N__34495),
            .I(N__34479));
    InMux I__7702 (
            .O(N__34494),
            .I(N__34476));
    Span4Mux_v I__7701 (
            .O(N__34489),
            .I(N__34470));
    InMux I__7700 (
            .O(N__34488),
            .I(N__34465));
    Span4Mux_v I__7699 (
            .O(N__34485),
            .I(N__34462));
    LocalMux I__7698 (
            .O(N__34482),
            .I(N__34459));
    LocalMux I__7697 (
            .O(N__34479),
            .I(N__34454));
    LocalMux I__7696 (
            .O(N__34476),
            .I(N__34454));
    InMux I__7695 (
            .O(N__34475),
            .I(N__34447));
    InMux I__7694 (
            .O(N__34474),
            .I(N__34447));
    InMux I__7693 (
            .O(N__34473),
            .I(N__34447));
    Span4Mux_h I__7692 (
            .O(N__34470),
            .I(N__34444));
    InMux I__7691 (
            .O(N__34469),
            .I(N__34439));
    InMux I__7690 (
            .O(N__34468),
            .I(N__34439));
    LocalMux I__7689 (
            .O(N__34465),
            .I(N__34434));
    Span4Mux_h I__7688 (
            .O(N__34462),
            .I(N__34434));
    Span4Mux_h I__7687 (
            .O(N__34459),
            .I(N__34431));
    Span4Mux_h I__7686 (
            .O(N__34454),
            .I(N__34424));
    LocalMux I__7685 (
            .O(N__34447),
            .I(N__34424));
    Span4Mux_h I__7684 (
            .O(N__34444),
            .I(N__34424));
    LocalMux I__7683 (
            .O(N__34439),
            .I(aluOperand2_1));
    Odrv4 I__7682 (
            .O(N__34434),
            .I(aluOperand2_1));
    Odrv4 I__7681 (
            .O(N__34431),
            .I(aluOperand2_1));
    Odrv4 I__7680 (
            .O(N__34424),
            .I(aluOperand2_1));
    CascadeMux I__7679 (
            .O(N__34415),
            .I(N__34412));
    InMux I__7678 (
            .O(N__34412),
            .I(N__34408));
    InMux I__7677 (
            .O(N__34411),
            .I(N__34405));
    LocalMux I__7676 (
            .O(N__34408),
            .I(N__34399));
    LocalMux I__7675 (
            .O(N__34405),
            .I(N__34396));
    InMux I__7674 (
            .O(N__34404),
            .I(N__34391));
    InMux I__7673 (
            .O(N__34403),
            .I(N__34388));
    InMux I__7672 (
            .O(N__34402),
            .I(N__34385));
    Span4Mux_v I__7671 (
            .O(N__34399),
            .I(N__34381));
    Span4Mux_h I__7670 (
            .O(N__34396),
            .I(N__34378));
    InMux I__7669 (
            .O(N__34395),
            .I(N__34375));
    InMux I__7668 (
            .O(N__34394),
            .I(N__34372));
    LocalMux I__7667 (
            .O(N__34391),
            .I(N__34369));
    LocalMux I__7666 (
            .O(N__34388),
            .I(N__34364));
    LocalMux I__7665 (
            .O(N__34385),
            .I(N__34364));
    InMux I__7664 (
            .O(N__34384),
            .I(N__34361));
    Odrv4 I__7663 (
            .O(N__34381),
            .I(\ALU.mult_10 ));
    Odrv4 I__7662 (
            .O(N__34378),
            .I(\ALU.mult_10 ));
    LocalMux I__7661 (
            .O(N__34375),
            .I(\ALU.mult_10 ));
    LocalMux I__7660 (
            .O(N__34372),
            .I(\ALU.mult_10 ));
    Odrv4 I__7659 (
            .O(N__34369),
            .I(\ALU.mult_10 ));
    Odrv12 I__7658 (
            .O(N__34364),
            .I(\ALU.mult_10 ));
    LocalMux I__7657 (
            .O(N__34361),
            .I(\ALU.mult_10 ));
    InMux I__7656 (
            .O(N__34346),
            .I(N__34339));
    InMux I__7655 (
            .O(N__34345),
            .I(N__34336));
    InMux I__7654 (
            .O(N__34344),
            .I(N__34333));
    InMux I__7653 (
            .O(N__34343),
            .I(N__34330));
    InMux I__7652 (
            .O(N__34342),
            .I(N__34327));
    LocalMux I__7651 (
            .O(N__34339),
            .I(N__34317));
    LocalMux I__7650 (
            .O(N__34336),
            .I(N__34317));
    LocalMux I__7649 (
            .O(N__34333),
            .I(N__34317));
    LocalMux I__7648 (
            .O(N__34330),
            .I(N__34317));
    LocalMux I__7647 (
            .O(N__34327),
            .I(N__34314));
    InMux I__7646 (
            .O(N__34326),
            .I(N__34311));
    Span4Mux_v I__7645 (
            .O(N__34317),
            .I(N__34307));
    Span4Mux_v I__7644 (
            .O(N__34314),
            .I(N__34304));
    LocalMux I__7643 (
            .O(N__34311),
            .I(N__34301));
    InMux I__7642 (
            .O(N__34310),
            .I(N__34298));
    Span4Mux_h I__7641 (
            .O(N__34307),
            .I(N__34295));
    Sp12to4 I__7640 (
            .O(N__34304),
            .I(N__34288));
    Span12Mux_v I__7639 (
            .O(N__34301),
            .I(N__34288));
    LocalMux I__7638 (
            .O(N__34298),
            .I(N__34288));
    Odrv4 I__7637 (
            .O(N__34295),
            .I(aluOperation_RNINNN4N3_0));
    Odrv12 I__7636 (
            .O(N__34288),
            .I(aluOperation_RNINNN4N3_0));
    InMux I__7635 (
            .O(N__34283),
            .I(N__34279));
    InMux I__7634 (
            .O(N__34282),
            .I(N__34276));
    LocalMux I__7633 (
            .O(N__34279),
            .I(N__34273));
    LocalMux I__7632 (
            .O(N__34276),
            .I(N__34270));
    Span4Mux_v I__7631 (
            .O(N__34273),
            .I(N__34264));
    Span4Mux_h I__7630 (
            .O(N__34270),
            .I(N__34264));
    CascadeMux I__7629 (
            .O(N__34269),
            .I(N__34261));
    Span4Mux_h I__7628 (
            .O(N__34264),
            .I(N__34258));
    InMux I__7627 (
            .O(N__34261),
            .I(N__34255));
    Odrv4 I__7626 (
            .O(N__34258),
            .I(\ALU.gZ0Z_10 ));
    LocalMux I__7625 (
            .O(N__34255),
            .I(\ALU.gZ0Z_10 ));
    InMux I__7624 (
            .O(N__34250),
            .I(N__34242));
    InMux I__7623 (
            .O(N__34249),
            .I(N__34239));
    InMux I__7622 (
            .O(N__34248),
            .I(N__34236));
    InMux I__7621 (
            .O(N__34247),
            .I(N__34233));
    InMux I__7620 (
            .O(N__34246),
            .I(N__34230));
    InMux I__7619 (
            .O(N__34245),
            .I(N__34227));
    LocalMux I__7618 (
            .O(N__34242),
            .I(N__34224));
    LocalMux I__7617 (
            .O(N__34239),
            .I(N__34215));
    LocalMux I__7616 (
            .O(N__34236),
            .I(N__34215));
    LocalMux I__7615 (
            .O(N__34233),
            .I(N__34215));
    LocalMux I__7614 (
            .O(N__34230),
            .I(N__34215));
    LocalMux I__7613 (
            .O(N__34227),
            .I(N__34211));
    Span4Mux_h I__7612 (
            .O(N__34224),
            .I(N__34208));
    Span4Mux_v I__7611 (
            .O(N__34215),
            .I(N__34205));
    InMux I__7610 (
            .O(N__34214),
            .I(N__34202));
    Span4Mux_h I__7609 (
            .O(N__34211),
            .I(N__34199));
    Span4Mux_h I__7608 (
            .O(N__34208),
            .I(N__34196));
    Sp12to4 I__7607 (
            .O(N__34205),
            .I(N__34193));
    LocalMux I__7606 (
            .O(N__34202),
            .I(N__34190));
    Odrv4 I__7605 (
            .O(N__34199),
            .I(aluOperation_RNI5QD2L3_0));
    Odrv4 I__7604 (
            .O(N__34196),
            .I(aluOperation_RNI5QD2L3_0));
    Odrv12 I__7603 (
            .O(N__34193),
            .I(aluOperation_RNI5QD2L3_0));
    Odrv12 I__7602 (
            .O(N__34190),
            .I(aluOperation_RNI5QD2L3_0));
    InMux I__7601 (
            .O(N__34181),
            .I(N__34176));
    InMux I__7600 (
            .O(N__34180),
            .I(N__34171));
    InMux I__7599 (
            .O(N__34179),
            .I(N__34168));
    LocalMux I__7598 (
            .O(N__34176),
            .I(N__34164));
    InMux I__7597 (
            .O(N__34175),
            .I(N__34161));
    InMux I__7596 (
            .O(N__34174),
            .I(N__34157));
    LocalMux I__7595 (
            .O(N__34171),
            .I(N__34154));
    LocalMux I__7594 (
            .O(N__34168),
            .I(N__34151));
    InMux I__7593 (
            .O(N__34167),
            .I(N__34148));
    Span4Mux_h I__7592 (
            .O(N__34164),
            .I(N__34144));
    LocalMux I__7591 (
            .O(N__34161),
            .I(N__34141));
    InMux I__7590 (
            .O(N__34160),
            .I(N__34138));
    LocalMux I__7589 (
            .O(N__34157),
            .I(N__34135));
    Span4Mux_v I__7588 (
            .O(N__34154),
            .I(N__34128));
    Span4Mux_h I__7587 (
            .O(N__34151),
            .I(N__34128));
    LocalMux I__7586 (
            .O(N__34148),
            .I(N__34128));
    InMux I__7585 (
            .O(N__34147),
            .I(N__34125));
    Odrv4 I__7584 (
            .O(N__34144),
            .I(\ALU.mult_11 ));
    Odrv4 I__7583 (
            .O(N__34141),
            .I(\ALU.mult_11 ));
    LocalMux I__7582 (
            .O(N__34138),
            .I(\ALU.mult_11 ));
    Odrv4 I__7581 (
            .O(N__34135),
            .I(\ALU.mult_11 ));
    Odrv4 I__7580 (
            .O(N__34128),
            .I(\ALU.mult_11 ));
    LocalMux I__7579 (
            .O(N__34125),
            .I(\ALU.mult_11 ));
    InMux I__7578 (
            .O(N__34112),
            .I(N__34109));
    LocalMux I__7577 (
            .O(N__34109),
            .I(N__34106));
    Span4Mux_v I__7576 (
            .O(N__34106),
            .I(N__34102));
    InMux I__7575 (
            .O(N__34105),
            .I(N__34099));
    Span4Mux_h I__7574 (
            .O(N__34102),
            .I(N__34094));
    LocalMux I__7573 (
            .O(N__34099),
            .I(N__34094));
    Odrv4 I__7572 (
            .O(N__34094),
            .I(\ALU.gZ0Z_11 ));
    InMux I__7571 (
            .O(N__34091),
            .I(N__34083));
    InMux I__7570 (
            .O(N__34090),
            .I(N__34080));
    InMux I__7569 (
            .O(N__34089),
            .I(N__34077));
    CascadeMux I__7568 (
            .O(N__34088),
            .I(N__34073));
    InMux I__7567 (
            .O(N__34087),
            .I(N__34070));
    InMux I__7566 (
            .O(N__34086),
            .I(N__34067));
    LocalMux I__7565 (
            .O(N__34083),
            .I(N__34064));
    LocalMux I__7564 (
            .O(N__34080),
            .I(N__34059));
    LocalMux I__7563 (
            .O(N__34077),
            .I(N__34059));
    InMux I__7562 (
            .O(N__34076),
            .I(N__34056));
    InMux I__7561 (
            .O(N__34073),
            .I(N__34053));
    LocalMux I__7560 (
            .O(N__34070),
            .I(N__34048));
    LocalMux I__7559 (
            .O(N__34067),
            .I(N__34048));
    Span4Mux_v I__7558 (
            .O(N__34064),
            .I(N__34045));
    Span4Mux_v I__7557 (
            .O(N__34059),
            .I(N__34042));
    LocalMux I__7556 (
            .O(N__34056),
            .I(aluOperation_RNIGPL5M3_0));
    LocalMux I__7555 (
            .O(N__34053),
            .I(aluOperation_RNIGPL5M3_0));
    Odrv4 I__7554 (
            .O(N__34048),
            .I(aluOperation_RNIGPL5M3_0));
    Odrv4 I__7553 (
            .O(N__34045),
            .I(aluOperation_RNIGPL5M3_0));
    Odrv4 I__7552 (
            .O(N__34042),
            .I(aluOperation_RNIGPL5M3_0));
    InMux I__7551 (
            .O(N__34031),
            .I(N__34027));
    InMux I__7550 (
            .O(N__34030),
            .I(N__34022));
    LocalMux I__7549 (
            .O(N__34027),
            .I(N__34017));
    InMux I__7548 (
            .O(N__34026),
            .I(N__34014));
    InMux I__7547 (
            .O(N__34025),
            .I(N__34011));
    LocalMux I__7546 (
            .O(N__34022),
            .I(N__34007));
    InMux I__7545 (
            .O(N__34021),
            .I(N__34004));
    InMux I__7544 (
            .O(N__34020),
            .I(N__34001));
    Span4Mux_h I__7543 (
            .O(N__34017),
            .I(N__33997));
    LocalMux I__7542 (
            .O(N__34014),
            .I(N__33994));
    LocalMux I__7541 (
            .O(N__34011),
            .I(N__33991));
    InMux I__7540 (
            .O(N__34010),
            .I(N__33988));
    Span4Mux_v I__7539 (
            .O(N__34007),
            .I(N__33983));
    LocalMux I__7538 (
            .O(N__34004),
            .I(N__33983));
    LocalMux I__7537 (
            .O(N__34001),
            .I(N__33980));
    InMux I__7536 (
            .O(N__34000),
            .I(N__33977));
    Odrv4 I__7535 (
            .O(N__33997),
            .I(\ALU.mult_12 ));
    Odrv4 I__7534 (
            .O(N__33994),
            .I(\ALU.mult_12 ));
    Odrv4 I__7533 (
            .O(N__33991),
            .I(\ALU.mult_12 ));
    LocalMux I__7532 (
            .O(N__33988),
            .I(\ALU.mult_12 ));
    Odrv4 I__7531 (
            .O(N__33983),
            .I(\ALU.mult_12 ));
    Odrv4 I__7530 (
            .O(N__33980),
            .I(\ALU.mult_12 ));
    LocalMux I__7529 (
            .O(N__33977),
            .I(\ALU.mult_12 ));
    InMux I__7528 (
            .O(N__33962),
            .I(N__33959));
    LocalMux I__7527 (
            .O(N__33959),
            .I(N__33955));
    InMux I__7526 (
            .O(N__33958),
            .I(N__33952));
    Span4Mux_h I__7525 (
            .O(N__33955),
            .I(N__33947));
    LocalMux I__7524 (
            .O(N__33952),
            .I(N__33947));
    Span4Mux_h I__7523 (
            .O(N__33947),
            .I(N__33944));
    Odrv4 I__7522 (
            .O(N__33944),
            .I(\ALU.gZ0Z_12 ));
    CascadeMux I__7521 (
            .O(N__33941),
            .I(N__33936));
    InMux I__7520 (
            .O(N__33940),
            .I(N__33931));
    InMux I__7519 (
            .O(N__33939),
            .I(N__33928));
    InMux I__7518 (
            .O(N__33936),
            .I(N__33925));
    InMux I__7517 (
            .O(N__33935),
            .I(N__33922));
    InMux I__7516 (
            .O(N__33934),
            .I(N__33917));
    LocalMux I__7515 (
            .O(N__33931),
            .I(N__33914));
    LocalMux I__7514 (
            .O(N__33928),
            .I(N__33911));
    LocalMux I__7513 (
            .O(N__33925),
            .I(N__33906));
    LocalMux I__7512 (
            .O(N__33922),
            .I(N__33906));
    InMux I__7511 (
            .O(N__33921),
            .I(N__33903));
    InMux I__7510 (
            .O(N__33920),
            .I(N__33900));
    LocalMux I__7509 (
            .O(N__33917),
            .I(N__33895));
    Span4Mux_h I__7508 (
            .O(N__33914),
            .I(N__33895));
    Span4Mux_h I__7507 (
            .O(N__33911),
            .I(N__33890));
    Span4Mux_v I__7506 (
            .O(N__33906),
            .I(N__33890));
    LocalMux I__7505 (
            .O(N__33903),
            .I(aluOperation_RNI2J9SL3_0));
    LocalMux I__7504 (
            .O(N__33900),
            .I(aluOperation_RNI2J9SL3_0));
    Odrv4 I__7503 (
            .O(N__33895),
            .I(aluOperation_RNI2J9SL3_0));
    Odrv4 I__7502 (
            .O(N__33890),
            .I(aluOperation_RNI2J9SL3_0));
    InMux I__7501 (
            .O(N__33881),
            .I(N__33877));
    InMux I__7500 (
            .O(N__33880),
            .I(N__33874));
    LocalMux I__7499 (
            .O(N__33877),
            .I(N__33868));
    LocalMux I__7498 (
            .O(N__33874),
            .I(N__33865));
    InMux I__7497 (
            .O(N__33873),
            .I(N__33860));
    InMux I__7496 (
            .O(N__33872),
            .I(N__33857));
    InMux I__7495 (
            .O(N__33871),
            .I(N__33854));
    Span4Mux_h I__7494 (
            .O(N__33868),
            .I(N__33848));
    Span4Mux_h I__7493 (
            .O(N__33865),
            .I(N__33848));
    InMux I__7492 (
            .O(N__33864),
            .I(N__33845));
    InMux I__7491 (
            .O(N__33863),
            .I(N__33842));
    LocalMux I__7490 (
            .O(N__33860),
            .I(N__33839));
    LocalMux I__7489 (
            .O(N__33857),
            .I(N__33834));
    LocalMux I__7488 (
            .O(N__33854),
            .I(N__33834));
    InMux I__7487 (
            .O(N__33853),
            .I(N__33831));
    Odrv4 I__7486 (
            .O(N__33848),
            .I(\ALU.mult_13 ));
    LocalMux I__7485 (
            .O(N__33845),
            .I(\ALU.mult_13 ));
    LocalMux I__7484 (
            .O(N__33842),
            .I(\ALU.mult_13 ));
    Odrv4 I__7483 (
            .O(N__33839),
            .I(\ALU.mult_13 ));
    Odrv4 I__7482 (
            .O(N__33834),
            .I(\ALU.mult_13 ));
    LocalMux I__7481 (
            .O(N__33831),
            .I(\ALU.mult_13 ));
    InMux I__7480 (
            .O(N__33818),
            .I(N__33809));
    InMux I__7479 (
            .O(N__33817),
            .I(N__33806));
    InMux I__7478 (
            .O(N__33816),
            .I(N__33803));
    InMux I__7477 (
            .O(N__33815),
            .I(N__33800));
    InMux I__7476 (
            .O(N__33814),
            .I(N__33797));
    InMux I__7475 (
            .O(N__33813),
            .I(N__33794));
    InMux I__7474 (
            .O(N__33812),
            .I(N__33791));
    LocalMux I__7473 (
            .O(N__33809),
            .I(N__33788));
    LocalMux I__7472 (
            .O(N__33806),
            .I(N__33785));
    LocalMux I__7471 (
            .O(N__33803),
            .I(N__33782));
    LocalMux I__7470 (
            .O(N__33800),
            .I(N__33769));
    LocalMux I__7469 (
            .O(N__33797),
            .I(N__33769));
    LocalMux I__7468 (
            .O(N__33794),
            .I(N__33769));
    LocalMux I__7467 (
            .O(N__33791),
            .I(N__33769));
    Span4Mux_h I__7466 (
            .O(N__33788),
            .I(N__33769));
    Span4Mux_v I__7465 (
            .O(N__33785),
            .I(N__33769));
    Span4Mux_h I__7464 (
            .O(N__33782),
            .I(N__33766));
    Span4Mux_v I__7463 (
            .O(N__33769),
            .I(N__33763));
    Odrv4 I__7462 (
            .O(N__33766),
            .I(aluOperation_RNIR872K3_0));
    Odrv4 I__7461 (
            .O(N__33763),
            .I(aluOperation_RNIR872K3_0));
    InMux I__7460 (
            .O(N__33758),
            .I(N__33753));
    InMux I__7459 (
            .O(N__33757),
            .I(N__33750));
    InMux I__7458 (
            .O(N__33756),
            .I(N__33744));
    LocalMux I__7457 (
            .O(N__33753),
            .I(N__33741));
    LocalMux I__7456 (
            .O(N__33750),
            .I(N__33737));
    InMux I__7455 (
            .O(N__33749),
            .I(N__33734));
    InMux I__7454 (
            .O(N__33748),
            .I(N__33731));
    InMux I__7453 (
            .O(N__33747),
            .I(N__33728));
    LocalMux I__7452 (
            .O(N__33744),
            .I(N__33724));
    Span4Mux_h I__7451 (
            .O(N__33741),
            .I(N__33721));
    InMux I__7450 (
            .O(N__33740),
            .I(N__33718));
    Span4Mux_h I__7449 (
            .O(N__33737),
            .I(N__33713));
    LocalMux I__7448 (
            .O(N__33734),
            .I(N__33713));
    LocalMux I__7447 (
            .O(N__33731),
            .I(N__33708));
    LocalMux I__7446 (
            .O(N__33728),
            .I(N__33708));
    InMux I__7445 (
            .O(N__33727),
            .I(N__33705));
    Odrv4 I__7444 (
            .O(N__33724),
            .I(\ALU.mult_14 ));
    Odrv4 I__7443 (
            .O(N__33721),
            .I(\ALU.mult_14 ));
    LocalMux I__7442 (
            .O(N__33718),
            .I(\ALU.mult_14 ));
    Odrv4 I__7441 (
            .O(N__33713),
            .I(\ALU.mult_14 ));
    Odrv4 I__7440 (
            .O(N__33708),
            .I(\ALU.mult_14 ));
    LocalMux I__7439 (
            .O(N__33705),
            .I(\ALU.mult_14 ));
    InMux I__7438 (
            .O(N__33692),
            .I(N__33689));
    LocalMux I__7437 (
            .O(N__33689),
            .I(N__33686));
    Span4Mux_h I__7436 (
            .O(N__33686),
            .I(N__33682));
    InMux I__7435 (
            .O(N__33685),
            .I(N__33679));
    Span4Mux_v I__7434 (
            .O(N__33682),
            .I(N__33676));
    LocalMux I__7433 (
            .O(N__33679),
            .I(N__33673));
    Span4Mux_h I__7432 (
            .O(N__33676),
            .I(N__33670));
    Span12Mux_s11_h I__7431 (
            .O(N__33673),
            .I(N__33667));
    Odrv4 I__7430 (
            .O(N__33670),
            .I(\ALU.gZ0Z_14 ));
    Odrv12 I__7429 (
            .O(N__33667),
            .I(\ALU.gZ0Z_14 ));
    InMux I__7428 (
            .O(N__33662),
            .I(N__33656));
    InMux I__7427 (
            .O(N__33661),
            .I(N__33650));
    InMux I__7426 (
            .O(N__33660),
            .I(N__33647));
    InMux I__7425 (
            .O(N__33659),
            .I(N__33644));
    LocalMux I__7424 (
            .O(N__33656),
            .I(N__33641));
    InMux I__7423 (
            .O(N__33655),
            .I(N__33638));
    InMux I__7422 (
            .O(N__33654),
            .I(N__33635));
    InMux I__7421 (
            .O(N__33653),
            .I(N__33632));
    LocalMux I__7420 (
            .O(N__33650),
            .I(N__33623));
    LocalMux I__7419 (
            .O(N__33647),
            .I(N__33623));
    LocalMux I__7418 (
            .O(N__33644),
            .I(N__33623));
    Span4Mux_h I__7417 (
            .O(N__33641),
            .I(N__33623));
    LocalMux I__7416 (
            .O(N__33638),
            .I(N__33620));
    LocalMux I__7415 (
            .O(N__33635),
            .I(N__33615));
    LocalMux I__7414 (
            .O(N__33632),
            .I(N__33615));
    Span4Mux_v I__7413 (
            .O(N__33623),
            .I(N__33612));
    Odrv4 I__7412 (
            .O(N__33620),
            .I(\ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93 ));
    Odrv4 I__7411 (
            .O(N__33615),
            .I(\ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93 ));
    Odrv4 I__7410 (
            .O(N__33612),
            .I(\ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93 ));
    InMux I__7409 (
            .O(N__33605),
            .I(N__33598));
    InMux I__7408 (
            .O(N__33604),
            .I(N__33595));
    InMux I__7407 (
            .O(N__33603),
            .I(N__33592));
    InMux I__7406 (
            .O(N__33602),
            .I(N__33586));
    InMux I__7405 (
            .O(N__33601),
            .I(N__33583));
    LocalMux I__7404 (
            .O(N__33598),
            .I(N__33580));
    LocalMux I__7403 (
            .O(N__33595),
            .I(N__33577));
    LocalMux I__7402 (
            .O(N__33592),
            .I(N__33574));
    InMux I__7401 (
            .O(N__33591),
            .I(N__33571));
    InMux I__7400 (
            .O(N__33590),
            .I(N__33568));
    InMux I__7399 (
            .O(N__33589),
            .I(N__33565));
    LocalMux I__7398 (
            .O(N__33586),
            .I(N__33562));
    LocalMux I__7397 (
            .O(N__33583),
            .I(N__33557));
    Span4Mux_h I__7396 (
            .O(N__33580),
            .I(N__33557));
    Span4Mux_h I__7395 (
            .O(N__33577),
            .I(N__33552));
    Span4Mux_h I__7394 (
            .O(N__33574),
            .I(N__33552));
    LocalMux I__7393 (
            .O(N__33571),
            .I(\ALU.mult_15 ));
    LocalMux I__7392 (
            .O(N__33568),
            .I(\ALU.mult_15 ));
    LocalMux I__7391 (
            .O(N__33565),
            .I(\ALU.mult_15 ));
    Odrv4 I__7390 (
            .O(N__33562),
            .I(\ALU.mult_15 ));
    Odrv4 I__7389 (
            .O(N__33557),
            .I(\ALU.mult_15 ));
    Odrv4 I__7388 (
            .O(N__33552),
            .I(\ALU.mult_15 ));
    InMux I__7387 (
            .O(N__33539),
            .I(N__33536));
    LocalMux I__7386 (
            .O(N__33536),
            .I(N__33532));
    InMux I__7385 (
            .O(N__33535),
            .I(N__33529));
    Span4Mux_v I__7384 (
            .O(N__33532),
            .I(N__33526));
    LocalMux I__7383 (
            .O(N__33529),
            .I(\ALU.gZ0Z_15 ));
    Odrv4 I__7382 (
            .O(N__33526),
            .I(\ALU.gZ0Z_15 ));
    CascadeMux I__7381 (
            .O(N__33521),
            .I(\ALU.a_15_m4_15_cascade_ ));
    InMux I__7380 (
            .O(N__33518),
            .I(N__33515));
    LocalMux I__7379 (
            .O(N__33515),
            .I(N__33512));
    Span4Mux_v I__7378 (
            .O(N__33512),
            .I(N__33509));
    Odrv4 I__7377 (
            .O(N__33509),
            .I(\ALU.a_15_m3_15 ));
    CascadeMux I__7376 (
            .O(N__33506),
            .I(\ALU.c_RNIR4QHM2Z0Z_15_cascade_ ));
    CascadeMux I__7375 (
            .O(N__33503),
            .I(\ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93_cascade_ ));
    InMux I__7374 (
            .O(N__33500),
            .I(N__33497));
    LocalMux I__7373 (
            .O(N__33497),
            .I(N__33494));
    Span4Mux_h I__7372 (
            .O(N__33494),
            .I(N__33491));
    Span4Mux_h I__7371 (
            .O(N__33491),
            .I(N__33488));
    Span4Mux_v I__7370 (
            .O(N__33488),
            .I(N__33484));
    InMux I__7369 (
            .O(N__33487),
            .I(N__33481));
    Odrv4 I__7368 (
            .O(N__33484),
            .I(\ALU.hZ0Z_15 ));
    LocalMux I__7367 (
            .O(N__33481),
            .I(\ALU.hZ0Z_15 ));
    InMux I__7366 (
            .O(N__33476),
            .I(N__33473));
    LocalMux I__7365 (
            .O(N__33473),
            .I(N__33469));
    InMux I__7364 (
            .O(N__33472),
            .I(N__33466));
    Span4Mux_h I__7363 (
            .O(N__33469),
            .I(N__33463));
    LocalMux I__7362 (
            .O(N__33466),
            .I(N__33460));
    Span4Mux_v I__7361 (
            .O(N__33463),
            .I(N__33457));
    Span4Mux_v I__7360 (
            .O(N__33460),
            .I(N__33454));
    Odrv4 I__7359 (
            .O(N__33457),
            .I(\ALU.dZ0Z_15 ));
    Odrv4 I__7358 (
            .O(N__33454),
            .I(\ALU.dZ0Z_15 ));
    InMux I__7357 (
            .O(N__33449),
            .I(N__33446));
    LocalMux I__7356 (
            .O(N__33446),
            .I(\ALU.d_RNISBLUZ0Z_15 ));
    InMux I__7355 (
            .O(N__33443),
            .I(N__33439));
    CEMux I__7354 (
            .O(N__33442),
            .I(N__33435));
    LocalMux I__7353 (
            .O(N__33439),
            .I(N__33431));
    InMux I__7352 (
            .O(N__33438),
            .I(N__33428));
    LocalMux I__7351 (
            .O(N__33435),
            .I(N__33425));
    InMux I__7350 (
            .O(N__33434),
            .I(N__33422));
    Sp12to4 I__7349 (
            .O(N__33431),
            .I(N__33419));
    LocalMux I__7348 (
            .O(N__33428),
            .I(N__33416));
    Span4Mux_h I__7347 (
            .O(N__33425),
            .I(N__33411));
    LocalMux I__7346 (
            .O(N__33422),
            .I(N__33411));
    Span12Mux_v I__7345 (
            .O(N__33419),
            .I(N__33408));
    Span12Mux_s4_v I__7344 (
            .O(N__33416),
            .I(N__33405));
    Span4Mux_s0_v I__7343 (
            .O(N__33411),
            .I(N__33402));
    Odrv12 I__7342 (
            .O(N__33408),
            .I(\CONTROL.aluOperation_cnvZ0Z_0 ));
    Odrv12 I__7341 (
            .O(N__33405),
            .I(\CONTROL.aluOperation_cnvZ0Z_0 ));
    Odrv4 I__7340 (
            .O(N__33402),
            .I(\CONTROL.aluOperation_cnvZ0Z_0 ));
    CascadeMux I__7339 (
            .O(N__33395),
            .I(N__33392));
    InMux I__7338 (
            .O(N__33392),
            .I(N__33389));
    LocalMux I__7337 (
            .O(N__33389),
            .I(N__33386));
    Span4Mux_h I__7336 (
            .O(N__33386),
            .I(N__33381));
    InMux I__7335 (
            .O(N__33385),
            .I(N__33376));
    InMux I__7334 (
            .O(N__33384),
            .I(N__33376));
    Span4Mux_h I__7333 (
            .O(N__33381),
            .I(N__33373));
    LocalMux I__7332 (
            .O(N__33376),
            .I(N__33370));
    Span4Mux_v I__7331 (
            .O(N__33373),
            .I(N__33367));
    Span4Mux_h I__7330 (
            .O(N__33370),
            .I(N__33362));
    Span4Mux_h I__7329 (
            .O(N__33367),
            .I(N__33362));
    Odrv4 I__7328 (
            .O(N__33362),
            .I(N_723));
    InMux I__7327 (
            .O(N__33359),
            .I(N__33351));
    InMux I__7326 (
            .O(N__33358),
            .I(N__33342));
    InMux I__7325 (
            .O(N__33357),
            .I(N__33342));
    InMux I__7324 (
            .O(N__33356),
            .I(N__33342));
    InMux I__7323 (
            .O(N__33355),
            .I(N__33342));
    InMux I__7322 (
            .O(N__33354),
            .I(N__33339));
    LocalMux I__7321 (
            .O(N__33351),
            .I(N__33336));
    LocalMux I__7320 (
            .O(N__33342),
            .I(N__33332));
    LocalMux I__7319 (
            .O(N__33339),
            .I(N__33325));
    Span4Mux_v I__7318 (
            .O(N__33336),
            .I(N__33325));
    CascadeMux I__7317 (
            .O(N__33335),
            .I(N__33322));
    Span4Mux_h I__7316 (
            .O(N__33332),
            .I(N__33319));
    InMux I__7315 (
            .O(N__33331),
            .I(N__33313));
    InMux I__7314 (
            .O(N__33330),
            .I(N__33310));
    Span4Mux_h I__7313 (
            .O(N__33325),
            .I(N__33307));
    InMux I__7312 (
            .O(N__33322),
            .I(N__33304));
    Span4Mux_v I__7311 (
            .O(N__33319),
            .I(N__33297));
    InMux I__7310 (
            .O(N__33318),
            .I(N__33287));
    InMux I__7309 (
            .O(N__33317),
            .I(N__33287));
    InMux I__7308 (
            .O(N__33316),
            .I(N__33287));
    LocalMux I__7307 (
            .O(N__33313),
            .I(N__33282));
    LocalMux I__7306 (
            .O(N__33310),
            .I(N__33282));
    Span4Mux_h I__7305 (
            .O(N__33307),
            .I(N__33279));
    LocalMux I__7304 (
            .O(N__33304),
            .I(N__33276));
    CascadeMux I__7303 (
            .O(N__33303),
            .I(N__33272));
    CascadeMux I__7302 (
            .O(N__33302),
            .I(N__33268));
    CascadeMux I__7301 (
            .O(N__33301),
            .I(N__33265));
    CascadeMux I__7300 (
            .O(N__33300),
            .I(N__33256));
    IoSpan4Mux I__7299 (
            .O(N__33297),
            .I(N__33253));
    InMux I__7298 (
            .O(N__33296),
            .I(N__33246));
    InMux I__7297 (
            .O(N__33295),
            .I(N__33246));
    InMux I__7296 (
            .O(N__33294),
            .I(N__33246));
    LocalMux I__7295 (
            .O(N__33287),
            .I(N__33240));
    Span4Mux_v I__7294 (
            .O(N__33282),
            .I(N__33240));
    Span4Mux_h I__7293 (
            .O(N__33279),
            .I(N__33237));
    Span4Mux_h I__7292 (
            .O(N__33276),
            .I(N__33234));
    InMux I__7291 (
            .O(N__33275),
            .I(N__33227));
    InMux I__7290 (
            .O(N__33272),
            .I(N__33227));
    InMux I__7289 (
            .O(N__33271),
            .I(N__33227));
    InMux I__7288 (
            .O(N__33268),
            .I(N__33220));
    InMux I__7287 (
            .O(N__33265),
            .I(N__33220));
    InMux I__7286 (
            .O(N__33264),
            .I(N__33220));
    InMux I__7285 (
            .O(N__33263),
            .I(N__33213));
    InMux I__7284 (
            .O(N__33262),
            .I(N__33213));
    InMux I__7283 (
            .O(N__33261),
            .I(N__33213));
    InMux I__7282 (
            .O(N__33260),
            .I(N__33210));
    InMux I__7281 (
            .O(N__33259),
            .I(N__33205));
    InMux I__7280 (
            .O(N__33256),
            .I(N__33205));
    Span4Mux_s0_v I__7279 (
            .O(N__33253),
            .I(N__33200));
    LocalMux I__7278 (
            .O(N__33246),
            .I(N__33200));
    InMux I__7277 (
            .O(N__33245),
            .I(N__33197));
    Span4Mux_h I__7276 (
            .O(N__33240),
            .I(N__33192));
    Span4Mux_v I__7275 (
            .O(N__33237),
            .I(N__33192));
    Odrv4 I__7274 (
            .O(N__33234),
            .I(testWordZ0Z_5));
    LocalMux I__7273 (
            .O(N__33227),
            .I(testWordZ0Z_5));
    LocalMux I__7272 (
            .O(N__33220),
            .I(testWordZ0Z_5));
    LocalMux I__7271 (
            .O(N__33213),
            .I(testWordZ0Z_5));
    LocalMux I__7270 (
            .O(N__33210),
            .I(testWordZ0Z_5));
    LocalMux I__7269 (
            .O(N__33205),
            .I(testWordZ0Z_5));
    Odrv4 I__7268 (
            .O(N__33200),
            .I(testWordZ0Z_5));
    LocalMux I__7267 (
            .O(N__33197),
            .I(testWordZ0Z_5));
    Odrv4 I__7266 (
            .O(N__33192),
            .I(testWordZ0Z_5));
    InMux I__7265 (
            .O(N__33173),
            .I(N__33170));
    LocalMux I__7264 (
            .O(N__33170),
            .I(N__33167));
    Span4Mux_h I__7263 (
            .O(N__33167),
            .I(N__33164));
    Span4Mux_h I__7262 (
            .O(N__33164),
            .I(N__33160));
    InMux I__7261 (
            .O(N__33163),
            .I(N__33157));
    Span4Mux_v I__7260 (
            .O(N__33160),
            .I(N__33154));
    LocalMux I__7259 (
            .O(N__33157),
            .I(aluOperation_5));
    Odrv4 I__7258 (
            .O(N__33154),
            .I(aluOperation_5));
    InMux I__7257 (
            .O(N__33149),
            .I(N__33145));
    CascadeMux I__7256 (
            .O(N__33148),
            .I(N__33142));
    LocalMux I__7255 (
            .O(N__33145),
            .I(N__33139));
    InMux I__7254 (
            .O(N__33142),
            .I(N__33136));
    Span4Mux_v I__7253 (
            .O(N__33139),
            .I(N__33133));
    LocalMux I__7252 (
            .O(N__33136),
            .I(N__33130));
    Span4Mux_v I__7251 (
            .O(N__33133),
            .I(N__33127));
    Span4Mux_h I__7250 (
            .O(N__33130),
            .I(N__33124));
    Span4Mux_h I__7249 (
            .O(N__33127),
            .I(N__33121));
    Span4Mux_v I__7248 (
            .O(N__33124),
            .I(N__33118));
    Odrv4 I__7247 (
            .O(N__33121),
            .I(\ALU.a2_b_0 ));
    Odrv4 I__7246 (
            .O(N__33118),
            .I(\ALU.a2_b_0 ));
    InMux I__7245 (
            .O(N__33113),
            .I(N__33110));
    LocalMux I__7244 (
            .O(N__33110),
            .I(N__33107));
    Odrv12 I__7243 (
            .O(N__33107),
            .I(\ALU.madd_axb_1_l_ofx ));
    CascadeMux I__7242 (
            .O(N__33104),
            .I(N__33100));
    CascadeMux I__7241 (
            .O(N__33103),
            .I(N__33097));
    InMux I__7240 (
            .O(N__33100),
            .I(N__33093));
    InMux I__7239 (
            .O(N__33097),
            .I(N__33090));
    CascadeMux I__7238 (
            .O(N__33096),
            .I(N__33086));
    LocalMux I__7237 (
            .O(N__33093),
            .I(N__33081));
    LocalMux I__7236 (
            .O(N__33090),
            .I(N__33078));
    InMux I__7235 (
            .O(N__33089),
            .I(N__33075));
    InMux I__7234 (
            .O(N__33086),
            .I(N__33072));
    InMux I__7233 (
            .O(N__33085),
            .I(N__33069));
    InMux I__7232 (
            .O(N__33084),
            .I(N__33066));
    Span4Mux_v I__7231 (
            .O(N__33081),
            .I(N__33055));
    Span4Mux_v I__7230 (
            .O(N__33078),
            .I(N__33055));
    LocalMux I__7229 (
            .O(N__33075),
            .I(N__33055));
    LocalMux I__7228 (
            .O(N__33072),
            .I(N__33052));
    LocalMux I__7227 (
            .O(N__33069),
            .I(N__33049));
    LocalMux I__7226 (
            .O(N__33066),
            .I(N__33045));
    InMux I__7225 (
            .O(N__33065),
            .I(N__33042));
    InMux I__7224 (
            .O(N__33064),
            .I(N__33037));
    InMux I__7223 (
            .O(N__33063),
            .I(N__33037));
    InMux I__7222 (
            .O(N__33062),
            .I(N__33034));
    Span4Mux_h I__7221 (
            .O(N__33055),
            .I(N__33031));
    Sp12to4 I__7220 (
            .O(N__33052),
            .I(N__33026));
    Sp12to4 I__7219 (
            .O(N__33049),
            .I(N__33026));
    InMux I__7218 (
            .O(N__33048),
            .I(N__33023));
    Span4Mux_v I__7217 (
            .O(N__33045),
            .I(N__33020));
    LocalMux I__7216 (
            .O(N__33042),
            .I(N__33013));
    LocalMux I__7215 (
            .O(N__33037),
            .I(N__33013));
    LocalMux I__7214 (
            .O(N__33034),
            .I(N__33013));
    Span4Mux_v I__7213 (
            .O(N__33031),
            .I(N__33010));
    Span12Mux_v I__7212 (
            .O(N__33026),
            .I(N__33007));
    LocalMux I__7211 (
            .O(N__33023),
            .I(aluOperand2_0_rep2));
    Odrv4 I__7210 (
            .O(N__33020),
            .I(aluOperand2_0_rep2));
    Odrv4 I__7209 (
            .O(N__33013),
            .I(aluOperand2_0_rep2));
    Odrv4 I__7208 (
            .O(N__33010),
            .I(aluOperand2_0_rep2));
    Odrv12 I__7207 (
            .O(N__33007),
            .I(aluOperand2_0_rep2));
    InMux I__7206 (
            .O(N__32996),
            .I(N__32987));
    InMux I__7205 (
            .O(N__32995),
            .I(N__32984));
    InMux I__7204 (
            .O(N__32994),
            .I(N__32980));
    InMux I__7203 (
            .O(N__32993),
            .I(N__32975));
    InMux I__7202 (
            .O(N__32992),
            .I(N__32975));
    InMux I__7201 (
            .O(N__32991),
            .I(N__32972));
    InMux I__7200 (
            .O(N__32990),
            .I(N__32967));
    LocalMux I__7199 (
            .O(N__32987),
            .I(N__32964));
    LocalMux I__7198 (
            .O(N__32984),
            .I(N__32960));
    InMux I__7197 (
            .O(N__32983),
            .I(N__32956));
    LocalMux I__7196 (
            .O(N__32980),
            .I(N__32953));
    LocalMux I__7195 (
            .O(N__32975),
            .I(N__32950));
    LocalMux I__7194 (
            .O(N__32972),
            .I(N__32947));
    InMux I__7193 (
            .O(N__32971),
            .I(N__32943));
    InMux I__7192 (
            .O(N__32970),
            .I(N__32940));
    LocalMux I__7191 (
            .O(N__32967),
            .I(N__32935));
    Span4Mux_s3_h I__7190 (
            .O(N__32964),
            .I(N__32935));
    InMux I__7189 (
            .O(N__32963),
            .I(N__32932));
    Span4Mux_h I__7188 (
            .O(N__32960),
            .I(N__32929));
    CascadeMux I__7187 (
            .O(N__32959),
            .I(N__32926));
    LocalMux I__7186 (
            .O(N__32956),
            .I(N__32921));
    Span4Mux_h I__7185 (
            .O(N__32953),
            .I(N__32921));
    Span4Mux_v I__7184 (
            .O(N__32950),
            .I(N__32918));
    Span4Mux_v I__7183 (
            .O(N__32947),
            .I(N__32915));
    InMux I__7182 (
            .O(N__32946),
            .I(N__32912));
    LocalMux I__7181 (
            .O(N__32943),
            .I(N__32909));
    LocalMux I__7180 (
            .O(N__32940),
            .I(N__32906));
    Span4Mux_h I__7179 (
            .O(N__32935),
            .I(N__32903));
    LocalMux I__7178 (
            .O(N__32932),
            .I(N__32899));
    Span4Mux_h I__7177 (
            .O(N__32929),
            .I(N__32896));
    InMux I__7176 (
            .O(N__32926),
            .I(N__32893));
    Span4Mux_h I__7175 (
            .O(N__32921),
            .I(N__32890));
    Span4Mux_h I__7174 (
            .O(N__32918),
            .I(N__32885));
    Span4Mux_h I__7173 (
            .O(N__32915),
            .I(N__32885));
    LocalMux I__7172 (
            .O(N__32912),
            .I(N__32876));
    Span4Mux_v I__7171 (
            .O(N__32909),
            .I(N__32876));
    Span4Mux_h I__7170 (
            .O(N__32906),
            .I(N__32876));
    Span4Mux_h I__7169 (
            .O(N__32903),
            .I(N__32876));
    InMux I__7168 (
            .O(N__32902),
            .I(N__32873));
    Span12Mux_v I__7167 (
            .O(N__32899),
            .I(N__32870));
    Span4Mux_v I__7166 (
            .O(N__32896),
            .I(N__32867));
    LocalMux I__7165 (
            .O(N__32893),
            .I(aluOperand2_0));
    Odrv4 I__7164 (
            .O(N__32890),
            .I(aluOperand2_0));
    Odrv4 I__7163 (
            .O(N__32885),
            .I(aluOperand2_0));
    Odrv4 I__7162 (
            .O(N__32876),
            .I(aluOperand2_0));
    LocalMux I__7161 (
            .O(N__32873),
            .I(aluOperand2_0));
    Odrv12 I__7160 (
            .O(N__32870),
            .I(aluOperand2_0));
    Odrv4 I__7159 (
            .O(N__32867),
            .I(aluOperand2_0));
    CascadeMux I__7158 (
            .O(N__32852),
            .I(\ALU.g_RNIVGLLZ0Z_9_cascade_ ));
    InMux I__7157 (
            .O(N__32849),
            .I(N__32846));
    LocalMux I__7156 (
            .O(N__32846),
            .I(N__32843));
    Odrv12 I__7155 (
            .O(N__32843),
            .I(\ALU.operand2_7_ns_1_9 ));
    InMux I__7154 (
            .O(N__32840),
            .I(N__32836));
    InMux I__7153 (
            .O(N__32839),
            .I(N__32833));
    LocalMux I__7152 (
            .O(N__32836),
            .I(N__32830));
    LocalMux I__7151 (
            .O(N__32833),
            .I(N__32827));
    Span4Mux_v I__7150 (
            .O(N__32830),
            .I(N__32824));
    Span4Mux_h I__7149 (
            .O(N__32827),
            .I(N__32821));
    Span4Mux_v I__7148 (
            .O(N__32824),
            .I(N__32818));
    Span4Mux_v I__7147 (
            .O(N__32821),
            .I(N__32814));
    Span4Mux_h I__7146 (
            .O(N__32818),
            .I(N__32811));
    InMux I__7145 (
            .O(N__32817),
            .I(N__32808));
    Span4Mux_h I__7144 (
            .O(N__32814),
            .I(N__32805));
    Odrv4 I__7143 (
            .O(N__32811),
            .I(\ALU.hZ0Z_9 ));
    LocalMux I__7142 (
            .O(N__32808),
            .I(\ALU.hZ0Z_9 ));
    Odrv4 I__7141 (
            .O(N__32805),
            .I(\ALU.hZ0Z_9 ));
    InMux I__7140 (
            .O(N__32798),
            .I(N__32793));
    InMux I__7139 (
            .O(N__32797),
            .I(N__32790));
    InMux I__7138 (
            .O(N__32796),
            .I(N__32787));
    LocalMux I__7137 (
            .O(N__32793),
            .I(N__32784));
    LocalMux I__7136 (
            .O(N__32790),
            .I(N__32781));
    LocalMux I__7135 (
            .O(N__32787),
            .I(N__32778));
    Span4Mux_v I__7134 (
            .O(N__32784),
            .I(N__32775));
    Span4Mux_h I__7133 (
            .O(N__32781),
            .I(N__32772));
    Span4Mux_v I__7132 (
            .O(N__32778),
            .I(N__32767));
    Span4Mux_v I__7131 (
            .O(N__32775),
            .I(N__32767));
    Span4Mux_h I__7130 (
            .O(N__32772),
            .I(N__32764));
    Odrv4 I__7129 (
            .O(N__32767),
            .I(\ALU.dZ0Z_9 ));
    Odrv4 I__7128 (
            .O(N__32764),
            .I(\ALU.dZ0Z_9 ));
    CascadeMux I__7127 (
            .O(N__32759),
            .I(N__32756));
    InMux I__7126 (
            .O(N__32756),
            .I(N__32753));
    LocalMux I__7125 (
            .O(N__32753),
            .I(N__32750));
    Span4Mux_h I__7124 (
            .O(N__32750),
            .I(N__32747));
    Span4Mux_h I__7123 (
            .O(N__32747),
            .I(N__32744));
    Odrv4 I__7122 (
            .O(N__32744),
            .I(\ALU.g0_0_0_m2_1 ));
    CascadeMux I__7121 (
            .O(N__32741),
            .I(\ALU.N_11_cascade_ ));
    InMux I__7120 (
            .O(N__32738),
            .I(N__32735));
    LocalMux I__7119 (
            .O(N__32735),
            .I(N__32732));
    Span4Mux_s3_h I__7118 (
            .O(N__32732),
            .I(N__32729));
    Span4Mux_h I__7117 (
            .O(N__32729),
            .I(N__32726));
    Span4Mux_h I__7116 (
            .O(N__32726),
            .I(N__32723));
    Odrv4 I__7115 (
            .O(N__32723),
            .I(\ALU.N_13 ));
    InMux I__7114 (
            .O(N__32720),
            .I(N__32717));
    LocalMux I__7113 (
            .O(N__32717),
            .I(N__32712));
    InMux I__7112 (
            .O(N__32716),
            .I(N__32707));
    InMux I__7111 (
            .O(N__32715),
            .I(N__32707));
    Span4Mux_h I__7110 (
            .O(N__32712),
            .I(N__32704));
    LocalMux I__7109 (
            .O(N__32707),
            .I(N__32701));
    Span4Mux_h I__7108 (
            .O(N__32704),
            .I(N__32696));
    Span4Mux_h I__7107 (
            .O(N__32701),
            .I(N__32696));
    Odrv4 I__7106 (
            .O(N__32696),
            .I(\ALU.cZ0Z_9 ));
    CascadeMux I__7105 (
            .O(N__32693),
            .I(N__32690));
    InMux I__7104 (
            .O(N__32690),
            .I(N__32687));
    LocalMux I__7103 (
            .O(N__32687),
            .I(\ALU.g0_0_0_m2_0_1 ));
    InMux I__7102 (
            .O(N__32684),
            .I(N__32681));
    LocalMux I__7101 (
            .O(N__32681),
            .I(N__32678));
    Odrv4 I__7100 (
            .O(N__32678),
            .I(\ALU.N_12 ));
    InMux I__7099 (
            .O(N__32675),
            .I(N__32671));
    InMux I__7098 (
            .O(N__32674),
            .I(N__32667));
    LocalMux I__7097 (
            .O(N__32671),
            .I(N__32662));
    CascadeMux I__7096 (
            .O(N__32670),
            .I(N__32658));
    LocalMux I__7095 (
            .O(N__32667),
            .I(N__32655));
    InMux I__7094 (
            .O(N__32666),
            .I(N__32652));
    CascadeMux I__7093 (
            .O(N__32665),
            .I(N__32649));
    Span4Mux_h I__7092 (
            .O(N__32662),
            .I(N__32646));
    InMux I__7091 (
            .O(N__32661),
            .I(N__32641));
    InMux I__7090 (
            .O(N__32658),
            .I(N__32641));
    Span12Mux_h I__7089 (
            .O(N__32655),
            .I(N__32638));
    LocalMux I__7088 (
            .O(N__32652),
            .I(N__32635));
    InMux I__7087 (
            .O(N__32649),
            .I(N__32632));
    Span4Mux_v I__7086 (
            .O(N__32646),
            .I(N__32627));
    LocalMux I__7085 (
            .O(N__32641),
            .I(N__32627));
    Odrv12 I__7084 (
            .O(N__32638),
            .I(\ALU.aluOut_15 ));
    Odrv12 I__7083 (
            .O(N__32635),
            .I(\ALU.aluOut_15 ));
    LocalMux I__7082 (
            .O(N__32632),
            .I(\ALU.aluOut_15 ));
    Odrv4 I__7081 (
            .O(N__32627),
            .I(\ALU.aluOut_15 ));
    CascadeMux I__7080 (
            .O(N__32618),
            .I(\ALU.a_15_m2_ns_1Z0Z_15_cascade_ ));
    InMux I__7079 (
            .O(N__32615),
            .I(N__32612));
    LocalMux I__7078 (
            .O(N__32612),
            .I(N__32609));
    Span4Mux_h I__7077 (
            .O(N__32609),
            .I(N__32605));
    InMux I__7076 (
            .O(N__32608),
            .I(N__32601));
    Span4Mux_h I__7075 (
            .O(N__32605),
            .I(N__32598));
    InMux I__7074 (
            .O(N__32604),
            .I(N__32595));
    LocalMux I__7073 (
            .O(N__32601),
            .I(N__32592));
    Odrv4 I__7072 (
            .O(N__32598),
            .I(\ALU.N_7_0 ));
    LocalMux I__7071 (
            .O(N__32595),
            .I(\ALU.N_7_0 ));
    Odrv12 I__7070 (
            .O(N__32592),
            .I(\ALU.N_7_0 ));
    CascadeMux I__7069 (
            .O(N__32585),
            .I(\ALU.a_15_m2_15_cascade_ ));
    InMux I__7068 (
            .O(N__32582),
            .I(N__32579));
    LocalMux I__7067 (
            .O(N__32579),
            .I(N__32576));
    Span4Mux_h I__7066 (
            .O(N__32576),
            .I(N__32573));
    Span4Mux_h I__7065 (
            .O(N__32573),
            .I(N__32570));
    Odrv4 I__7064 (
            .O(N__32570),
            .I(\ALU.lshift_15 ));
    InMux I__7063 (
            .O(N__32567),
            .I(N__32564));
    LocalMux I__7062 (
            .O(N__32564),
            .I(N__32561));
    Odrv12 I__7061 (
            .O(N__32561),
            .I(TXbufferZ0Z_7));
    InMux I__7060 (
            .O(N__32558),
            .I(N__32555));
    LocalMux I__7059 (
            .O(N__32555),
            .I(\FTDI.TXshiftZ0Z_7 ));
    InMux I__7058 (
            .O(N__32552),
            .I(N__32549));
    LocalMux I__7057 (
            .O(N__32549),
            .I(N__32546));
    Span4Mux_h I__7056 (
            .O(N__32546),
            .I(N__32543));
    Span4Mux_h I__7055 (
            .O(N__32543),
            .I(N__32540));
    Odrv4 I__7054 (
            .O(N__32540),
            .I(\ALU.un2_addsub_cry_10_c_RNIUS1OJZ0 ));
    CascadeMux I__7053 (
            .O(N__32537),
            .I(\ALU.a_15_m2_ns_1Z0Z_11_cascade_ ));
    CascadeMux I__7052 (
            .O(N__32534),
            .I(\ALU.a_15_m2_11_cascade_ ));
    InMux I__7051 (
            .O(N__32531),
            .I(N__32528));
    LocalMux I__7050 (
            .O(N__32528),
            .I(N__32525));
    Span4Mux_h I__7049 (
            .O(N__32525),
            .I(N__32522));
    Span4Mux_h I__7048 (
            .O(N__32522),
            .I(N__32519));
    Odrv4 I__7047 (
            .O(N__32519),
            .I(\ALU.lshift_11 ));
    CascadeMux I__7046 (
            .O(N__32516),
            .I(\ALU.a_15_m4_11_cascade_ ));
    InMux I__7045 (
            .O(N__32513),
            .I(N__32510));
    LocalMux I__7044 (
            .O(N__32510),
            .I(N__32507));
    Span4Mux_h I__7043 (
            .O(N__32507),
            .I(N__32504));
    Odrv4 I__7042 (
            .O(N__32504),
            .I(\ALU.a_15_m3_11 ));
    CascadeMux I__7041 (
            .O(N__32501),
            .I(c_RNID7K8N2_11_cascade_));
    InMux I__7040 (
            .O(N__32498),
            .I(N__32495));
    LocalMux I__7039 (
            .O(N__32495),
            .I(un2_addsub_cry_10_c_RNIEBKOT));
    CascadeMux I__7038 (
            .O(N__32492),
            .I(aluOperation_RNI5QD2L3_0_cascade_));
    InMux I__7037 (
            .O(N__32489),
            .I(N__32486));
    LocalMux I__7036 (
            .O(N__32486),
            .I(N__32483));
    Span4Mux_v I__7035 (
            .O(N__32483),
            .I(N__32479));
    InMux I__7034 (
            .O(N__32482),
            .I(N__32476));
    Span4Mux_h I__7033 (
            .O(N__32479),
            .I(N__32471));
    LocalMux I__7032 (
            .O(N__32476),
            .I(N__32471));
    Odrv4 I__7031 (
            .O(N__32471),
            .I(\ALU.aZ0Z_11 ));
    CEMux I__7030 (
            .O(N__32468),
            .I(N__32464));
    CEMux I__7029 (
            .O(N__32467),
            .I(N__32461));
    LocalMux I__7028 (
            .O(N__32464),
            .I(N__32458));
    LocalMux I__7027 (
            .O(N__32461),
            .I(N__32454));
    Span4Mux_v I__7026 (
            .O(N__32458),
            .I(N__32451));
    CEMux I__7025 (
            .O(N__32457),
            .I(N__32448));
    Span4Mux_v I__7024 (
            .O(N__32454),
            .I(N__32445));
    Span4Mux_v I__7023 (
            .O(N__32451),
            .I(N__32439));
    LocalMux I__7022 (
            .O(N__32448),
            .I(N__32439));
    Span4Mux_h I__7021 (
            .O(N__32445),
            .I(N__32436));
    CEMux I__7020 (
            .O(N__32444),
            .I(N__32432));
    Span4Mux_h I__7019 (
            .O(N__32439),
            .I(N__32429));
    Span4Mux_v I__7018 (
            .O(N__32436),
            .I(N__32426));
    CEMux I__7017 (
            .O(N__32435),
            .I(N__32423));
    LocalMux I__7016 (
            .O(N__32432),
            .I(N__32420));
    Span4Mux_h I__7015 (
            .O(N__32429),
            .I(N__32417));
    Span4Mux_v I__7014 (
            .O(N__32426),
            .I(N__32414));
    LocalMux I__7013 (
            .O(N__32423),
            .I(N__32411));
    Span4Mux_h I__7012 (
            .O(N__32420),
            .I(N__32408));
    Span4Mux_v I__7011 (
            .O(N__32417),
            .I(N__32405));
    IoSpan4Mux I__7010 (
            .O(N__32414),
            .I(N__32402));
    Span4Mux_v I__7009 (
            .O(N__32411),
            .I(N__32399));
    Sp12to4 I__7008 (
            .O(N__32408),
            .I(N__32396));
    Span4Mux_v I__7007 (
            .O(N__32405),
            .I(N__32393));
    Span4Mux_s1_v I__7006 (
            .O(N__32402),
            .I(N__32390));
    Span4Mux_h I__7005 (
            .O(N__32399),
            .I(N__32387));
    Span12Mux_s10_h I__7004 (
            .O(N__32396),
            .I(N__32384));
    Span4Mux_h I__7003 (
            .O(N__32393),
            .I(N__32379));
    Span4Mux_h I__7002 (
            .O(N__32390),
            .I(N__32379));
    Span4Mux_h I__7001 (
            .O(N__32387),
            .I(N__32376));
    Span12Mux_v I__7000 (
            .O(N__32384),
            .I(N__32373));
    Span4Mux_h I__6999 (
            .O(N__32379),
            .I(N__32370));
    Odrv4 I__6998 (
            .O(N__32376),
            .I(\ALU.e_cnvZ0Z_0 ));
    Odrv12 I__6997 (
            .O(N__32373),
            .I(\ALU.e_cnvZ0Z_0 ));
    Odrv4 I__6996 (
            .O(N__32370),
            .I(\ALU.e_cnvZ0Z_0 ));
    InMux I__6995 (
            .O(N__32363),
            .I(N__32359));
    IoInMux I__6994 (
            .O(N__32362),
            .I(N__32356));
    LocalMux I__6993 (
            .O(N__32359),
            .I(N__32353));
    LocalMux I__6992 (
            .O(N__32356),
            .I(N__32350));
    Span4Mux_h I__6991 (
            .O(N__32353),
            .I(N__32347));
    Span4Mux_s3_v I__6990 (
            .O(N__32350),
            .I(N__32344));
    Sp12to4 I__6989 (
            .O(N__32347),
            .I(N__32341));
    Span4Mux_h I__6988 (
            .O(N__32344),
            .I(N__32338));
    Span12Mux_s10_v I__6987 (
            .O(N__32341),
            .I(N__32335));
    Sp12to4 I__6986 (
            .O(N__32338),
            .I(N__32332));
    Odrv12 I__6985 (
            .O(N__32335),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6984 (
            .O(N__32332),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__6983 (
            .O(N__32327),
            .I(N__32323));
    InMux I__6982 (
            .O(N__32326),
            .I(N__32316));
    InMux I__6981 (
            .O(N__32323),
            .I(N__32313));
    InMux I__6980 (
            .O(N__32322),
            .I(N__32308));
    InMux I__6979 (
            .O(N__32321),
            .I(N__32308));
    InMux I__6978 (
            .O(N__32320),
            .I(N__32303));
    InMux I__6977 (
            .O(N__32319),
            .I(N__32303));
    LocalMux I__6976 (
            .O(N__32316),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__6975 (
            .O(N__32313),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__6974 (
            .O(N__32308),
            .I(\FTDI.un3_TX_0 ));
    LocalMux I__6973 (
            .O(N__32303),
            .I(\FTDI.un3_TX_0 ));
    InMux I__6972 (
            .O(N__32294),
            .I(N__32288));
    InMux I__6971 (
            .O(N__32293),
            .I(N__32285));
    InMux I__6970 (
            .O(N__32292),
            .I(N__32282));
    CascadeMux I__6969 (
            .O(N__32291),
            .I(N__32279));
    LocalMux I__6968 (
            .O(N__32288),
            .I(N__32276));
    LocalMux I__6967 (
            .O(N__32285),
            .I(N__32273));
    LocalMux I__6966 (
            .O(N__32282),
            .I(N__32270));
    InMux I__6965 (
            .O(N__32279),
            .I(N__32267));
    Span4Mux_v I__6964 (
            .O(N__32276),
            .I(N__32263));
    Span4Mux_v I__6963 (
            .O(N__32273),
            .I(N__32260));
    Span4Mux_h I__6962 (
            .O(N__32270),
            .I(N__32257));
    LocalMux I__6961 (
            .O(N__32267),
            .I(N__32254));
    InMux I__6960 (
            .O(N__32266),
            .I(N__32251));
    Sp12to4 I__6959 (
            .O(N__32263),
            .I(N__32248));
    Span4Mux_h I__6958 (
            .O(N__32260),
            .I(N__32245));
    Span4Mux_v I__6957 (
            .O(N__32257),
            .I(N__32242));
    Span4Mux_v I__6956 (
            .O(N__32254),
            .I(N__32239));
    LocalMux I__6955 (
            .O(N__32251),
            .I(RXbuffer_4));
    Odrv12 I__6954 (
            .O(N__32248),
            .I(RXbuffer_4));
    Odrv4 I__6953 (
            .O(N__32245),
            .I(RXbuffer_4));
    Odrv4 I__6952 (
            .O(N__32242),
            .I(RXbuffer_4));
    Odrv4 I__6951 (
            .O(N__32239),
            .I(RXbuffer_4));
    InMux I__6950 (
            .O(N__32228),
            .I(N__32225));
    LocalMux I__6949 (
            .O(N__32225),
            .I(N__32221));
    InMux I__6948 (
            .O(N__32224),
            .I(N__32218));
    Span4Mux_v I__6947 (
            .O(N__32221),
            .I(N__32215));
    LocalMux I__6946 (
            .O(N__32218),
            .I(N__32210));
    Span4Mux_h I__6945 (
            .O(N__32215),
            .I(N__32207));
    InMux I__6944 (
            .O(N__32214),
            .I(N__32204));
    InMux I__6943 (
            .O(N__32213),
            .I(N__32201));
    Span4Mux_v I__6942 (
            .O(N__32210),
            .I(N__32198));
    Span4Mux_h I__6941 (
            .O(N__32207),
            .I(N__32193));
    LocalMux I__6940 (
            .O(N__32204),
            .I(N__32193));
    LocalMux I__6939 (
            .O(N__32201),
            .I(N__32188));
    Span4Mux_v I__6938 (
            .O(N__32198),
            .I(N__32188));
    Span4Mux_v I__6937 (
            .O(N__32193),
            .I(N__32185));
    Span4Mux_v I__6936 (
            .O(N__32188),
            .I(N__32181));
    Span4Mux_h I__6935 (
            .O(N__32185),
            .I(N__32178));
    CascadeMux I__6934 (
            .O(N__32184),
            .I(N__32175));
    Span4Mux_h I__6933 (
            .O(N__32181),
            .I(N__32172));
    Span4Mux_h I__6932 (
            .O(N__32178),
            .I(N__32169));
    InMux I__6931 (
            .O(N__32175),
            .I(N__32166));
    Span4Mux_h I__6930 (
            .O(N__32172),
            .I(N__32163));
    Span4Mux_v I__6929 (
            .O(N__32169),
            .I(N__32160));
    LocalMux I__6928 (
            .O(N__32166),
            .I(testWordZ0Z_12));
    Odrv4 I__6927 (
            .O(N__32163),
            .I(testWordZ0Z_12));
    Odrv4 I__6926 (
            .O(N__32160),
            .I(testWordZ0Z_12));
    InMux I__6925 (
            .O(N__32153),
            .I(N__32150));
    LocalMux I__6924 (
            .O(N__32150),
            .I(N__32147));
    Odrv4 I__6923 (
            .O(N__32147),
            .I(TXbufferZ0Z_0));
    InMux I__6922 (
            .O(N__32144),
            .I(N__32141));
    LocalMux I__6921 (
            .O(N__32141),
            .I(N__32138));
    Odrv4 I__6920 (
            .O(N__32138),
            .I(TXbufferZ0Z_3));
    InMux I__6919 (
            .O(N__32135),
            .I(N__32132));
    LocalMux I__6918 (
            .O(N__32132),
            .I(\FTDI.TXshiftZ0Z_5 ));
    InMux I__6917 (
            .O(N__32129),
            .I(N__32126));
    LocalMux I__6916 (
            .O(N__32126),
            .I(N__32123));
    Odrv12 I__6915 (
            .O(N__32123),
            .I(TXbufferZ0Z_4));
    InMux I__6914 (
            .O(N__32120),
            .I(N__32117));
    LocalMux I__6913 (
            .O(N__32117),
            .I(N__32114));
    Odrv4 I__6912 (
            .O(N__32114),
            .I(\FTDI.TXshiftZ0Z_4 ));
    InMux I__6911 (
            .O(N__32111),
            .I(N__32108));
    LocalMux I__6910 (
            .O(N__32108),
            .I(\FTDI.TXshiftZ0Z_3 ));
    InMux I__6909 (
            .O(N__32105),
            .I(N__32102));
    LocalMux I__6908 (
            .O(N__32102),
            .I(N__32099));
    Odrv4 I__6907 (
            .O(N__32099),
            .I(TXbufferZ0Z_2));
    InMux I__6906 (
            .O(N__32096),
            .I(N__32093));
    LocalMux I__6905 (
            .O(N__32093),
            .I(N__32090));
    Odrv4 I__6904 (
            .O(N__32090),
            .I(TXbufferZ0Z_6));
    InMux I__6903 (
            .O(N__32087),
            .I(N__32084));
    LocalMux I__6902 (
            .O(N__32084),
            .I(\FTDI.TXshiftZ0Z_6 ));
    InMux I__6901 (
            .O(N__32081),
            .I(N__32074));
    InMux I__6900 (
            .O(N__32080),
            .I(N__32074));
    InMux I__6899 (
            .O(N__32079),
            .I(N__32070));
    LocalMux I__6898 (
            .O(N__32074),
            .I(N__32062));
    InMux I__6897 (
            .O(N__32073),
            .I(N__32059));
    LocalMux I__6896 (
            .O(N__32070),
            .I(N__32056));
    InMux I__6895 (
            .O(N__32069),
            .I(N__32053));
    InMux I__6894 (
            .O(N__32068),
            .I(N__32050));
    InMux I__6893 (
            .O(N__32067),
            .I(N__32044));
    InMux I__6892 (
            .O(N__32066),
            .I(N__32044));
    CascadeMux I__6891 (
            .O(N__32065),
            .I(N__32041));
    Span4Mux_v I__6890 (
            .O(N__32062),
            .I(N__32036));
    LocalMux I__6889 (
            .O(N__32059),
            .I(N__32033));
    Span4Mux_h I__6888 (
            .O(N__32056),
            .I(N__32028));
    LocalMux I__6887 (
            .O(N__32053),
            .I(N__32028));
    LocalMux I__6886 (
            .O(N__32050),
            .I(N__32022));
    InMux I__6885 (
            .O(N__32049),
            .I(N__32019));
    LocalMux I__6884 (
            .O(N__32044),
            .I(N__32016));
    InMux I__6883 (
            .O(N__32041),
            .I(N__32011));
    InMux I__6882 (
            .O(N__32040),
            .I(N__32006));
    InMux I__6881 (
            .O(N__32039),
            .I(N__32006));
    Span4Mux_h I__6880 (
            .O(N__32036),
            .I(N__31999));
    Span4Mux_v I__6879 (
            .O(N__32033),
            .I(N__31999));
    Span4Mux_h I__6878 (
            .O(N__32028),
            .I(N__31999));
    InMux I__6877 (
            .O(N__32027),
            .I(N__31992));
    InMux I__6876 (
            .O(N__32026),
            .I(N__31992));
    InMux I__6875 (
            .O(N__32025),
            .I(N__31992));
    Sp12to4 I__6874 (
            .O(N__32022),
            .I(N__31987));
    LocalMux I__6873 (
            .O(N__32019),
            .I(N__31987));
    Span4Mux_v I__6872 (
            .O(N__32016),
            .I(N__31984));
    InMux I__6871 (
            .O(N__32015),
            .I(N__31979));
    InMux I__6870 (
            .O(N__32014),
            .I(N__31979));
    LocalMux I__6869 (
            .O(N__32011),
            .I(aluOperand2_2_rep1));
    LocalMux I__6868 (
            .O(N__32006),
            .I(aluOperand2_2_rep1));
    Odrv4 I__6867 (
            .O(N__31999),
            .I(aluOperand2_2_rep1));
    LocalMux I__6866 (
            .O(N__31992),
            .I(aluOperand2_2_rep1));
    Odrv12 I__6865 (
            .O(N__31987),
            .I(aluOperand2_2_rep1));
    Odrv4 I__6864 (
            .O(N__31984),
            .I(aluOperand2_2_rep1));
    LocalMux I__6863 (
            .O(N__31979),
            .I(aluOperand2_2_rep1));
    InMux I__6862 (
            .O(N__31964),
            .I(N__31960));
    InMux I__6861 (
            .O(N__31963),
            .I(N__31957));
    LocalMux I__6860 (
            .O(N__31960),
            .I(N__31954));
    LocalMux I__6859 (
            .O(N__31957),
            .I(\ALU.bZ0Z_2 ));
    Odrv4 I__6858 (
            .O(N__31954),
            .I(\ALU.bZ0Z_2 ));
    InMux I__6857 (
            .O(N__31949),
            .I(N__31946));
    LocalMux I__6856 (
            .O(N__31946),
            .I(\ALU.f_RNIESEJZ0Z_2 ));
    InMux I__6855 (
            .O(N__31943),
            .I(N__31940));
    LocalMux I__6854 (
            .O(N__31940),
            .I(N__31937));
    Span4Mux_h I__6853 (
            .O(N__31937),
            .I(N__31934));
    Span4Mux_h I__6852 (
            .O(N__31934),
            .I(N__31930));
    InMux I__6851 (
            .O(N__31933),
            .I(N__31927));
    Odrv4 I__6850 (
            .O(N__31930),
            .I(\ALU.gZ0Z_0 ));
    LocalMux I__6849 (
            .O(N__31927),
            .I(\ALU.gZ0Z_0 ));
    CascadeMux I__6848 (
            .O(N__31922),
            .I(N__31918));
    InMux I__6847 (
            .O(N__31921),
            .I(N__31915));
    InMux I__6846 (
            .O(N__31918),
            .I(N__31912));
    LocalMux I__6845 (
            .O(N__31915),
            .I(N__31909));
    LocalMux I__6844 (
            .O(N__31912),
            .I(N__31906));
    Odrv4 I__6843 (
            .O(N__31909),
            .I(\ALU.gZ0Z_1 ));
    Odrv12 I__6842 (
            .O(N__31906),
            .I(\ALU.gZ0Z_1 ));
    InMux I__6841 (
            .O(N__31901),
            .I(N__31898));
    LocalMux I__6840 (
            .O(N__31898),
            .I(N__31895));
    Span4Mux_h I__6839 (
            .O(N__31895),
            .I(N__31891));
    InMux I__6838 (
            .O(N__31894),
            .I(N__31888));
    Odrv4 I__6837 (
            .O(N__31891),
            .I(\ALU.gZ0Z_2 ));
    LocalMux I__6836 (
            .O(N__31888),
            .I(\ALU.gZ0Z_2 ));
    InMux I__6835 (
            .O(N__31883),
            .I(N__31880));
    LocalMux I__6834 (
            .O(N__31880),
            .I(N__31876));
    InMux I__6833 (
            .O(N__31879),
            .I(N__31873));
    Span4Mux_h I__6832 (
            .O(N__31876),
            .I(N__31870));
    LocalMux I__6831 (
            .O(N__31873),
            .I(N__31867));
    Odrv4 I__6830 (
            .O(N__31870),
            .I(\ALU.gZ0Z_3 ));
    Odrv12 I__6829 (
            .O(N__31867),
            .I(\ALU.gZ0Z_3 ));
    InMux I__6828 (
            .O(N__31862),
            .I(N__31858));
    InMux I__6827 (
            .O(N__31861),
            .I(N__31855));
    LocalMux I__6826 (
            .O(N__31858),
            .I(N__31852));
    LocalMux I__6825 (
            .O(N__31855),
            .I(N__31849));
    Span4Mux_h I__6824 (
            .O(N__31852),
            .I(N__31846));
    Span4Mux_v I__6823 (
            .O(N__31849),
            .I(N__31843));
    Span4Mux_h I__6822 (
            .O(N__31846),
            .I(N__31840));
    Odrv4 I__6821 (
            .O(N__31843),
            .I(\ALU.gZ0Z_4 ));
    Odrv4 I__6820 (
            .O(N__31840),
            .I(\ALU.gZ0Z_4 ));
    InMux I__6819 (
            .O(N__31835),
            .I(N__31832));
    LocalMux I__6818 (
            .O(N__31832),
            .I(N__31829));
    Span4Mux_v I__6817 (
            .O(N__31829),
            .I(N__31826));
    Span4Mux_h I__6816 (
            .O(N__31826),
            .I(N__31822));
    InMux I__6815 (
            .O(N__31825),
            .I(N__31819));
    Odrv4 I__6814 (
            .O(N__31822),
            .I(\ALU.gZ0Z_5 ));
    LocalMux I__6813 (
            .O(N__31819),
            .I(\ALU.gZ0Z_5 ));
    InMux I__6812 (
            .O(N__31814),
            .I(N__31811));
    LocalMux I__6811 (
            .O(N__31811),
            .I(N__31808));
    Span4Mux_h I__6810 (
            .O(N__31808),
            .I(N__31804));
    InMux I__6809 (
            .O(N__31807),
            .I(N__31801));
    Span4Mux_h I__6808 (
            .O(N__31804),
            .I(N__31798));
    LocalMux I__6807 (
            .O(N__31801),
            .I(N__31795));
    Odrv4 I__6806 (
            .O(N__31798),
            .I(\ALU.gZ0Z_7 ));
    Odrv4 I__6805 (
            .O(N__31795),
            .I(\ALU.gZ0Z_7 ));
    InMux I__6804 (
            .O(N__31790),
            .I(N__31787));
    LocalMux I__6803 (
            .O(N__31787),
            .I(N__31784));
    Span4Mux_h I__6802 (
            .O(N__31784),
            .I(N__31780));
    InMux I__6801 (
            .O(N__31783),
            .I(N__31777));
    Odrv4 I__6800 (
            .O(N__31780),
            .I(\ALU.N_578 ));
    LocalMux I__6799 (
            .O(N__31777),
            .I(\ALU.N_578 ));
    InMux I__6798 (
            .O(N__31772),
            .I(N__31768));
    InMux I__6797 (
            .O(N__31771),
            .I(N__31764));
    LocalMux I__6796 (
            .O(N__31768),
            .I(N__31761));
    InMux I__6795 (
            .O(N__31767),
            .I(N__31758));
    LocalMux I__6794 (
            .O(N__31764),
            .I(\ALU.N_477 ));
    Odrv12 I__6793 (
            .O(N__31761),
            .I(\ALU.N_477 ));
    LocalMux I__6792 (
            .O(N__31758),
            .I(\ALU.N_477 ));
    InMux I__6791 (
            .O(N__31751),
            .I(N__31748));
    LocalMux I__6790 (
            .O(N__31748),
            .I(\ALU.N_634 ));
    InMux I__6789 (
            .O(N__31745),
            .I(N__31742));
    LocalMux I__6788 (
            .O(N__31742),
            .I(N__31738));
    InMux I__6787 (
            .O(N__31741),
            .I(N__31735));
    Span4Mux_h I__6786 (
            .O(N__31738),
            .I(N__31732));
    LocalMux I__6785 (
            .O(N__31735),
            .I(N__31729));
    Odrv4 I__6784 (
            .O(N__31732),
            .I(\ALU.aZ0Z_15 ));
    Odrv4 I__6783 (
            .O(N__31729),
            .I(\ALU.aZ0Z_15 ));
    InMux I__6782 (
            .O(N__31724),
            .I(N__31721));
    LocalMux I__6781 (
            .O(N__31721),
            .I(N__31718));
    Span4Mux_v I__6780 (
            .O(N__31718),
            .I(N__31715));
    Span4Mux_h I__6779 (
            .O(N__31715),
            .I(N__31712));
    Odrv4 I__6778 (
            .O(N__31712),
            .I(\ALU.f_RNI0P6LZ0Z_1 ));
    InMux I__6777 (
            .O(N__31709),
            .I(N__31706));
    LocalMux I__6776 (
            .O(N__31706),
            .I(N__31703));
    Span4Mux_h I__6775 (
            .O(N__31703),
            .I(N__31700));
    Span4Mux_h I__6774 (
            .O(N__31700),
            .I(N__31697));
    Odrv4 I__6773 (
            .O(N__31697),
            .I(\ALU.f_RNICQEJZ0Z_1 ));
    InMux I__6772 (
            .O(N__31694),
            .I(N__31691));
    LocalMux I__6771 (
            .O(N__31691),
            .I(N__31687));
    InMux I__6770 (
            .O(N__31690),
            .I(N__31684));
    Span4Mux_v I__6769 (
            .O(N__31687),
            .I(N__31681));
    LocalMux I__6768 (
            .O(N__31684),
            .I(N__31678));
    Span4Mux_h I__6767 (
            .O(N__31681),
            .I(N__31673));
    Span4Mux_h I__6766 (
            .O(N__31678),
            .I(N__31673));
    Odrv4 I__6765 (
            .O(N__31673),
            .I(\ALU.cZ0Z_7 ));
    InMux I__6764 (
            .O(N__31670),
            .I(N__31667));
    LocalMux I__6763 (
            .O(N__31667),
            .I(N__31664));
    Span4Mux_h I__6762 (
            .O(N__31664),
            .I(N__31661));
    Span4Mux_h I__6761 (
            .O(N__31661),
            .I(N__31658));
    Odrv4 I__6760 (
            .O(N__31658),
            .I(\ALU.g_RNIQCLLZ0Z_7 ));
    InMux I__6759 (
            .O(N__31655),
            .I(N__31652));
    LocalMux I__6758 (
            .O(N__31652),
            .I(N__31649));
    Odrv12 I__6757 (
            .O(N__31649),
            .I(\ALU.f_RNIL2FJZ0Z_5 ));
    InMux I__6756 (
            .O(N__31646),
            .I(N__31643));
    LocalMux I__6755 (
            .O(N__31643),
            .I(N__31640));
    Span4Mux_v I__6754 (
            .O(N__31640),
            .I(N__31637));
    Span4Mux_h I__6753 (
            .O(N__31637),
            .I(N__31634));
    Span4Mux_v I__6752 (
            .O(N__31634),
            .I(N__31631));
    Odrv4 I__6751 (
            .O(N__31631),
            .I(\ALU.m286_bmZ0 ));
    InMux I__6750 (
            .O(N__31628),
            .I(N__31625));
    LocalMux I__6749 (
            .O(N__31625),
            .I(N__31622));
    Span4Mux_v I__6748 (
            .O(N__31622),
            .I(N__31619));
    Span4Mux_h I__6747 (
            .O(N__31619),
            .I(N__31616));
    Span4Mux_v I__6746 (
            .O(N__31616),
            .I(N__31613));
    Span4Mux_v I__6745 (
            .O(N__31613),
            .I(N__31610));
    Odrv4 I__6744 (
            .O(N__31610),
            .I(\ALU.m286_amZ0 ));
    InMux I__6743 (
            .O(N__31607),
            .I(N__31604));
    LocalMux I__6742 (
            .O(N__31604),
            .I(N__31601));
    Odrv12 I__6741 (
            .O(N__31601),
            .I(\ALU.f_RNIAOEJZ0Z_0 ));
    InMux I__6740 (
            .O(N__31598),
            .I(N__31594));
    InMux I__6739 (
            .O(N__31597),
            .I(N__31590));
    LocalMux I__6738 (
            .O(N__31594),
            .I(N__31587));
    CascadeMux I__6737 (
            .O(N__31593),
            .I(N__31584));
    LocalMux I__6736 (
            .O(N__31590),
            .I(N__31581));
    Span4Mux_h I__6735 (
            .O(N__31587),
            .I(N__31578));
    InMux I__6734 (
            .O(N__31584),
            .I(N__31574));
    Span4Mux_h I__6733 (
            .O(N__31581),
            .I(N__31571));
    Span4Mux_h I__6732 (
            .O(N__31578),
            .I(N__31568));
    InMux I__6731 (
            .O(N__31577),
            .I(N__31565));
    LocalMux I__6730 (
            .O(N__31574),
            .I(aluOperand2_fast_0));
    Odrv4 I__6729 (
            .O(N__31571),
            .I(aluOperand2_fast_0));
    Odrv4 I__6728 (
            .O(N__31568),
            .I(aluOperand2_fast_0));
    LocalMux I__6727 (
            .O(N__31565),
            .I(aluOperand2_fast_0));
    InMux I__6726 (
            .O(N__31556),
            .I(N__31553));
    LocalMux I__6725 (
            .O(N__31553),
            .I(N__31550));
    Span4Mux_h I__6724 (
            .O(N__31550),
            .I(N__31547));
    Span4Mux_v I__6723 (
            .O(N__31547),
            .I(N__31544));
    Span4Mux_h I__6722 (
            .O(N__31544),
            .I(N__31540));
    InMux I__6721 (
            .O(N__31543),
            .I(N__31537));
    Odrv4 I__6720 (
            .O(N__31540),
            .I(\ALU.cZ0Z_14 ));
    LocalMux I__6719 (
            .O(N__31537),
            .I(\ALU.cZ0Z_14 ));
    InMux I__6718 (
            .O(N__31532),
            .I(N__31529));
    LocalMux I__6717 (
            .O(N__31529),
            .I(N__31526));
    Odrv12 I__6716 (
            .O(N__31526),
            .I(\ALU.c_RNIND49Z0Z_14 ));
    InMux I__6715 (
            .O(N__31523),
            .I(N__31519));
    InMux I__6714 (
            .O(N__31522),
            .I(N__31516));
    LocalMux I__6713 (
            .O(N__31519),
            .I(N__31513));
    LocalMux I__6712 (
            .O(N__31516),
            .I(N__31510));
    Span4Mux_h I__6711 (
            .O(N__31513),
            .I(N__31507));
    Odrv4 I__6710 (
            .O(N__31510),
            .I(\ALU.cZ0Z_15 ));
    Odrv4 I__6709 (
            .O(N__31507),
            .I(\ALU.cZ0Z_15 ));
    CEMux I__6708 (
            .O(N__31502),
            .I(N__31499));
    LocalMux I__6707 (
            .O(N__31499),
            .I(N__31494));
    CEMux I__6706 (
            .O(N__31498),
            .I(N__31491));
    CEMux I__6705 (
            .O(N__31497),
            .I(N__31488));
    Span4Mux_h I__6704 (
            .O(N__31494),
            .I(N__31485));
    LocalMux I__6703 (
            .O(N__31491),
            .I(N__31482));
    LocalMux I__6702 (
            .O(N__31488),
            .I(N__31479));
    Span4Mux_v I__6701 (
            .O(N__31485),
            .I(N__31476));
    Span4Mux_s1_v I__6700 (
            .O(N__31482),
            .I(N__31473));
    Span4Mux_h I__6699 (
            .O(N__31479),
            .I(N__31470));
    Span4Mux_v I__6698 (
            .O(N__31476),
            .I(N__31467));
    Span4Mux_v I__6697 (
            .O(N__31473),
            .I(N__31464));
    Span4Mux_v I__6696 (
            .O(N__31470),
            .I(N__31461));
    Span4Mux_v I__6695 (
            .O(N__31467),
            .I(N__31458));
    Span4Mux_h I__6694 (
            .O(N__31464),
            .I(N__31455));
    Span4Mux_v I__6693 (
            .O(N__31461),
            .I(N__31452));
    Span4Mux_h I__6692 (
            .O(N__31458),
            .I(N__31449));
    Odrv4 I__6691 (
            .O(N__31455),
            .I(\ALU.c_cnvZ0Z_0 ));
    Odrv4 I__6690 (
            .O(N__31452),
            .I(\ALU.c_cnvZ0Z_0 ));
    Odrv4 I__6689 (
            .O(N__31449),
            .I(\ALU.c_cnvZ0Z_0 ));
    InMux I__6688 (
            .O(N__31442),
            .I(N__31436));
    InMux I__6687 (
            .O(N__31441),
            .I(N__31436));
    LocalMux I__6686 (
            .O(N__31436),
            .I(N__31433));
    Span4Mux_v I__6685 (
            .O(N__31433),
            .I(N__31430));
    Odrv4 I__6684 (
            .O(N__31430),
            .I(\ALU.hZ0Z_1 ));
    InMux I__6683 (
            .O(N__31427),
            .I(N__31424));
    LocalMux I__6682 (
            .O(N__31424),
            .I(N__31420));
    InMux I__6681 (
            .O(N__31423),
            .I(N__31417));
    Span4Mux_h I__6680 (
            .O(N__31420),
            .I(N__31412));
    LocalMux I__6679 (
            .O(N__31417),
            .I(N__31412));
    Span4Mux_v I__6678 (
            .O(N__31412),
            .I(N__31409));
    Odrv4 I__6677 (
            .O(N__31409),
            .I(\ALU.hZ0Z_2 ));
    InMux I__6676 (
            .O(N__31406),
            .I(N__31403));
    LocalMux I__6675 (
            .O(N__31403),
            .I(N__31400));
    Span4Mux_h I__6674 (
            .O(N__31400),
            .I(N__31397));
    Span4Mux_v I__6673 (
            .O(N__31397),
            .I(N__31393));
    InMux I__6672 (
            .O(N__31396),
            .I(N__31390));
    Odrv4 I__6671 (
            .O(N__31393),
            .I(\ALU.hZ0Z_5 ));
    LocalMux I__6670 (
            .O(N__31390),
            .I(\ALU.hZ0Z_5 ));
    InMux I__6669 (
            .O(N__31385),
            .I(N__31382));
    LocalMux I__6668 (
            .O(N__31382),
            .I(N__31379));
    Span4Mux_h I__6667 (
            .O(N__31379),
            .I(N__31375));
    InMux I__6666 (
            .O(N__31378),
            .I(N__31372));
    Span4Mux_h I__6665 (
            .O(N__31375),
            .I(N__31367));
    LocalMux I__6664 (
            .O(N__31372),
            .I(N__31367));
    Span4Mux_v I__6663 (
            .O(N__31367),
            .I(N__31364));
    Odrv4 I__6662 (
            .O(N__31364),
            .I(\ALU.aZ0Z_14 ));
    InMux I__6661 (
            .O(N__31361),
            .I(N__31357));
    InMux I__6660 (
            .O(N__31360),
            .I(N__31354));
    LocalMux I__6659 (
            .O(N__31357),
            .I(\ALU.eZ0Z_15 ));
    LocalMux I__6658 (
            .O(N__31354),
            .I(\ALU.eZ0Z_15 ));
    CascadeMux I__6657 (
            .O(N__31349),
            .I(\ALU.a_RNILVBOZ0Z_15_cascade_ ));
    InMux I__6656 (
            .O(N__31346),
            .I(N__31343));
    LocalMux I__6655 (
            .O(N__31343),
            .I(\ALU.c_RNIPF49Z0Z_15 ));
    CascadeMux I__6654 (
            .O(N__31340),
            .I(\ALU.operand2_7_ns_1_15_cascade_ ));
    InMux I__6653 (
            .O(N__31337),
            .I(N__31334));
    LocalMux I__6652 (
            .O(N__31334),
            .I(N__31331));
    Span4Mux_v I__6651 (
            .O(N__31331),
            .I(N__31328));
    Span4Mux_v I__6650 (
            .O(N__31328),
            .I(N__31325));
    Odrv4 I__6649 (
            .O(N__31325),
            .I(\ALU.b_RNIORSD1Z0Z_15 ));
    InMux I__6648 (
            .O(N__31322),
            .I(N__31319));
    LocalMux I__6647 (
            .O(N__31319),
            .I(N__31316));
    Span4Mux_h I__6646 (
            .O(N__31316),
            .I(N__31313));
    Span4Mux_h I__6645 (
            .O(N__31313),
            .I(N__31310));
    Odrv4 I__6644 (
            .O(N__31310),
            .I(\ALU.operand2_15 ));
    InMux I__6643 (
            .O(N__31307),
            .I(N__31304));
    LocalMux I__6642 (
            .O(N__31304),
            .I(N__31301));
    Span4Mux_v I__6641 (
            .O(N__31301),
            .I(N__31297));
    InMux I__6640 (
            .O(N__31300),
            .I(N__31294));
    Span4Mux_h I__6639 (
            .O(N__31297),
            .I(N__31289));
    LocalMux I__6638 (
            .O(N__31294),
            .I(N__31289));
    Odrv4 I__6637 (
            .O(N__31289),
            .I(\ALU.cZ0Z_11 ));
    InMux I__6636 (
            .O(N__31286),
            .I(N__31283));
    LocalMux I__6635 (
            .O(N__31283),
            .I(N__31279));
    InMux I__6634 (
            .O(N__31282),
            .I(N__31276));
    Span4Mux_h I__6633 (
            .O(N__31279),
            .I(N__31271));
    LocalMux I__6632 (
            .O(N__31276),
            .I(N__31271));
    Span4Mux_h I__6631 (
            .O(N__31271),
            .I(N__31268));
    Odrv4 I__6630 (
            .O(N__31268),
            .I(\ALU.cZ0Z_12 ));
    InMux I__6629 (
            .O(N__31265),
            .I(N__31257));
    InMux I__6628 (
            .O(N__31264),
            .I(N__31254));
    InMux I__6627 (
            .O(N__31263),
            .I(N__31251));
    InMux I__6626 (
            .O(N__31262),
            .I(N__31246));
    InMux I__6625 (
            .O(N__31261),
            .I(N__31243));
    InMux I__6624 (
            .O(N__31260),
            .I(N__31240));
    LocalMux I__6623 (
            .O(N__31257),
            .I(N__31237));
    LocalMux I__6622 (
            .O(N__31254),
            .I(N__31234));
    LocalMux I__6621 (
            .O(N__31251),
            .I(N__31231));
    CascadeMux I__6620 (
            .O(N__31250),
            .I(N__31228));
    InMux I__6619 (
            .O(N__31249),
            .I(N__31225));
    LocalMux I__6618 (
            .O(N__31246),
            .I(N__31212));
    LocalMux I__6617 (
            .O(N__31243),
            .I(N__31212));
    LocalMux I__6616 (
            .O(N__31240),
            .I(N__31212));
    Span4Mux_h I__6615 (
            .O(N__31237),
            .I(N__31212));
    Span4Mux_v I__6614 (
            .O(N__31234),
            .I(N__31212));
    Span4Mux_h I__6613 (
            .O(N__31231),
            .I(N__31212));
    InMux I__6612 (
            .O(N__31228),
            .I(N__31209));
    LocalMux I__6611 (
            .O(N__31225),
            .I(N__31206));
    Span4Mux_v I__6610 (
            .O(N__31212),
            .I(N__31203));
    LocalMux I__6609 (
            .O(N__31209),
            .I(N__31198));
    Span12Mux_h I__6608 (
            .O(N__31206),
            .I(N__31198));
    Odrv4 I__6607 (
            .O(N__31203),
            .I(aluOperand2_0_rep1));
    Odrv12 I__6606 (
            .O(N__31198),
            .I(aluOperand2_0_rep1));
    CascadeMux I__6605 (
            .O(N__31193),
            .I(\ALU.a_RNICNBOZ0Z_11_cascade_ ));
    CascadeMux I__6604 (
            .O(N__31190),
            .I(\ALU.operand2_7_ns_1_11_cascade_ ));
    InMux I__6603 (
            .O(N__31187),
            .I(N__31184));
    LocalMux I__6602 (
            .O(N__31184),
            .I(\ALU.b_RNIGJSD1Z0Z_11 ));
    InMux I__6601 (
            .O(N__31181),
            .I(N__31177));
    CascadeMux I__6600 (
            .O(N__31180),
            .I(N__31174));
    LocalMux I__6599 (
            .O(N__31177),
            .I(N__31171));
    InMux I__6598 (
            .O(N__31174),
            .I(N__31168));
    Span4Mux_h I__6597 (
            .O(N__31171),
            .I(N__31165));
    LocalMux I__6596 (
            .O(N__31168),
            .I(N__31162));
    Odrv4 I__6595 (
            .O(N__31165),
            .I(\ALU.operand2_11 ));
    Odrv12 I__6594 (
            .O(N__31162),
            .I(\ALU.operand2_11 ));
    InMux I__6593 (
            .O(N__31157),
            .I(N__31154));
    LocalMux I__6592 (
            .O(N__31154),
            .I(N__31150));
    InMux I__6591 (
            .O(N__31153),
            .I(N__31147));
    Odrv12 I__6590 (
            .O(N__31150),
            .I(\ALU.dZ0Z_11 ));
    LocalMux I__6589 (
            .O(N__31147),
            .I(\ALU.dZ0Z_11 ));
    InMux I__6588 (
            .O(N__31142),
            .I(N__31139));
    LocalMux I__6587 (
            .O(N__31139),
            .I(\ALU.d_RNIK3LUZ0Z_11 ));
    InMux I__6586 (
            .O(N__31136),
            .I(N__31133));
    LocalMux I__6585 (
            .O(N__31133),
            .I(N__31130));
    Span4Mux_v I__6584 (
            .O(N__31130),
            .I(N__31126));
    InMux I__6583 (
            .O(N__31129),
            .I(N__31123));
    Odrv4 I__6582 (
            .O(N__31126),
            .I(\ALU.hZ0Z_11 ));
    LocalMux I__6581 (
            .O(N__31123),
            .I(\ALU.hZ0Z_11 ));
    InMux I__6580 (
            .O(N__31118),
            .I(N__31115));
    LocalMux I__6579 (
            .O(N__31115),
            .I(\ALU.c_RNIG749Z0Z_11 ));
    CascadeMux I__6578 (
            .O(N__31112),
            .I(\ALU.a_RNIHRBOZ0Z_13_cascade_ ));
    InMux I__6577 (
            .O(N__31109),
            .I(N__31106));
    LocalMux I__6576 (
            .O(N__31106),
            .I(\ALU.c_RNILB49Z0Z_13 ));
    InMux I__6575 (
            .O(N__31103),
            .I(N__31100));
    LocalMux I__6574 (
            .O(N__31100),
            .I(N__31097));
    Span4Mux_v I__6573 (
            .O(N__31097),
            .I(N__31093));
    InMux I__6572 (
            .O(N__31096),
            .I(N__31090));
    Span4Mux_h I__6571 (
            .O(N__31093),
            .I(N__31087));
    LocalMux I__6570 (
            .O(N__31090),
            .I(\ALU.operand2_7_ns_1_13 ));
    Odrv4 I__6569 (
            .O(N__31087),
            .I(\ALU.operand2_7_ns_1_13 ));
    InMux I__6568 (
            .O(N__31082),
            .I(N__31079));
    LocalMux I__6567 (
            .O(N__31079),
            .I(N__31076));
    Span4Mux_h I__6566 (
            .O(N__31076),
            .I(N__31073));
    Span4Mux_h I__6565 (
            .O(N__31073),
            .I(N__31070));
    Odrv4 I__6564 (
            .O(N__31070),
            .I(\ALU.un2_addsub_cry_7_c_RNIL8JHGZ0 ));
    InMux I__6563 (
            .O(N__31067),
            .I(N__31064));
    LocalMux I__6562 (
            .O(N__31064),
            .I(N__31061));
    Span4Mux_h I__6561 (
            .O(N__31061),
            .I(N__31057));
    InMux I__6560 (
            .O(N__31060),
            .I(N__31054));
    Span4Mux_h I__6559 (
            .O(N__31057),
            .I(N__31051));
    LocalMux I__6558 (
            .O(N__31054),
            .I(\ALU.aZ0Z_8 ));
    Odrv4 I__6557 (
            .O(N__31051),
            .I(\ALU.aZ0Z_8 ));
    InMux I__6556 (
            .O(N__31046),
            .I(N__31038));
    CascadeMux I__6555 (
            .O(N__31045),
            .I(N__31035));
    CascadeMux I__6554 (
            .O(N__31044),
            .I(N__31032));
    InMux I__6553 (
            .O(N__31043),
            .I(N__31029));
    InMux I__6552 (
            .O(N__31042),
            .I(N__31026));
    InMux I__6551 (
            .O(N__31041),
            .I(N__31023));
    LocalMux I__6550 (
            .O(N__31038),
            .I(N__31020));
    InMux I__6549 (
            .O(N__31035),
            .I(N__31015));
    InMux I__6548 (
            .O(N__31032),
            .I(N__31015));
    LocalMux I__6547 (
            .O(N__31029),
            .I(N__31010));
    LocalMux I__6546 (
            .O(N__31026),
            .I(N__31007));
    LocalMux I__6545 (
            .O(N__31023),
            .I(N__31004));
    Span4Mux_v I__6544 (
            .O(N__31020),
            .I(N__30999));
    LocalMux I__6543 (
            .O(N__31015),
            .I(N__30999));
    InMux I__6542 (
            .O(N__31014),
            .I(N__30994));
    InMux I__6541 (
            .O(N__31013),
            .I(N__30994));
    Span4Mux_v I__6540 (
            .O(N__31010),
            .I(N__30991));
    Span4Mux_v I__6539 (
            .O(N__31007),
            .I(N__30988));
    Span4Mux_h I__6538 (
            .O(N__31004),
            .I(N__30983));
    Span4Mux_h I__6537 (
            .O(N__30999),
            .I(N__30983));
    LocalMux I__6536 (
            .O(N__30994),
            .I(aluOperand2_fast_1));
    Odrv4 I__6535 (
            .O(N__30991),
            .I(aluOperand2_fast_1));
    Odrv4 I__6534 (
            .O(N__30988),
            .I(aluOperand2_fast_1));
    Odrv4 I__6533 (
            .O(N__30983),
            .I(aluOperand2_fast_1));
    CascadeMux I__6532 (
            .O(N__30974),
            .I(N__30970));
    CascadeMux I__6531 (
            .O(N__30973),
            .I(N__30967));
    InMux I__6530 (
            .O(N__30970),
            .I(N__30964));
    InMux I__6529 (
            .O(N__30967),
            .I(N__30961));
    LocalMux I__6528 (
            .O(N__30964),
            .I(N__30958));
    LocalMux I__6527 (
            .O(N__30961),
            .I(N__30955));
    Span4Mux_v I__6526 (
            .O(N__30958),
            .I(N__30952));
    Span4Mux_v I__6525 (
            .O(N__30955),
            .I(N__30949));
    Span4Mux_h I__6524 (
            .O(N__30952),
            .I(N__30946));
    Odrv4 I__6523 (
            .O(N__30949),
            .I(\ALU.eZ0Z_8 ));
    Odrv4 I__6522 (
            .O(N__30946),
            .I(\ALU.eZ0Z_8 ));
    CascadeMux I__6521 (
            .O(N__30941),
            .I(N__30938));
    InMux I__6520 (
            .O(N__30938),
            .I(N__30934));
    InMux I__6519 (
            .O(N__30937),
            .I(N__30931));
    LocalMux I__6518 (
            .O(N__30934),
            .I(N__30928));
    LocalMux I__6517 (
            .O(N__30931),
            .I(N__30925));
    Span4Mux_h I__6516 (
            .O(N__30928),
            .I(N__30922));
    Span4Mux_v I__6515 (
            .O(N__30925),
            .I(N__30919));
    Span4Mux_v I__6514 (
            .O(N__30922),
            .I(N__30916));
    Sp12to4 I__6513 (
            .O(N__30919),
            .I(N__30913));
    Odrv4 I__6512 (
            .O(N__30916),
            .I(\ALU.gZ0Z_8 ));
    Odrv12 I__6511 (
            .O(N__30913),
            .I(\ALU.gZ0Z_8 ));
    InMux I__6510 (
            .O(N__30908),
            .I(N__30905));
    LocalMux I__6509 (
            .O(N__30905),
            .I(N__30902));
    Span4Mux_h I__6508 (
            .O(N__30902),
            .I(N__30898));
    InMux I__6507 (
            .O(N__30901),
            .I(N__30895));
    Span4Mux_v I__6506 (
            .O(N__30898),
            .I(N__30892));
    LocalMux I__6505 (
            .O(N__30895),
            .I(N__30889));
    Span4Mux_v I__6504 (
            .O(N__30892),
            .I(N__30886));
    Span4Mux_v I__6503 (
            .O(N__30889),
            .I(N__30883));
    Odrv4 I__6502 (
            .O(N__30886),
            .I(\ALU.cZ0Z_8 ));
    Odrv4 I__6501 (
            .O(N__30883),
            .I(\ALU.cZ0Z_8 ));
    CascadeMux I__6500 (
            .O(N__30878),
            .I(\ALU.operand2_3_ns_1_8_cascade_ ));
    InMux I__6499 (
            .O(N__30875),
            .I(N__30872));
    LocalMux I__6498 (
            .O(N__30872),
            .I(N__30869));
    Span4Mux_s3_h I__6497 (
            .O(N__30869),
            .I(N__30866));
    Span4Mux_h I__6496 (
            .O(N__30866),
            .I(N__30863));
    Odrv4 I__6495 (
            .O(N__30863),
            .I(\ALU.N_819 ));
    CascadeMux I__6494 (
            .O(N__30860),
            .I(\ALU.addsub_0_sqmuxa_cascade_ ));
    InMux I__6493 (
            .O(N__30857),
            .I(N__30854));
    LocalMux I__6492 (
            .O(N__30854),
            .I(N__30851));
    Span12Mux_h I__6491 (
            .O(N__30851),
            .I(N__30848));
    Odrv12 I__6490 (
            .O(N__30848),
            .I(\ALU.un2_addsub_cry_8_c_RNIKR81JZ0 ));
    CascadeMux I__6489 (
            .O(N__30845),
            .I(\ALU.un9_addsub_cry_8_c_RNIKTS9SZ0_cascade_ ));
    InMux I__6488 (
            .O(N__30842),
            .I(N__30839));
    LocalMux I__6487 (
            .O(N__30839),
            .I(N__30836));
    Odrv4 I__6486 (
            .O(N__30836),
            .I(\ALU.a_15_m5_9 ));
    CascadeMux I__6485 (
            .O(N__30833),
            .I(\ALU.a_15_ns_1_9_cascade_ ));
    InMux I__6484 (
            .O(N__30830),
            .I(N__30827));
    LocalMux I__6483 (
            .O(N__30827),
            .I(N__30823));
    InMux I__6482 (
            .O(N__30826),
            .I(N__30820));
    Span4Mux_v I__6481 (
            .O(N__30823),
            .I(N__30817));
    LocalMux I__6480 (
            .O(N__30820),
            .I(N__30814));
    Odrv4 I__6479 (
            .O(N__30817),
            .I(\ALU.eZ0Z_11 ));
    Odrv4 I__6478 (
            .O(N__30814),
            .I(\ALU.eZ0Z_11 ));
    CascadeMux I__6477 (
            .O(N__30809),
            .I(N__30802));
    InMux I__6476 (
            .O(N__30808),
            .I(N__30797));
    InMux I__6475 (
            .O(N__30807),
            .I(N__30797));
    InMux I__6474 (
            .O(N__30806),
            .I(N__30794));
    InMux I__6473 (
            .O(N__30805),
            .I(N__30789));
    InMux I__6472 (
            .O(N__30802),
            .I(N__30789));
    LocalMux I__6471 (
            .O(N__30797),
            .I(N__30784));
    LocalMux I__6470 (
            .O(N__30794),
            .I(N__30784));
    LocalMux I__6469 (
            .O(N__30789),
            .I(N__30775));
    Span4Mux_v I__6468 (
            .O(N__30784),
            .I(N__30775));
    CascadeMux I__6467 (
            .O(N__30783),
            .I(N__30772));
    CascadeMux I__6466 (
            .O(N__30782),
            .I(N__30769));
    CascadeMux I__6465 (
            .O(N__30781),
            .I(N__30766));
    CascadeMux I__6464 (
            .O(N__30780),
            .I(N__30763));
    Span4Mux_h I__6463 (
            .O(N__30775),
            .I(N__30760));
    InMux I__6462 (
            .O(N__30772),
            .I(N__30757));
    InMux I__6461 (
            .O(N__30769),
            .I(N__30750));
    InMux I__6460 (
            .O(N__30766),
            .I(N__30750));
    InMux I__6459 (
            .O(N__30763),
            .I(N__30750));
    Odrv4 I__6458 (
            .O(N__30760),
            .I(testStateZ0Z_2));
    LocalMux I__6457 (
            .O(N__30757),
            .I(testStateZ0Z_2));
    LocalMux I__6456 (
            .O(N__30750),
            .I(testStateZ0Z_2));
    IoInMux I__6455 (
            .O(N__30743),
            .I(N__30740));
    LocalMux I__6454 (
            .O(N__30740),
            .I(N__30737));
    Span12Mux_s0_h I__6453 (
            .O(N__30737),
            .I(N__30734));
    Span12Mux_v I__6452 (
            .O(N__30734),
            .I(N__30731));
    Odrv12 I__6451 (
            .O(N__30731),
            .I(testState_i_2));
    InMux I__6450 (
            .O(N__30728),
            .I(N__30725));
    LocalMux I__6449 (
            .O(N__30725),
            .I(N__30722));
    Span4Mux_h I__6448 (
            .O(N__30722),
            .I(N__30718));
    InMux I__6447 (
            .O(N__30721),
            .I(N__30715));
    Span4Mux_h I__6446 (
            .O(N__30718),
            .I(N__30710));
    LocalMux I__6445 (
            .O(N__30715),
            .I(N__30710));
    Span4Mux_v I__6444 (
            .O(N__30710),
            .I(N__30707));
    Odrv4 I__6443 (
            .O(N__30707),
            .I(\ALU.eZ0Z_14 ));
    InMux I__6442 (
            .O(N__30704),
            .I(N__30701));
    LocalMux I__6441 (
            .O(N__30701),
            .I(N__30698));
    Span4Mux_v I__6440 (
            .O(N__30698),
            .I(N__30695));
    Span4Mux_h I__6439 (
            .O(N__30695),
            .I(N__30692));
    Span4Mux_h I__6438 (
            .O(N__30692),
            .I(N__30689));
    Odrv4 I__6437 (
            .O(N__30689),
            .I(\ALU.un2_addsub_cry_13_c_RNINVE5KZ0 ));
    CascadeMux I__6436 (
            .O(N__30686),
            .I(un2_addsub_cry_13_c_RNI2LH1U_cascade_));
    InMux I__6435 (
            .O(N__30683),
            .I(N__30680));
    LocalMux I__6434 (
            .O(N__30680),
            .I(N__30677));
    Span4Mux_v I__6433 (
            .O(N__30677),
            .I(N__30674));
    Span4Mux_h I__6432 (
            .O(N__30674),
            .I(N__30671));
    Odrv4 I__6431 (
            .O(N__30671),
            .I(c_RNIFCGVL2_14));
    CascadeMux I__6430 (
            .O(N__30668),
            .I(aluOperation_RNIR872K3_0_cascade_));
    CascadeMux I__6429 (
            .O(N__30665),
            .I(N__30662));
    InMux I__6428 (
            .O(N__30662),
            .I(N__30659));
    LocalMux I__6427 (
            .O(N__30659),
            .I(\ALU.a_RNIJTBOZ0Z_14 ));
    CascadeMux I__6426 (
            .O(N__30656),
            .I(\ALU.operand2_7_ns_1_14_cascade_ ));
    InMux I__6425 (
            .O(N__30653),
            .I(N__30650));
    LocalMux I__6424 (
            .O(N__30650),
            .I(\ALU.b_RNIMPSD1Z0Z_14 ));
    CascadeMux I__6423 (
            .O(N__30647),
            .I(N__30643));
    CascadeMux I__6422 (
            .O(N__30646),
            .I(N__30640));
    InMux I__6421 (
            .O(N__30643),
            .I(N__30635));
    InMux I__6420 (
            .O(N__30640),
            .I(N__30635));
    LocalMux I__6419 (
            .O(N__30635),
            .I(N__30631));
    InMux I__6418 (
            .O(N__30634),
            .I(N__30628));
    Span12Mux_s5_v I__6417 (
            .O(N__30631),
            .I(N__30623));
    LocalMux I__6416 (
            .O(N__30628),
            .I(N__30623));
    Odrv12 I__6415 (
            .O(N__30623),
            .I(\ALU.operand2_14 ));
    InMux I__6414 (
            .O(N__30620),
            .I(N__30617));
    LocalMux I__6413 (
            .O(N__30617),
            .I(N__30614));
    Span4Mux_v I__6412 (
            .O(N__30614),
            .I(N__30611));
    Span4Mux_s3_h I__6411 (
            .O(N__30611),
            .I(N__30607));
    InMux I__6410 (
            .O(N__30610),
            .I(N__30604));
    Span4Mux_h I__6409 (
            .O(N__30607),
            .I(N__30601));
    LocalMux I__6408 (
            .O(N__30604),
            .I(\ALU.hZ0Z_14 ));
    Odrv4 I__6407 (
            .O(N__30601),
            .I(\ALU.hZ0Z_14 ));
    InMux I__6406 (
            .O(N__30596),
            .I(N__30593));
    LocalMux I__6405 (
            .O(N__30593),
            .I(N__30590));
    Span4Mux_h I__6404 (
            .O(N__30590),
            .I(N__30586));
    InMux I__6403 (
            .O(N__30589),
            .I(N__30583));
    Span4Mux_h I__6402 (
            .O(N__30586),
            .I(N__30580));
    LocalMux I__6401 (
            .O(N__30583),
            .I(N__30577));
    Span4Mux_v I__6400 (
            .O(N__30580),
            .I(N__30574));
    Span4Mux_h I__6399 (
            .O(N__30577),
            .I(N__30571));
    Odrv4 I__6398 (
            .O(N__30574),
            .I(\ALU.dZ0Z_14 ));
    Odrv4 I__6397 (
            .O(N__30571),
            .I(\ALU.dZ0Z_14 ));
    InMux I__6396 (
            .O(N__30566),
            .I(N__30563));
    LocalMux I__6395 (
            .O(N__30563),
            .I(\ALU.d_RNIQ9LUZ0Z_14 ));
    CascadeMux I__6394 (
            .O(N__30560),
            .I(\ALU.c_RNI1OCN4Z0Z_15_cascade_ ));
    InMux I__6393 (
            .O(N__30557),
            .I(N__30553));
    InMux I__6392 (
            .O(N__30556),
            .I(N__30550));
    LocalMux I__6391 (
            .O(N__30553),
            .I(N__30547));
    LocalMux I__6390 (
            .O(N__30550),
            .I(N__30544));
    Span12Mux_h I__6389 (
            .O(N__30547),
            .I(N__30539));
    Span12Mux_s5_h I__6388 (
            .O(N__30544),
            .I(N__30539));
    Odrv12 I__6387 (
            .O(N__30539),
            .I(\ALU.N_762 ));
    InMux I__6386 (
            .O(N__30536),
            .I(N__30532));
    InMux I__6385 (
            .O(N__30535),
            .I(N__30529));
    LocalMux I__6384 (
            .O(N__30532),
            .I(N__30526));
    LocalMux I__6383 (
            .O(N__30529),
            .I(N__30523));
    Span4Mux_h I__6382 (
            .O(N__30526),
            .I(N__30520));
    Span4Mux_h I__6381 (
            .O(N__30523),
            .I(N__30517));
    Span4Mux_v I__6380 (
            .O(N__30520),
            .I(N__30514));
    Span4Mux_v I__6379 (
            .O(N__30517),
            .I(N__30509));
    Span4Mux_h I__6378 (
            .O(N__30514),
            .I(N__30509));
    Odrv4 I__6377 (
            .O(N__30509),
            .I(\ALU.N_714 ));
    CascadeMux I__6376 (
            .O(N__30506),
            .I(\ALU.N_621_1_cascade_ ));
    InMux I__6375 (
            .O(N__30503),
            .I(N__30499));
    InMux I__6374 (
            .O(N__30502),
            .I(N__30496));
    LocalMux I__6373 (
            .O(N__30499),
            .I(N__30492));
    LocalMux I__6372 (
            .O(N__30496),
            .I(N__30489));
    InMux I__6371 (
            .O(N__30495),
            .I(N__30486));
    Odrv4 I__6370 (
            .O(N__30492),
            .I(\ALU.N_589 ));
    Odrv4 I__6369 (
            .O(N__30489),
            .I(\ALU.N_589 ));
    LocalMux I__6368 (
            .O(N__30486),
            .I(\ALU.N_589 ));
    InMux I__6367 (
            .O(N__30479),
            .I(N__30472));
    InMux I__6366 (
            .O(N__30478),
            .I(N__30472));
    InMux I__6365 (
            .O(N__30477),
            .I(N__30466));
    LocalMux I__6364 (
            .O(N__30472),
            .I(N__30463));
    InMux I__6363 (
            .O(N__30471),
            .I(N__30460));
    InMux I__6362 (
            .O(N__30470),
            .I(N__30455));
    InMux I__6361 (
            .O(N__30469),
            .I(N__30455));
    LocalMux I__6360 (
            .O(N__30466),
            .I(N__30452));
    Odrv4 I__6359 (
            .O(N__30463),
            .I(\ALU.N_621_1 ));
    LocalMux I__6358 (
            .O(N__30460),
            .I(\ALU.N_621_1 ));
    LocalMux I__6357 (
            .O(N__30455),
            .I(\ALU.N_621_1 ));
    Odrv4 I__6356 (
            .O(N__30452),
            .I(\ALU.N_621_1 ));
    InMux I__6355 (
            .O(N__30443),
            .I(N__30440));
    LocalMux I__6354 (
            .O(N__30440),
            .I(\ALU.c_RNI4JFV4_0Z0Z_15 ));
    InMux I__6353 (
            .O(N__30437),
            .I(N__30434));
    LocalMux I__6352 (
            .O(N__30434),
            .I(N__30431));
    Odrv12 I__6351 (
            .O(N__30431),
            .I(\ALU.N_274_0 ));
    InMux I__6350 (
            .O(N__30428),
            .I(N__30425));
    LocalMux I__6349 (
            .O(N__30425),
            .I(\ALU.d_RNI36KJ21Z0Z_9 ));
    InMux I__6348 (
            .O(N__30422),
            .I(N__30419));
    LocalMux I__6347 (
            .O(N__30419),
            .I(N__30414));
    InMux I__6346 (
            .O(N__30418),
            .I(N__30411));
    InMux I__6345 (
            .O(N__30417),
            .I(N__30407));
    Span4Mux_s2_v I__6344 (
            .O(N__30414),
            .I(N__30404));
    LocalMux I__6343 (
            .O(N__30411),
            .I(N__30401));
    InMux I__6342 (
            .O(N__30410),
            .I(N__30398));
    LocalMux I__6341 (
            .O(N__30407),
            .I(N__30395));
    Odrv4 I__6340 (
            .O(N__30404),
            .I(\FTDI.TXready ));
    Odrv4 I__6339 (
            .O(N__30401),
            .I(\FTDI.TXready ));
    LocalMux I__6338 (
            .O(N__30398),
            .I(\FTDI.TXready ));
    Odrv12 I__6337 (
            .O(N__30395),
            .I(\FTDI.TXready ));
    InMux I__6336 (
            .O(N__30386),
            .I(N__30381));
    InMux I__6335 (
            .O(N__30385),
            .I(N__30372));
    InMux I__6334 (
            .O(N__30384),
            .I(N__30372));
    LocalMux I__6333 (
            .O(N__30381),
            .I(N__30369));
    InMux I__6332 (
            .O(N__30380),
            .I(N__30366));
    InMux I__6331 (
            .O(N__30379),
            .I(N__30359));
    InMux I__6330 (
            .O(N__30378),
            .I(N__30359));
    InMux I__6329 (
            .O(N__30377),
            .I(N__30359));
    LocalMux I__6328 (
            .O(N__30372),
            .I(N__30356));
    Span4Mux_v I__6327 (
            .O(N__30369),
            .I(N__30349));
    LocalMux I__6326 (
            .O(N__30366),
            .I(N__30349));
    LocalMux I__6325 (
            .O(N__30359),
            .I(N__30349));
    Span4Mux_h I__6324 (
            .O(N__30356),
            .I(N__30346));
    Odrv4 I__6323 (
            .O(N__30349),
            .I(\FTDI.baudAccZ0Z_2 ));
    Odrv4 I__6322 (
            .O(N__30346),
            .I(\FTDI.baudAccZ0Z_2 ));
    InMux I__6321 (
            .O(N__30341),
            .I(N__30338));
    LocalMux I__6320 (
            .O(N__30338),
            .I(N__30333));
    InMux I__6319 (
            .O(N__30337),
            .I(N__30328));
    InMux I__6318 (
            .O(N__30336),
            .I(N__30328));
    Odrv4 I__6317 (
            .O(N__30333),
            .I(TXstartZ0));
    LocalMux I__6316 (
            .O(N__30328),
            .I(TXstartZ0));
    InMux I__6315 (
            .O(N__30323),
            .I(N__30319));
    CascadeMux I__6314 (
            .O(N__30322),
            .I(N__30316));
    LocalMux I__6313 (
            .O(N__30319),
            .I(N__30311));
    InMux I__6312 (
            .O(N__30316),
            .I(N__30306));
    InMux I__6311 (
            .O(N__30315),
            .I(N__30306));
    InMux I__6310 (
            .O(N__30314),
            .I(N__30303));
    Span4Mux_v I__6309 (
            .O(N__30311),
            .I(N__30299));
    LocalMux I__6308 (
            .O(N__30306),
            .I(N__30296));
    LocalMux I__6307 (
            .O(N__30303),
            .I(N__30293));
    CascadeMux I__6306 (
            .O(N__30302),
            .I(N__30286));
    Sp12to4 I__6305 (
            .O(N__30299),
            .I(N__30282));
    Span4Mux_v I__6304 (
            .O(N__30296),
            .I(N__30279));
    Span4Mux_s2_v I__6303 (
            .O(N__30293),
            .I(N__30276));
    InMux I__6302 (
            .O(N__30292),
            .I(N__30269));
    InMux I__6301 (
            .O(N__30291),
            .I(N__30269));
    InMux I__6300 (
            .O(N__30290),
            .I(N__30269));
    InMux I__6299 (
            .O(N__30289),
            .I(N__30264));
    InMux I__6298 (
            .O(N__30286),
            .I(N__30264));
    InMux I__6297 (
            .O(N__30285),
            .I(N__30261));
    Span12Mux_s6_h I__6296 (
            .O(N__30282),
            .I(N__30258));
    Span4Mux_h I__6295 (
            .O(N__30279),
            .I(N__30253));
    Span4Mux_h I__6294 (
            .O(N__30276),
            .I(N__30253));
    LocalMux I__6293 (
            .O(N__30269),
            .I(N__30250));
    LocalMux I__6292 (
            .O(N__30264),
            .I(testStateZ0Z_0));
    LocalMux I__6291 (
            .O(N__30261),
            .I(testStateZ0Z_0));
    Odrv12 I__6290 (
            .O(N__30258),
            .I(testStateZ0Z_0));
    Odrv4 I__6289 (
            .O(N__30253),
            .I(testStateZ0Z_0));
    Odrv12 I__6288 (
            .O(N__30250),
            .I(testStateZ0Z_0));
    InMux I__6287 (
            .O(N__30239),
            .I(N__30235));
    CascadeMux I__6286 (
            .O(N__30238),
            .I(N__30231));
    LocalMux I__6285 (
            .O(N__30235),
            .I(N__30228));
    InMux I__6284 (
            .O(N__30234),
            .I(N__30223));
    InMux I__6283 (
            .O(N__30231),
            .I(N__30223));
    Odrv12 I__6282 (
            .O(N__30228),
            .I(ctrlOut_13));
    LocalMux I__6281 (
            .O(N__30223),
            .I(ctrlOut_13));
    InMux I__6280 (
            .O(N__30218),
            .I(N__30212));
    CascadeMux I__6279 (
            .O(N__30217),
            .I(N__30208));
    CascadeMux I__6278 (
            .O(N__30216),
            .I(N__30202));
    InMux I__6277 (
            .O(N__30215),
            .I(N__30197));
    LocalMux I__6276 (
            .O(N__30212),
            .I(N__30189));
    InMux I__6275 (
            .O(N__30211),
            .I(N__30186));
    InMux I__6274 (
            .O(N__30208),
            .I(N__30181));
    InMux I__6273 (
            .O(N__30207),
            .I(N__30181));
    InMux I__6272 (
            .O(N__30206),
            .I(N__30176));
    InMux I__6271 (
            .O(N__30205),
            .I(N__30176));
    InMux I__6270 (
            .O(N__30202),
            .I(N__30173));
    InMux I__6269 (
            .O(N__30201),
            .I(N__30167));
    InMux I__6268 (
            .O(N__30200),
            .I(N__30164));
    LocalMux I__6267 (
            .O(N__30197),
            .I(N__30161));
    InMux I__6266 (
            .O(N__30196),
            .I(N__30158));
    InMux I__6265 (
            .O(N__30195),
            .I(N__30153));
    InMux I__6264 (
            .O(N__30194),
            .I(N__30153));
    InMux I__6263 (
            .O(N__30193),
            .I(N__30148));
    InMux I__6262 (
            .O(N__30192),
            .I(N__30148));
    Span4Mux_h I__6261 (
            .O(N__30189),
            .I(N__30143));
    LocalMux I__6260 (
            .O(N__30186),
            .I(N__30143));
    LocalMux I__6259 (
            .O(N__30181),
            .I(N__30140));
    LocalMux I__6258 (
            .O(N__30176),
            .I(N__30137));
    LocalMux I__6257 (
            .O(N__30173),
            .I(N__30132));
    InMux I__6256 (
            .O(N__30172),
            .I(N__30122));
    InMux I__6255 (
            .O(N__30171),
            .I(N__30122));
    InMux I__6254 (
            .O(N__30170),
            .I(N__30122));
    LocalMux I__6253 (
            .O(N__30167),
            .I(N__30117));
    LocalMux I__6252 (
            .O(N__30164),
            .I(N__30117));
    Span4Mux_v I__6251 (
            .O(N__30161),
            .I(N__30112));
    LocalMux I__6250 (
            .O(N__30158),
            .I(N__30112));
    LocalMux I__6249 (
            .O(N__30153),
            .I(N__30109));
    LocalMux I__6248 (
            .O(N__30148),
            .I(N__30106));
    Span4Mux_h I__6247 (
            .O(N__30143),
            .I(N__30103));
    Span4Mux_v I__6246 (
            .O(N__30140),
            .I(N__30098));
    Span4Mux_s1_h I__6245 (
            .O(N__30137),
            .I(N__30098));
    InMux I__6244 (
            .O(N__30136),
            .I(N__30093));
    InMux I__6243 (
            .O(N__30135),
            .I(N__30093));
    Span4Mux_v I__6242 (
            .O(N__30132),
            .I(N__30090));
    InMux I__6241 (
            .O(N__30131),
            .I(N__30083));
    InMux I__6240 (
            .O(N__30130),
            .I(N__30083));
    InMux I__6239 (
            .O(N__30129),
            .I(N__30083));
    LocalMux I__6238 (
            .O(N__30122),
            .I(N__30074));
    Span4Mux_h I__6237 (
            .O(N__30117),
            .I(N__30074));
    Span4Mux_v I__6236 (
            .O(N__30112),
            .I(N__30074));
    Span4Mux_h I__6235 (
            .O(N__30109),
            .I(N__30074));
    Odrv4 I__6234 (
            .O(N__30106),
            .I(busState_2));
    Odrv4 I__6233 (
            .O(N__30103),
            .I(busState_2));
    Odrv4 I__6232 (
            .O(N__30098),
            .I(busState_2));
    LocalMux I__6231 (
            .O(N__30093),
            .I(busState_2));
    Odrv4 I__6230 (
            .O(N__30090),
            .I(busState_2));
    LocalMux I__6229 (
            .O(N__30083),
            .I(busState_2));
    Odrv4 I__6228 (
            .O(N__30074),
            .I(busState_2));
    CascadeMux I__6227 (
            .O(N__30059),
            .I(N__30051));
    CascadeMux I__6226 (
            .O(N__30058),
            .I(N__30046));
    CascadeMux I__6225 (
            .O(N__30057),
            .I(N__30042));
    CascadeMux I__6224 (
            .O(N__30056),
            .I(N__30039));
    CascadeMux I__6223 (
            .O(N__30055),
            .I(N__30036));
    CascadeMux I__6222 (
            .O(N__30054),
            .I(N__30033));
    InMux I__6221 (
            .O(N__30051),
            .I(N__30027));
    CascadeMux I__6220 (
            .O(N__30050),
            .I(N__30018));
    InMux I__6219 (
            .O(N__30049),
            .I(N__30015));
    InMux I__6218 (
            .O(N__30046),
            .I(N__30007));
    InMux I__6217 (
            .O(N__30045),
            .I(N__30007));
    InMux I__6216 (
            .O(N__30042),
            .I(N__30002));
    InMux I__6215 (
            .O(N__30039),
            .I(N__30002));
    InMux I__6214 (
            .O(N__30036),
            .I(N__29995));
    InMux I__6213 (
            .O(N__30033),
            .I(N__29995));
    InMux I__6212 (
            .O(N__30032),
            .I(N__29995));
    CascadeMux I__6211 (
            .O(N__30031),
            .I(N__29990));
    CascadeMux I__6210 (
            .O(N__30030),
            .I(N__29987));
    LocalMux I__6209 (
            .O(N__30027),
            .I(N__29984));
    InMux I__6208 (
            .O(N__30026),
            .I(N__29981));
    CascadeMux I__6207 (
            .O(N__30025),
            .I(N__29977));
    CascadeMux I__6206 (
            .O(N__30024),
            .I(N__29974));
    CascadeMux I__6205 (
            .O(N__30023),
            .I(N__29971));
    CascadeMux I__6204 (
            .O(N__30022),
            .I(N__29968));
    InMux I__6203 (
            .O(N__30021),
            .I(N__29963));
    InMux I__6202 (
            .O(N__30018),
            .I(N__29960));
    LocalMux I__6201 (
            .O(N__30015),
            .I(N__29957));
    CascadeMux I__6200 (
            .O(N__30014),
            .I(N__29951));
    CascadeMux I__6199 (
            .O(N__30013),
            .I(N__29948));
    CascadeMux I__6198 (
            .O(N__30012),
            .I(N__29945));
    LocalMux I__6197 (
            .O(N__30007),
            .I(N__29942));
    LocalMux I__6196 (
            .O(N__30002),
            .I(N__29937));
    LocalMux I__6195 (
            .O(N__29995),
            .I(N__29937));
    CascadeMux I__6194 (
            .O(N__29994),
            .I(N__29934));
    CascadeMux I__6193 (
            .O(N__29993),
            .I(N__29931));
    InMux I__6192 (
            .O(N__29990),
            .I(N__29926));
    InMux I__6191 (
            .O(N__29987),
            .I(N__29926));
    Span4Mux_v I__6190 (
            .O(N__29984),
            .I(N__29921));
    LocalMux I__6189 (
            .O(N__29981),
            .I(N__29921));
    InMux I__6188 (
            .O(N__29980),
            .I(N__29918));
    InMux I__6187 (
            .O(N__29977),
            .I(N__29915));
    InMux I__6186 (
            .O(N__29974),
            .I(N__29911));
    InMux I__6185 (
            .O(N__29971),
            .I(N__29908));
    InMux I__6184 (
            .O(N__29968),
            .I(N__29905));
    CascadeMux I__6183 (
            .O(N__29967),
            .I(N__29902));
    InMux I__6182 (
            .O(N__29966),
            .I(N__29899));
    LocalMux I__6181 (
            .O(N__29963),
            .I(N__29891));
    LocalMux I__6180 (
            .O(N__29960),
            .I(N__29891));
    Span4Mux_h I__6179 (
            .O(N__29957),
            .I(N__29891));
    CascadeMux I__6178 (
            .O(N__29956),
            .I(N__29888));
    InMux I__6177 (
            .O(N__29955),
            .I(N__29883));
    InMux I__6176 (
            .O(N__29954),
            .I(N__29883));
    InMux I__6175 (
            .O(N__29951),
            .I(N__29880));
    InMux I__6174 (
            .O(N__29948),
            .I(N__29875));
    InMux I__6173 (
            .O(N__29945),
            .I(N__29875));
    Span4Mux_h I__6172 (
            .O(N__29942),
            .I(N__29870));
    Span4Mux_v I__6171 (
            .O(N__29937),
            .I(N__29870));
    InMux I__6170 (
            .O(N__29934),
            .I(N__29865));
    InMux I__6169 (
            .O(N__29931),
            .I(N__29865));
    LocalMux I__6168 (
            .O(N__29926),
            .I(N__29860));
    Span4Mux_v I__6167 (
            .O(N__29921),
            .I(N__29860));
    LocalMux I__6166 (
            .O(N__29918),
            .I(N__29857));
    LocalMux I__6165 (
            .O(N__29915),
            .I(N__29854));
    CascadeMux I__6164 (
            .O(N__29914),
            .I(N__29851));
    LocalMux I__6163 (
            .O(N__29911),
            .I(N__29844));
    LocalMux I__6162 (
            .O(N__29908),
            .I(N__29844));
    LocalMux I__6161 (
            .O(N__29905),
            .I(N__29844));
    InMux I__6160 (
            .O(N__29902),
            .I(N__29841));
    LocalMux I__6159 (
            .O(N__29899),
            .I(N__29838));
    CascadeMux I__6158 (
            .O(N__29898),
            .I(N__29833));
    Span4Mux_h I__6157 (
            .O(N__29891),
            .I(N__29830));
    InMux I__6156 (
            .O(N__29888),
            .I(N__29827));
    LocalMux I__6155 (
            .O(N__29883),
            .I(N__29818));
    LocalMux I__6154 (
            .O(N__29880),
            .I(N__29818));
    LocalMux I__6153 (
            .O(N__29875),
            .I(N__29818));
    Span4Mux_v I__6152 (
            .O(N__29870),
            .I(N__29818));
    LocalMux I__6151 (
            .O(N__29865),
            .I(N__29815));
    Span4Mux_h I__6150 (
            .O(N__29860),
            .I(N__29810));
    Span4Mux_v I__6149 (
            .O(N__29857),
            .I(N__29810));
    Span4Mux_h I__6148 (
            .O(N__29854),
            .I(N__29807));
    InMux I__6147 (
            .O(N__29851),
            .I(N__29804));
    Span4Mux_v I__6146 (
            .O(N__29844),
            .I(N__29801));
    LocalMux I__6145 (
            .O(N__29841),
            .I(N__29798));
    Span12Mux_v I__6144 (
            .O(N__29838),
            .I(N__29795));
    InMux I__6143 (
            .O(N__29837),
            .I(N__29788));
    InMux I__6142 (
            .O(N__29836),
            .I(N__29788));
    InMux I__6141 (
            .O(N__29833),
            .I(N__29788));
    Span4Mux_v I__6140 (
            .O(N__29830),
            .I(N__29785));
    LocalMux I__6139 (
            .O(N__29827),
            .I(N__29780));
    Span4Mux_h I__6138 (
            .O(N__29818),
            .I(N__29780));
    Span4Mux_v I__6137 (
            .O(N__29815),
            .I(N__29773));
    Span4Mux_v I__6136 (
            .O(N__29810),
            .I(N__29773));
    Span4Mux_h I__6135 (
            .O(N__29807),
            .I(N__29773));
    LocalMux I__6134 (
            .O(N__29804),
            .I(aluReadBus_rep2));
    Odrv4 I__6133 (
            .O(N__29801),
            .I(aluReadBus_rep2));
    Odrv12 I__6132 (
            .O(N__29798),
            .I(aluReadBus_rep2));
    Odrv12 I__6131 (
            .O(N__29795),
            .I(aluReadBus_rep2));
    LocalMux I__6130 (
            .O(N__29788),
            .I(aluReadBus_rep2));
    Odrv4 I__6129 (
            .O(N__29785),
            .I(aluReadBus_rep2));
    Odrv4 I__6128 (
            .O(N__29780),
            .I(aluReadBus_rep2));
    Odrv4 I__6127 (
            .O(N__29773),
            .I(aluReadBus_rep2));
    CascadeMux I__6126 (
            .O(N__29756),
            .I(N__29750));
    CascadeMux I__6125 (
            .O(N__29755),
            .I(N__29747));
    InMux I__6124 (
            .O(N__29754),
            .I(N__29742));
    InMux I__6123 (
            .O(N__29753),
            .I(N__29736));
    InMux I__6122 (
            .O(N__29750),
            .I(N__29730));
    InMux I__6121 (
            .O(N__29747),
            .I(N__29730));
    InMux I__6120 (
            .O(N__29746),
            .I(N__29723));
    InMux I__6119 (
            .O(N__29745),
            .I(N__29723));
    LocalMux I__6118 (
            .O(N__29742),
            .I(N__29720));
    InMux I__6117 (
            .O(N__29741),
            .I(N__29717));
    InMux I__6116 (
            .O(N__29740),
            .I(N__29714));
    InMux I__6115 (
            .O(N__29739),
            .I(N__29711));
    LocalMux I__6114 (
            .O(N__29736),
            .I(N__29708));
    InMux I__6113 (
            .O(N__29735),
            .I(N__29705));
    LocalMux I__6112 (
            .O(N__29730),
            .I(N__29698));
    InMux I__6111 (
            .O(N__29729),
            .I(N__29693));
    InMux I__6110 (
            .O(N__29728),
            .I(N__29693));
    LocalMux I__6109 (
            .O(N__29723),
            .I(N__29688));
    Span4Mux_h I__6108 (
            .O(N__29720),
            .I(N__29683));
    LocalMux I__6107 (
            .O(N__29717),
            .I(N__29683));
    LocalMux I__6106 (
            .O(N__29714),
            .I(N__29673));
    LocalMux I__6105 (
            .O(N__29711),
            .I(N__29673));
    Span4Mux_v I__6104 (
            .O(N__29708),
            .I(N__29668));
    LocalMux I__6103 (
            .O(N__29705),
            .I(N__29668));
    InMux I__6102 (
            .O(N__29704),
            .I(N__29659));
    InMux I__6101 (
            .O(N__29703),
            .I(N__29659));
    InMux I__6100 (
            .O(N__29702),
            .I(N__29659));
    InMux I__6099 (
            .O(N__29701),
            .I(N__29659));
    Span4Mux_v I__6098 (
            .O(N__29698),
            .I(N__29654));
    LocalMux I__6097 (
            .O(N__29693),
            .I(N__29654));
    InMux I__6096 (
            .O(N__29692),
            .I(N__29649));
    InMux I__6095 (
            .O(N__29691),
            .I(N__29649));
    Span4Mux_h I__6094 (
            .O(N__29688),
            .I(N__29644));
    Span4Mux_h I__6093 (
            .O(N__29683),
            .I(N__29644));
    InMux I__6092 (
            .O(N__29682),
            .I(N__29639));
    InMux I__6091 (
            .O(N__29681),
            .I(N__29639));
    InMux I__6090 (
            .O(N__29680),
            .I(N__29632));
    InMux I__6089 (
            .O(N__29679),
            .I(N__29632));
    InMux I__6088 (
            .O(N__29678),
            .I(N__29632));
    Span4Mux_h I__6087 (
            .O(N__29673),
            .I(N__29623));
    Span4Mux_v I__6086 (
            .O(N__29668),
            .I(N__29623));
    LocalMux I__6085 (
            .O(N__29659),
            .I(N__29623));
    Span4Mux_h I__6084 (
            .O(N__29654),
            .I(N__29623));
    LocalMux I__6083 (
            .O(N__29649),
            .I(busState_0));
    Odrv4 I__6082 (
            .O(N__29644),
            .I(busState_0));
    LocalMux I__6081 (
            .O(N__29639),
            .I(busState_0));
    LocalMux I__6080 (
            .O(N__29632),
            .I(busState_0));
    Odrv4 I__6079 (
            .O(N__29623),
            .I(busState_0));
    InMux I__6078 (
            .O(N__29612),
            .I(N__29609));
    LocalMux I__6077 (
            .O(N__29609),
            .I(N__29606));
    Span4Mux_v I__6076 (
            .O(N__29606),
            .I(N__29603));
    Odrv4 I__6075 (
            .O(N__29603),
            .I(\ALU.N_9_1 ));
    CascadeMux I__6074 (
            .O(N__29600),
            .I(\FTDI.N_217_0_cascade_ ));
    InMux I__6073 (
            .O(N__29597),
            .I(N__29594));
    LocalMux I__6072 (
            .O(N__29594),
            .I(\FTDI.N_216_0 ));
    CascadeMux I__6071 (
            .O(N__29591),
            .I(\FTDI.TXready_cascade_ ));
    InMux I__6070 (
            .O(N__29588),
            .I(N__29583));
    InMux I__6069 (
            .O(N__29587),
            .I(N__29580));
    InMux I__6068 (
            .O(N__29586),
            .I(N__29577));
    LocalMux I__6067 (
            .O(N__29583),
            .I(\FTDI.baudAccZ0Z_0 ));
    LocalMux I__6066 (
            .O(N__29580),
            .I(\FTDI.baudAccZ0Z_0 ));
    LocalMux I__6065 (
            .O(N__29577),
            .I(\FTDI.baudAccZ0Z_0 ));
    InMux I__6064 (
            .O(N__29570),
            .I(N__29567));
    LocalMux I__6063 (
            .O(N__29567),
            .I(N__29564));
    Span4Mux_h I__6062 (
            .O(N__29564),
            .I(N__29560));
    InMux I__6061 (
            .O(N__29563),
            .I(N__29557));
    Odrv4 I__6060 (
            .O(N__29560),
            .I(\FTDI.baudAccZ0Z_1 ));
    LocalMux I__6059 (
            .O(N__29557),
            .I(\FTDI.baudAccZ0Z_1 ));
    InMux I__6058 (
            .O(N__29552),
            .I(N__29549));
    LocalMux I__6057 (
            .O(N__29549),
            .I(N__29546));
    Span4Mux_h I__6056 (
            .O(N__29546),
            .I(N__29543));
    Span4Mux_h I__6055 (
            .O(N__29543),
            .I(N__29540));
    Span4Mux_h I__6054 (
            .O(N__29540),
            .I(N__29537));
    Odrv4 I__6053 (
            .O(N__29537),
            .I(\ALU.N_290_0 ));
    InMux I__6052 (
            .O(N__29534),
            .I(N__29531));
    LocalMux I__6051 (
            .O(N__29531),
            .I(\ALU.rshift_5 ));
    InMux I__6050 (
            .O(N__29528),
            .I(N__29525));
    LocalMux I__6049 (
            .O(N__29525),
            .I(\ALU.a_15_m3_5 ));
    InMux I__6048 (
            .O(N__29522),
            .I(N__29514));
    InMux I__6047 (
            .O(N__29521),
            .I(N__29507));
    InMux I__6046 (
            .O(N__29520),
            .I(N__29507));
    InMux I__6045 (
            .O(N__29519),
            .I(N__29507));
    InMux I__6044 (
            .O(N__29518),
            .I(N__29502));
    InMux I__6043 (
            .O(N__29517),
            .I(N__29502));
    LocalMux I__6042 (
            .O(N__29514),
            .I(\FTDI.TXstateZ1Z_0 ));
    LocalMux I__6041 (
            .O(N__29507),
            .I(\FTDI.TXstateZ1Z_0 ));
    LocalMux I__6040 (
            .O(N__29502),
            .I(\FTDI.TXstateZ1Z_0 ));
    InMux I__6039 (
            .O(N__29495),
            .I(N__29483));
    InMux I__6038 (
            .O(N__29494),
            .I(N__29483));
    InMux I__6037 (
            .O(N__29493),
            .I(N__29483));
    InMux I__6036 (
            .O(N__29492),
            .I(N__29480));
    InMux I__6035 (
            .O(N__29491),
            .I(N__29475));
    InMux I__6034 (
            .O(N__29490),
            .I(N__29475));
    LocalMux I__6033 (
            .O(N__29483),
            .I(\FTDI.TXstateZ1Z_1 ));
    LocalMux I__6032 (
            .O(N__29480),
            .I(\FTDI.TXstateZ1Z_1 ));
    LocalMux I__6031 (
            .O(N__29475),
            .I(\FTDI.TXstateZ1Z_1 ));
    InMux I__6030 (
            .O(N__29468),
            .I(N__29464));
    InMux I__6029 (
            .O(N__29467),
            .I(N__29461));
    LocalMux I__6028 (
            .O(N__29464),
            .I(\FTDI.N_170_0 ));
    LocalMux I__6027 (
            .O(N__29461),
            .I(\FTDI.N_170_0 ));
    CascadeMux I__6026 (
            .O(N__29456),
            .I(\FTDI.TXstate_e_1_3_cascade_ ));
    InMux I__6025 (
            .O(N__29453),
            .I(N__29450));
    LocalMux I__6024 (
            .O(N__29450),
            .I(N__29447));
    Span4Mux_h I__6023 (
            .O(N__29447),
            .I(N__29444));
    Span4Mux_h I__6022 (
            .O(N__29444),
            .I(N__29441));
    Odrv4 I__6021 (
            .O(N__29441),
            .I(\ALU.N_11_0 ));
    CascadeMux I__6020 (
            .O(N__29438),
            .I(N__29430));
    InMux I__6019 (
            .O(N__29437),
            .I(N__29427));
    InMux I__6018 (
            .O(N__29436),
            .I(N__29423));
    InMux I__6017 (
            .O(N__29435),
            .I(N__29420));
    CascadeMux I__6016 (
            .O(N__29434),
            .I(N__29417));
    CascadeMux I__6015 (
            .O(N__29433),
            .I(N__29414));
    InMux I__6014 (
            .O(N__29430),
            .I(N__29409));
    LocalMux I__6013 (
            .O(N__29427),
            .I(N__29406));
    InMux I__6012 (
            .O(N__29426),
            .I(N__29399));
    LocalMux I__6011 (
            .O(N__29423),
            .I(N__29394));
    LocalMux I__6010 (
            .O(N__29420),
            .I(N__29394));
    InMux I__6009 (
            .O(N__29417),
            .I(N__29387));
    InMux I__6008 (
            .O(N__29414),
            .I(N__29387));
    InMux I__6007 (
            .O(N__29413),
            .I(N__29387));
    InMux I__6006 (
            .O(N__29412),
            .I(N__29384));
    LocalMux I__6005 (
            .O(N__29409),
            .I(N__29381));
    Span4Mux_h I__6004 (
            .O(N__29406),
            .I(N__29374));
    InMux I__6003 (
            .O(N__29405),
            .I(N__29371));
    InMux I__6002 (
            .O(N__29404),
            .I(N__29368));
    InMux I__6001 (
            .O(N__29403),
            .I(N__29362));
    InMux I__6000 (
            .O(N__29402),
            .I(N__29362));
    LocalMux I__5999 (
            .O(N__29399),
            .I(N__29355));
    Span4Mux_v I__5998 (
            .O(N__29394),
            .I(N__29355));
    LocalMux I__5997 (
            .O(N__29387),
            .I(N__29355));
    LocalMux I__5996 (
            .O(N__29384),
            .I(N__29352));
    Span4Mux_h I__5995 (
            .O(N__29381),
            .I(N__29349));
    InMux I__5994 (
            .O(N__29380),
            .I(N__29342));
    InMux I__5993 (
            .O(N__29379),
            .I(N__29342));
    InMux I__5992 (
            .O(N__29378),
            .I(N__29342));
    InMux I__5991 (
            .O(N__29377),
            .I(N__29339));
    Span4Mux_h I__5990 (
            .O(N__29374),
            .I(N__29334));
    LocalMux I__5989 (
            .O(N__29371),
            .I(N__29334));
    LocalMux I__5988 (
            .O(N__29368),
            .I(N__29331));
    InMux I__5987 (
            .O(N__29367),
            .I(N__29328));
    LocalMux I__5986 (
            .O(N__29362),
            .I(N__29325));
    Span4Mux_h I__5985 (
            .O(N__29355),
            .I(N__29316));
    Span4Mux_h I__5984 (
            .O(N__29352),
            .I(N__29316));
    Span4Mux_v I__5983 (
            .O(N__29349),
            .I(N__29316));
    LocalMux I__5982 (
            .O(N__29342),
            .I(N__29316));
    LocalMux I__5981 (
            .O(N__29339),
            .I(N__29311));
    Span4Mux_h I__5980 (
            .O(N__29334),
            .I(N__29311));
    Span4Mux_v I__5979 (
            .O(N__29331),
            .I(N__29306));
    LocalMux I__5978 (
            .O(N__29328),
            .I(N__29299));
    Span4Mux_v I__5977 (
            .O(N__29325),
            .I(N__29299));
    Span4Mux_v I__5976 (
            .O(N__29316),
            .I(N__29299));
    Sp12to4 I__5975 (
            .O(N__29311),
            .I(N__29296));
    InMux I__5974 (
            .O(N__29310),
            .I(N__29293));
    InMux I__5973 (
            .O(N__29309),
            .I(N__29289));
    Span4Mux_h I__5972 (
            .O(N__29306),
            .I(N__29284));
    Span4Mux_v I__5971 (
            .O(N__29299),
            .I(N__29284));
    Span12Mux_s6_v I__5970 (
            .O(N__29296),
            .I(N__29279));
    LocalMux I__5969 (
            .O(N__29293),
            .I(N__29279));
    InMux I__5968 (
            .O(N__29292),
            .I(N__29276));
    LocalMux I__5967 (
            .O(N__29289),
            .I(\ALU.N_5_0 ));
    Odrv4 I__5966 (
            .O(N__29284),
            .I(\ALU.N_5_0 ));
    Odrv12 I__5965 (
            .O(N__29279),
            .I(\ALU.N_5_0 ));
    LocalMux I__5964 (
            .O(N__29276),
            .I(\ALU.N_5_0 ));
    CascadeMux I__5963 (
            .O(N__29267),
            .I(N__29263));
    CascadeMux I__5962 (
            .O(N__29266),
            .I(N__29258));
    InMux I__5961 (
            .O(N__29263),
            .I(N__29251));
    InMux I__5960 (
            .O(N__29262),
            .I(N__29251));
    InMux I__5959 (
            .O(N__29261),
            .I(N__29251));
    InMux I__5958 (
            .O(N__29258),
            .I(N__29246));
    LocalMux I__5957 (
            .O(N__29251),
            .I(N__29243));
    InMux I__5956 (
            .O(N__29250),
            .I(N__29238));
    InMux I__5955 (
            .O(N__29249),
            .I(N__29238));
    LocalMux I__5954 (
            .O(N__29246),
            .I(N__29235));
    Span4Mux_v I__5953 (
            .O(N__29243),
            .I(N__29230));
    LocalMux I__5952 (
            .O(N__29238),
            .I(N__29230));
    Span4Mux_h I__5951 (
            .O(N__29235),
            .I(N__29227));
    Span4Mux_h I__5950 (
            .O(N__29230),
            .I(N__29224));
    Odrv4 I__5949 (
            .O(N__29227),
            .I(\FTDI.gapZ0Z_2 ));
    Odrv4 I__5948 (
            .O(N__29224),
            .I(\FTDI.gapZ0Z_2 ));
    CascadeMux I__5947 (
            .O(N__29219),
            .I(N__29216));
    InMux I__5946 (
            .O(N__29216),
            .I(N__29210));
    InMux I__5945 (
            .O(N__29215),
            .I(N__29210));
    LocalMux I__5944 (
            .O(N__29210),
            .I(N__29207));
    Span4Mux_s1_v I__5943 (
            .O(N__29207),
            .I(N__29203));
    InMux I__5942 (
            .O(N__29206),
            .I(N__29200));
    Odrv4 I__5941 (
            .O(N__29203),
            .I(\FTDI.gapZ0Z_0 ));
    LocalMux I__5940 (
            .O(N__29200),
            .I(\FTDI.gapZ0Z_0 ));
    InMux I__5939 (
            .O(N__29195),
            .I(N__29190));
    InMux I__5938 (
            .O(N__29194),
            .I(N__29185));
    InMux I__5937 (
            .O(N__29193),
            .I(N__29185));
    LocalMux I__5936 (
            .O(N__29190),
            .I(N__29182));
    LocalMux I__5935 (
            .O(N__29185),
            .I(N__29179));
    IoSpan4Mux I__5934 (
            .O(N__29182),
            .I(N__29176));
    Span4Mux_h I__5933 (
            .O(N__29179),
            .I(N__29171));
    Span4Mux_s0_v I__5932 (
            .O(N__29176),
            .I(N__29171));
    Odrv4 I__5931 (
            .O(N__29171),
            .I(\FTDI.gap8 ));
    InMux I__5930 (
            .O(N__29168),
            .I(N__29162));
    InMux I__5929 (
            .O(N__29167),
            .I(N__29162));
    LocalMux I__5928 (
            .O(N__29162),
            .I(\FTDI.gapZ0Z_1 ));
    InMux I__5927 (
            .O(N__29159),
            .I(N__29156));
    LocalMux I__5926 (
            .O(N__29156),
            .I(\FTDI.TXstate_e_1_0 ));
    CascadeMux I__5925 (
            .O(N__29153),
            .I(\FTDI.N_169_0_cascade_ ));
    CascadeMux I__5924 (
            .O(N__29150),
            .I(N__29147));
    InMux I__5923 (
            .O(N__29147),
            .I(N__29144));
    LocalMux I__5922 (
            .O(N__29144),
            .I(\FTDI.N_169_0 ));
    CascadeMux I__5921 (
            .O(N__29141),
            .I(\FTDI.TXstate_cnst_0_0_2_cascade_ ));
    InMux I__5920 (
            .O(N__29138),
            .I(N__29135));
    LocalMux I__5919 (
            .O(N__29135),
            .I(N__29131));
    InMux I__5918 (
            .O(N__29134),
            .I(N__29128));
    Span4Mux_h I__5917 (
            .O(N__29131),
            .I(N__29125));
    LocalMux I__5916 (
            .O(N__29128),
            .I(N__29122));
    Odrv4 I__5915 (
            .O(N__29125),
            .I(\ALU.cZ0Z_0 ));
    Odrv4 I__5914 (
            .O(N__29122),
            .I(\ALU.cZ0Z_0 ));
    InMux I__5913 (
            .O(N__29117),
            .I(N__29114));
    LocalMux I__5912 (
            .O(N__29114),
            .I(N__29111));
    Span4Mux_v I__5911 (
            .O(N__29111),
            .I(N__29107));
    InMux I__5910 (
            .O(N__29110),
            .I(N__29104));
    Span4Mux_h I__5909 (
            .O(N__29107),
            .I(N__29101));
    LocalMux I__5908 (
            .O(N__29104),
            .I(\ALU.cZ0Z_1 ));
    Odrv4 I__5907 (
            .O(N__29101),
            .I(\ALU.cZ0Z_1 ));
    CascadeMux I__5906 (
            .O(N__29096),
            .I(N__29093));
    InMux I__5905 (
            .O(N__29093),
            .I(N__29090));
    LocalMux I__5904 (
            .O(N__29090),
            .I(N__29086));
    InMux I__5903 (
            .O(N__29089),
            .I(N__29083));
    Span4Mux_v I__5902 (
            .O(N__29086),
            .I(N__29080));
    LocalMux I__5901 (
            .O(N__29083),
            .I(N__29077));
    Odrv4 I__5900 (
            .O(N__29080),
            .I(\ALU.cZ0Z_2 ));
    Odrv4 I__5899 (
            .O(N__29077),
            .I(\ALU.cZ0Z_2 ));
    InMux I__5898 (
            .O(N__29072),
            .I(N__29068));
    InMux I__5897 (
            .O(N__29071),
            .I(N__29065));
    LocalMux I__5896 (
            .O(N__29068),
            .I(N__29062));
    LocalMux I__5895 (
            .O(N__29065),
            .I(N__29059));
    Span4Mux_h I__5894 (
            .O(N__29062),
            .I(N__29056));
    Odrv4 I__5893 (
            .O(N__29059),
            .I(\ALU.cZ0Z_3 ));
    Odrv4 I__5892 (
            .O(N__29056),
            .I(\ALU.cZ0Z_3 ));
    InMux I__5891 (
            .O(N__29051),
            .I(N__29048));
    LocalMux I__5890 (
            .O(N__29048),
            .I(N__29044));
    InMux I__5889 (
            .O(N__29047),
            .I(N__29041));
    Span4Mux_v I__5888 (
            .O(N__29044),
            .I(N__29036));
    LocalMux I__5887 (
            .O(N__29041),
            .I(N__29036));
    Span4Mux_h I__5886 (
            .O(N__29036),
            .I(N__29033));
    Odrv4 I__5885 (
            .O(N__29033),
            .I(\ALU.cZ0Z_4 ));
    InMux I__5884 (
            .O(N__29030),
            .I(N__29027));
    LocalMux I__5883 (
            .O(N__29027),
            .I(N__29023));
    InMux I__5882 (
            .O(N__29026),
            .I(N__29020));
    Odrv12 I__5881 (
            .O(N__29023),
            .I(\ALU.cZ0Z_5 ));
    LocalMux I__5880 (
            .O(N__29020),
            .I(\ALU.cZ0Z_5 ));
    InMux I__5879 (
            .O(N__29015),
            .I(N__29012));
    LocalMux I__5878 (
            .O(N__29012),
            .I(N__29008));
    InMux I__5877 (
            .O(N__29011),
            .I(N__29005));
    Span4Mux_h I__5876 (
            .O(N__29008),
            .I(N__29002));
    LocalMux I__5875 (
            .O(N__29005),
            .I(\ALU.cZ0Z_6 ));
    Odrv4 I__5874 (
            .O(N__29002),
            .I(\ALU.cZ0Z_6 ));
    InMux I__5873 (
            .O(N__28997),
            .I(N__28994));
    LocalMux I__5872 (
            .O(N__28994),
            .I(N__28991));
    Span4Mux_h I__5871 (
            .O(N__28991),
            .I(N__28987));
    InMux I__5870 (
            .O(N__28990),
            .I(N__28984));
    Span4Mux_v I__5869 (
            .O(N__28987),
            .I(N__28979));
    LocalMux I__5868 (
            .O(N__28984),
            .I(N__28979));
    Odrv4 I__5867 (
            .O(N__28979),
            .I(\ALU.dZ0Z_4 ));
    InMux I__5866 (
            .O(N__28976),
            .I(N__28972));
    InMux I__5865 (
            .O(N__28975),
            .I(N__28969));
    LocalMux I__5864 (
            .O(N__28972),
            .I(N__28966));
    LocalMux I__5863 (
            .O(N__28969),
            .I(N__28963));
    Span4Mux_h I__5862 (
            .O(N__28966),
            .I(N__28960));
    Span4Mux_h I__5861 (
            .O(N__28963),
            .I(N__28957));
    Odrv4 I__5860 (
            .O(N__28960),
            .I(\ALU.gZ0Z_6 ));
    Odrv4 I__5859 (
            .O(N__28957),
            .I(\ALU.gZ0Z_6 ));
    InMux I__5858 (
            .O(N__28952),
            .I(N__28949));
    LocalMux I__5857 (
            .O(N__28949),
            .I(N__28945));
    InMux I__5856 (
            .O(N__28948),
            .I(N__28942));
    Odrv12 I__5855 (
            .O(N__28945),
            .I(\ALU.eZ0Z_0 ));
    LocalMux I__5854 (
            .O(N__28942),
            .I(\ALU.eZ0Z_0 ));
    InMux I__5853 (
            .O(N__28937),
            .I(N__28934));
    LocalMux I__5852 (
            .O(N__28934),
            .I(N__28930));
    InMux I__5851 (
            .O(N__28933),
            .I(N__28927));
    Span4Mux_v I__5850 (
            .O(N__28930),
            .I(N__28923));
    LocalMux I__5849 (
            .O(N__28927),
            .I(N__28920));
    InMux I__5848 (
            .O(N__28926),
            .I(N__28917));
    Span4Mux_v I__5847 (
            .O(N__28923),
            .I(N__28914));
    Span4Mux_v I__5846 (
            .O(N__28920),
            .I(N__28909));
    LocalMux I__5845 (
            .O(N__28917),
            .I(N__28909));
    Odrv4 I__5844 (
            .O(N__28914),
            .I(a_0));
    Odrv4 I__5843 (
            .O(N__28909),
            .I(a_0));
    CascadeMux I__5842 (
            .O(N__28904),
            .I(N__28901));
    InMux I__5841 (
            .O(N__28901),
            .I(N__28898));
    LocalMux I__5840 (
            .O(N__28898),
            .I(N__28895));
    Odrv12 I__5839 (
            .O(N__28895),
            .I(\ALU.e_RNINIVJZ0Z_0 ));
    InMux I__5838 (
            .O(N__28892),
            .I(N__28889));
    LocalMux I__5837 (
            .O(N__28889),
            .I(\ALU.g_RNIM8LLZ0Z_5 ));
    CascadeMux I__5836 (
            .O(N__28886),
            .I(\ALU.e_RNI1TVJZ0Z_5_cascade_ ));
    InMux I__5835 (
            .O(N__28883),
            .I(N__28880));
    LocalMux I__5834 (
            .O(N__28880),
            .I(N__28877));
    Span4Mux_v I__5833 (
            .O(N__28877),
            .I(N__28874));
    Span4Mux_h I__5832 (
            .O(N__28874),
            .I(N__28871));
    Odrv4 I__5831 (
            .O(N__28871),
            .I(\ALU.operand2_7_ns_1_5 ));
    InMux I__5830 (
            .O(N__28868),
            .I(N__28865));
    LocalMux I__5829 (
            .O(N__28865),
            .I(N__28862));
    Span4Mux_h I__5828 (
            .O(N__28862),
            .I(N__28858));
    InMux I__5827 (
            .O(N__28861),
            .I(N__28855));
    Odrv4 I__5826 (
            .O(N__28858),
            .I(\ALU.eZ0Z_5 ));
    LocalMux I__5825 (
            .O(N__28855),
            .I(\ALU.eZ0Z_5 ));
    InMux I__5824 (
            .O(N__28850),
            .I(N__28847));
    LocalMux I__5823 (
            .O(N__28847),
            .I(N__28844));
    Span4Mux_h I__5822 (
            .O(N__28844),
            .I(N__28841));
    Odrv4 I__5821 (
            .O(N__28841),
            .I(\ALU.g_RNIRUBOZ0Z_0 ));
    InMux I__5820 (
            .O(N__28838),
            .I(N__28835));
    LocalMux I__5819 (
            .O(N__28835),
            .I(N__28832));
    Span4Mux_h I__5818 (
            .O(N__28832),
            .I(N__28829));
    Odrv4 I__5817 (
            .O(N__28829),
            .I(\ALU.d_RNIG6R7Z0Z_1 ));
    InMux I__5816 (
            .O(N__28826),
            .I(N__28823));
    LocalMux I__5815 (
            .O(N__28823),
            .I(N__28820));
    Span4Mux_h I__5814 (
            .O(N__28820),
            .I(N__28817));
    Span4Mux_v I__5813 (
            .O(N__28817),
            .I(N__28814));
    Odrv4 I__5812 (
            .O(N__28814),
            .I(\ALU.d_RNI45J9Z0Z_1 ));
    InMux I__5811 (
            .O(N__28811),
            .I(N__28808));
    LocalMux I__5810 (
            .O(N__28808),
            .I(\ALU.d_RNII8R7Z0Z_2 ));
    InMux I__5809 (
            .O(N__28805),
            .I(N__28802));
    LocalMux I__5808 (
            .O(N__28802),
            .I(N__28799));
    Span4Mux_h I__5807 (
            .O(N__28799),
            .I(N__28795));
    InMux I__5806 (
            .O(N__28798),
            .I(N__28792));
    Span4Mux_h I__5805 (
            .O(N__28795),
            .I(N__28789));
    LocalMux I__5804 (
            .O(N__28792),
            .I(N__28786));
    Odrv4 I__5803 (
            .O(N__28789),
            .I(\ALU.eZ0Z_7 ));
    Odrv12 I__5802 (
            .O(N__28786),
            .I(\ALU.eZ0Z_7 ));
    InMux I__5801 (
            .O(N__28781),
            .I(N__28777));
    InMux I__5800 (
            .O(N__28780),
            .I(N__28774));
    LocalMux I__5799 (
            .O(N__28777),
            .I(\ALU.eZ0Z_2 ));
    LocalMux I__5798 (
            .O(N__28774),
            .I(\ALU.eZ0Z_2 ));
    InMux I__5797 (
            .O(N__28769),
            .I(N__28766));
    LocalMux I__5796 (
            .O(N__28766),
            .I(N__28763));
    Span4Mux_h I__5795 (
            .O(N__28763),
            .I(N__28760));
    Span4Mux_v I__5794 (
            .O(N__28760),
            .I(N__28755));
    InMux I__5793 (
            .O(N__28759),
            .I(N__28752));
    InMux I__5792 (
            .O(N__28758),
            .I(N__28749));
    Odrv4 I__5791 (
            .O(N__28755),
            .I(a_2));
    LocalMux I__5790 (
            .O(N__28752),
            .I(a_2));
    LocalMux I__5789 (
            .O(N__28749),
            .I(a_2));
    CascadeMux I__5788 (
            .O(N__28742),
            .I(\ALU.g_RNIV2COZ0Z_2_cascade_ ));
    InMux I__5787 (
            .O(N__28739),
            .I(N__28736));
    LocalMux I__5786 (
            .O(N__28736),
            .I(\ALU.e_RNIRMVJZ0Z_2 ));
    CascadeMux I__5785 (
            .O(N__28733),
            .I(\ALU.operand2_7_ns_1_2_cascade_ ));
    InMux I__5784 (
            .O(N__28730),
            .I(N__28727));
    LocalMux I__5783 (
            .O(N__28727),
            .I(N__28723));
    InMux I__5782 (
            .O(N__28726),
            .I(N__28720));
    Span4Mux_h I__5781 (
            .O(N__28723),
            .I(N__28717));
    LocalMux I__5780 (
            .O(N__28720),
            .I(N__28714));
    Span4Mux_h I__5779 (
            .O(N__28717),
            .I(N__28711));
    Span4Mux_h I__5778 (
            .O(N__28714),
            .I(N__28708));
    Span4Mux_v I__5777 (
            .O(N__28711),
            .I(N__28703));
    Span4Mux_h I__5776 (
            .O(N__28708),
            .I(N__28703));
    Odrv4 I__5775 (
            .O(N__28703),
            .I(\ALU.operand2_2 ));
    InMux I__5774 (
            .O(N__28700),
            .I(N__28697));
    LocalMux I__5773 (
            .O(N__28697),
            .I(N__28694));
    Span4Mux_v I__5772 (
            .O(N__28694),
            .I(N__28691));
    Odrv4 I__5771 (
            .O(N__28691),
            .I(\ALU.un2_addsub_cry_12_c_RNIUL1GKZ0 ));
    CascadeMux I__5770 (
            .O(N__28688),
            .I(un2_addsub_cry_12_c_RNIG3PMU_cascade_));
    InMux I__5769 (
            .O(N__28685),
            .I(N__28682));
    LocalMux I__5768 (
            .O(N__28682),
            .I(N__28679));
    Span4Mux_v I__5767 (
            .O(N__28679),
            .I(N__28676));
    Span4Mux_v I__5766 (
            .O(N__28676),
            .I(N__28673));
    Odrv4 I__5765 (
            .O(N__28673),
            .I(c_RNI88B4N2_13));
    CascadeMux I__5764 (
            .O(N__28670),
            .I(aluOperation_RNI2J9SL3_0_cascade_));
    InMux I__5763 (
            .O(N__28667),
            .I(N__28664));
    LocalMux I__5762 (
            .O(N__28664),
            .I(N__28661));
    Span4Mux_v I__5761 (
            .O(N__28661),
            .I(N__28658));
    Odrv4 I__5760 (
            .O(N__28658),
            .I(\ALU.mult_2 ));
    InMux I__5759 (
            .O(N__28655),
            .I(N__28652));
    LocalMux I__5758 (
            .O(N__28652),
            .I(N__28649));
    Span4Mux_v I__5757 (
            .O(N__28649),
            .I(N__28646));
    Span4Mux_v I__5756 (
            .O(N__28646),
            .I(N__28643));
    Odrv4 I__5755 (
            .O(N__28643),
            .I(\ALU.a_15_m5_2 ));
    CascadeMux I__5754 (
            .O(N__28640),
            .I(\ALU.d_RNIIFMN04Z0Z_2_cascade_ ));
    InMux I__5753 (
            .O(N__28637),
            .I(N__28631));
    InMux I__5752 (
            .O(N__28636),
            .I(N__28631));
    LocalMux I__5751 (
            .O(N__28631),
            .I(N__28628));
    Span4Mux_h I__5750 (
            .O(N__28628),
            .I(N__28625));
    Odrv4 I__5749 (
            .O(N__28625),
            .I(\ALU.eZ0Z_3 ));
    InMux I__5748 (
            .O(N__28622),
            .I(N__28618));
    InMux I__5747 (
            .O(N__28621),
            .I(N__28615));
    LocalMux I__5746 (
            .O(N__28618),
            .I(N__28612));
    LocalMux I__5745 (
            .O(N__28615),
            .I(N__28609));
    Span4Mux_h I__5744 (
            .O(N__28612),
            .I(N__28606));
    Odrv4 I__5743 (
            .O(N__28609),
            .I(\ALU.eZ0Z_6 ));
    Odrv4 I__5742 (
            .O(N__28606),
            .I(\ALU.eZ0Z_6 ));
    InMux I__5741 (
            .O(N__28601),
            .I(N__28597));
    InMux I__5740 (
            .O(N__28600),
            .I(N__28594));
    LocalMux I__5739 (
            .O(N__28597),
            .I(N__28590));
    LocalMux I__5738 (
            .O(N__28594),
            .I(N__28587));
    InMux I__5737 (
            .O(N__28593),
            .I(N__28584));
    Span4Mux_v I__5736 (
            .O(N__28590),
            .I(N__28581));
    Span4Mux_v I__5735 (
            .O(N__28587),
            .I(N__28576));
    LocalMux I__5734 (
            .O(N__28584),
            .I(N__28576));
    Span4Mux_h I__5733 (
            .O(N__28581),
            .I(N__28573));
    Span4Mux_h I__5732 (
            .O(N__28576),
            .I(N__28570));
    Odrv4 I__5731 (
            .O(N__28573),
            .I(\ALU.eZ0Z_10 ));
    Odrv4 I__5730 (
            .O(N__28570),
            .I(\ALU.eZ0Z_10 ));
    InMux I__5729 (
            .O(N__28565),
            .I(N__28562));
    LocalMux I__5728 (
            .O(N__28562),
            .I(N__28558));
    InMux I__5727 (
            .O(N__28561),
            .I(N__28555));
    Span4Mux_h I__5726 (
            .O(N__28558),
            .I(N__28552));
    LocalMux I__5725 (
            .O(N__28555),
            .I(N__28549));
    Span4Mux_h I__5724 (
            .O(N__28552),
            .I(N__28544));
    Span4Mux_h I__5723 (
            .O(N__28549),
            .I(N__28544));
    Odrv4 I__5722 (
            .O(N__28544),
            .I(\ALU.eZ0Z_12 ));
    InMux I__5721 (
            .O(N__28541),
            .I(N__28538));
    LocalMux I__5720 (
            .O(N__28538),
            .I(N__28535));
    Span4Mux_v I__5719 (
            .O(N__28535),
            .I(N__28532));
    Span4Mux_h I__5718 (
            .O(N__28532),
            .I(N__28529));
    Odrv4 I__5717 (
            .O(N__28529),
            .I(\ALU.d_RNIPER7Z0Z_5 ));
    InMux I__5716 (
            .O(N__28526),
            .I(N__28522));
    InMux I__5715 (
            .O(N__28525),
            .I(N__28519));
    LocalMux I__5714 (
            .O(N__28522),
            .I(N__28515));
    LocalMux I__5713 (
            .O(N__28519),
            .I(N__28512));
    InMux I__5712 (
            .O(N__28518),
            .I(N__28509));
    Span4Mux_h I__5711 (
            .O(N__28515),
            .I(N__28506));
    Span4Mux_h I__5710 (
            .O(N__28512),
            .I(N__28503));
    LocalMux I__5709 (
            .O(N__28509),
            .I(\ALU.bZ0Z_10 ));
    Odrv4 I__5708 (
            .O(N__28506),
            .I(\ALU.bZ0Z_10 ));
    Odrv4 I__5707 (
            .O(N__28503),
            .I(\ALU.bZ0Z_10 ));
    InMux I__5706 (
            .O(N__28496),
            .I(N__28492));
    InMux I__5705 (
            .O(N__28495),
            .I(N__28489));
    LocalMux I__5704 (
            .O(N__28492),
            .I(N__28484));
    LocalMux I__5703 (
            .O(N__28489),
            .I(N__28484));
    Span4Mux_v I__5702 (
            .O(N__28484),
            .I(N__28481));
    Span4Mux_h I__5701 (
            .O(N__28481),
            .I(N__28478));
    Odrv4 I__5700 (
            .O(N__28478),
            .I(\ALU.bZ0Z_15 ));
    InMux I__5699 (
            .O(N__28475),
            .I(N__28472));
    LocalMux I__5698 (
            .O(N__28472),
            .I(N__28469));
    Span4Mux_h I__5697 (
            .O(N__28469),
            .I(N__28465));
    InMux I__5696 (
            .O(N__28468),
            .I(N__28462));
    Odrv4 I__5695 (
            .O(N__28465),
            .I(\ALU.fZ0Z_11 ));
    LocalMux I__5694 (
            .O(N__28462),
            .I(\ALU.fZ0Z_11 ));
    InMux I__5693 (
            .O(N__28457),
            .I(N__28454));
    LocalMux I__5692 (
            .O(N__28454),
            .I(N__28451));
    Span4Mux_v I__5691 (
            .O(N__28451),
            .I(N__28447));
    InMux I__5690 (
            .O(N__28450),
            .I(N__28444));
    Odrv4 I__5689 (
            .O(N__28447),
            .I(\ALU.bZ0Z_11 ));
    LocalMux I__5688 (
            .O(N__28444),
            .I(\ALU.bZ0Z_11 ));
    InMux I__5687 (
            .O(N__28439),
            .I(N__28436));
    LocalMux I__5686 (
            .O(N__28436),
            .I(N__28433));
    Span4Mux_h I__5685 (
            .O(N__28433),
            .I(N__28430));
    Odrv4 I__5684 (
            .O(N__28430),
            .I(\ALU.b_RNIKNSD1Z0Z_13 ));
    InMux I__5683 (
            .O(N__28427),
            .I(N__28423));
    InMux I__5682 (
            .O(N__28426),
            .I(N__28419));
    LocalMux I__5681 (
            .O(N__28423),
            .I(N__28416));
    InMux I__5680 (
            .O(N__28422),
            .I(N__28413));
    LocalMux I__5679 (
            .O(N__28419),
            .I(N__28408));
    Span4Mux_v I__5678 (
            .O(N__28416),
            .I(N__28408));
    LocalMux I__5677 (
            .O(N__28413),
            .I(N__28405));
    Span4Mux_v I__5676 (
            .O(N__28408),
            .I(N__28402));
    Span4Mux_h I__5675 (
            .O(N__28405),
            .I(N__28399));
    Odrv4 I__5674 (
            .O(N__28402),
            .I(\ALU.dZ0Z_10 ));
    Odrv4 I__5673 (
            .O(N__28399),
            .I(\ALU.dZ0Z_10 ));
    InMux I__5672 (
            .O(N__28394),
            .I(N__28391));
    LocalMux I__5671 (
            .O(N__28391),
            .I(N__28387));
    InMux I__5670 (
            .O(N__28390),
            .I(N__28384));
    Span4Mux_h I__5669 (
            .O(N__28387),
            .I(N__28381));
    LocalMux I__5668 (
            .O(N__28384),
            .I(N__28378));
    Span4Mux_h I__5667 (
            .O(N__28381),
            .I(N__28373));
    Span4Mux_h I__5666 (
            .O(N__28378),
            .I(N__28373));
    Odrv4 I__5665 (
            .O(N__28373),
            .I(\ALU.dZ0Z_12 ));
    InMux I__5664 (
            .O(N__28370),
            .I(N__28367));
    LocalMux I__5663 (
            .O(N__28367),
            .I(N__28364));
    Span4Mux_v I__5662 (
            .O(N__28364),
            .I(N__28360));
    InMux I__5661 (
            .O(N__28363),
            .I(N__28357));
    Span4Mux_h I__5660 (
            .O(N__28360),
            .I(N__28354));
    LocalMux I__5659 (
            .O(N__28357),
            .I(\ALU.bZ0Z_12 ));
    Odrv4 I__5658 (
            .O(N__28354),
            .I(\ALU.bZ0Z_12 ));
    CascadeMux I__5657 (
            .O(N__28349),
            .I(N__28346));
    InMux I__5656 (
            .O(N__28346),
            .I(N__28343));
    LocalMux I__5655 (
            .O(N__28343),
            .I(N__28339));
    InMux I__5654 (
            .O(N__28342),
            .I(N__28336));
    Span12Mux_s8_h I__5653 (
            .O(N__28339),
            .I(N__28333));
    LocalMux I__5652 (
            .O(N__28336),
            .I(\ALU.fZ0Z_12 ));
    Odrv12 I__5651 (
            .O(N__28333),
            .I(\ALU.fZ0Z_12 ));
    InMux I__5650 (
            .O(N__28328),
            .I(N__28325));
    LocalMux I__5649 (
            .O(N__28325),
            .I(\ALU.b_RNIILSD1Z0Z_12 ));
    CascadeMux I__5648 (
            .O(N__28322),
            .I(N__28319));
    InMux I__5647 (
            .O(N__28319),
            .I(N__28316));
    LocalMux I__5646 (
            .O(N__28316),
            .I(N__28313));
    Span4Mux_h I__5645 (
            .O(N__28313),
            .I(N__28310));
    Span4Mux_h I__5644 (
            .O(N__28310),
            .I(N__28306));
    InMux I__5643 (
            .O(N__28309),
            .I(N__28303));
    Odrv4 I__5642 (
            .O(N__28306),
            .I(\ALU.fZ0Z_14 ));
    LocalMux I__5641 (
            .O(N__28303),
            .I(\ALU.fZ0Z_14 ));
    InMux I__5640 (
            .O(N__28298),
            .I(N__28295));
    LocalMux I__5639 (
            .O(N__28295),
            .I(N__28292));
    Span4Mux_h I__5638 (
            .O(N__28292),
            .I(N__28289));
    Span4Mux_h I__5637 (
            .O(N__28289),
            .I(N__28285));
    InMux I__5636 (
            .O(N__28288),
            .I(N__28282));
    Odrv4 I__5635 (
            .O(N__28285),
            .I(\ALU.bZ0Z_14 ));
    LocalMux I__5634 (
            .O(N__28282),
            .I(\ALU.bZ0Z_14 ));
    CascadeMux I__5633 (
            .O(N__28277),
            .I(\ALU.g0_3_1_cascade_ ));
    InMux I__5632 (
            .O(N__28274),
            .I(N__28271));
    LocalMux I__5631 (
            .O(N__28271),
            .I(N__28268));
    Span4Mux_v I__5630 (
            .O(N__28268),
            .I(N__28265));
    Span4Mux_h I__5629 (
            .O(N__28265),
            .I(N__28262));
    Span4Mux_h I__5628 (
            .O(N__28262),
            .I(N__28259));
    Odrv4 I__5627 (
            .O(N__28259),
            .I(\ALU.N_703_0_0 ));
    InMux I__5626 (
            .O(N__28256),
            .I(N__28253));
    LocalMux I__5625 (
            .O(N__28253),
            .I(\ALU.N_4 ));
    CascadeMux I__5624 (
            .O(N__28250),
            .I(N__28247));
    InMux I__5623 (
            .O(N__28247),
            .I(N__28244));
    LocalMux I__5622 (
            .O(N__28244),
            .I(N__28241));
    Odrv4 I__5621 (
            .O(N__28241),
            .I(\ALU.N_5 ));
    CascadeMux I__5620 (
            .O(N__28238),
            .I(\ALU.a_15_m4_12_cascade_ ));
    InMux I__5619 (
            .O(N__28235),
            .I(N__28232));
    LocalMux I__5618 (
            .O(N__28232),
            .I(N__28229));
    Span4Mux_h I__5617 (
            .O(N__28229),
            .I(N__28226));
    Odrv4 I__5616 (
            .O(N__28226),
            .I(\ALU.un2_addsub_cry_11_c_RNII7OFZ0Z9 ));
    CascadeMux I__5615 (
            .O(N__28223),
            .I(un2_addsub_cry_11_c_RNIQ9LMU_cascade_));
    InMux I__5614 (
            .O(N__28220),
            .I(N__28217));
    LocalMux I__5613 (
            .O(N__28217),
            .I(c_RNIC8RDN2_12));
    CascadeMux I__5612 (
            .O(N__28214),
            .I(aluOperation_RNIGPL5M3_0_cascade_));
    InMux I__5611 (
            .O(N__28211),
            .I(N__28208));
    LocalMux I__5610 (
            .O(N__28208),
            .I(N__28204));
    InMux I__5609 (
            .O(N__28207),
            .I(N__28201));
    Odrv12 I__5608 (
            .O(N__28204),
            .I(\ALU.aZ0Z_12 ));
    LocalMux I__5607 (
            .O(N__28201),
            .I(\ALU.aZ0Z_12 ));
    InMux I__5606 (
            .O(N__28196),
            .I(N__28193));
    LocalMux I__5605 (
            .O(N__28193),
            .I(N__28190));
    Odrv12 I__5604 (
            .O(N__28190),
            .I(\ALU.N_271_0 ));
    InMux I__5603 (
            .O(N__28187),
            .I(N__28184));
    LocalMux I__5602 (
            .O(N__28184),
            .I(\ALU.a_15_m3_12 ));
    InMux I__5601 (
            .O(N__28181),
            .I(N__28178));
    LocalMux I__5600 (
            .O(N__28178),
            .I(N__28175));
    Span4Mux_v I__5599 (
            .O(N__28175),
            .I(N__28172));
    Span4Mux_h I__5598 (
            .O(N__28172),
            .I(N__28169));
    Odrv4 I__5597 (
            .O(N__28169),
            .I(\ALU.N_314 ));
    InMux I__5596 (
            .O(N__28166),
            .I(N__28163));
    LocalMux I__5595 (
            .O(N__28163),
            .I(\ALU.lshift_12 ));
    InMux I__5594 (
            .O(N__28160),
            .I(N__28155));
    CascadeMux I__5593 (
            .O(N__28159),
            .I(N__28152));
    CascadeMux I__5592 (
            .O(N__28158),
            .I(N__28149));
    LocalMux I__5591 (
            .O(N__28155),
            .I(N__28146));
    InMux I__5590 (
            .O(N__28152),
            .I(N__28141));
    InMux I__5589 (
            .O(N__28149),
            .I(N__28141));
    Span4Mux_v I__5588 (
            .O(N__28146),
            .I(N__28138));
    LocalMux I__5587 (
            .O(N__28141),
            .I(\ALU.fZ0Z_9 ));
    Odrv4 I__5586 (
            .O(N__28138),
            .I(\ALU.fZ0Z_9 ));
    InMux I__5585 (
            .O(N__28133),
            .I(N__28130));
    LocalMux I__5584 (
            .O(N__28130),
            .I(N__28127));
    Span4Mux_v I__5583 (
            .O(N__28127),
            .I(N__28122));
    InMux I__5582 (
            .O(N__28126),
            .I(N__28117));
    InMux I__5581 (
            .O(N__28125),
            .I(N__28117));
    Span4Mux_h I__5580 (
            .O(N__28122),
            .I(N__28114));
    LocalMux I__5579 (
            .O(N__28117),
            .I(\ALU.bZ0Z_9 ));
    Odrv4 I__5578 (
            .O(N__28114),
            .I(\ALU.bZ0Z_9 ));
    InMux I__5577 (
            .O(N__28109),
            .I(N__28106));
    LocalMux I__5576 (
            .O(N__28106),
            .I(N__28103));
    Odrv12 I__5575 (
            .O(N__28103),
            .I(\ALU.f_RNIUUJ01Z0Z_9 ));
    CascadeMux I__5574 (
            .O(N__28100),
            .I(\ALU.a_15_m2_ns_1Z0Z_5_cascade_ ));
    InMux I__5573 (
            .O(N__28097),
            .I(N__28094));
    LocalMux I__5572 (
            .O(N__28094),
            .I(N__28091));
    Span4Mux_v I__5571 (
            .O(N__28091),
            .I(N__28081));
    InMux I__5570 (
            .O(N__28090),
            .I(N__28078));
    InMux I__5569 (
            .O(N__28089),
            .I(N__28075));
    CascadeMux I__5568 (
            .O(N__28088),
            .I(N__28072));
    InMux I__5567 (
            .O(N__28087),
            .I(N__28065));
    InMux I__5566 (
            .O(N__28086),
            .I(N__28060));
    InMux I__5565 (
            .O(N__28085),
            .I(N__28060));
    InMux I__5564 (
            .O(N__28084),
            .I(N__28057));
    Span4Mux_v I__5563 (
            .O(N__28081),
            .I(N__28050));
    LocalMux I__5562 (
            .O(N__28078),
            .I(N__28050));
    LocalMux I__5561 (
            .O(N__28075),
            .I(N__28050));
    InMux I__5560 (
            .O(N__28072),
            .I(N__28047));
    InMux I__5559 (
            .O(N__28071),
            .I(N__28044));
    InMux I__5558 (
            .O(N__28070),
            .I(N__28041));
    InMux I__5557 (
            .O(N__28069),
            .I(N__28036));
    InMux I__5556 (
            .O(N__28068),
            .I(N__28036));
    LocalMux I__5555 (
            .O(N__28065),
            .I(N__28031));
    LocalMux I__5554 (
            .O(N__28060),
            .I(N__28028));
    LocalMux I__5553 (
            .O(N__28057),
            .I(N__28020));
    Span4Mux_h I__5552 (
            .O(N__28050),
            .I(N__28020));
    LocalMux I__5551 (
            .O(N__28047),
            .I(N__28015));
    LocalMux I__5550 (
            .O(N__28044),
            .I(N__28015));
    LocalMux I__5549 (
            .O(N__28041),
            .I(N__28010));
    LocalMux I__5548 (
            .O(N__28036),
            .I(N__28010));
    InMux I__5547 (
            .O(N__28035),
            .I(N__28007));
    InMux I__5546 (
            .O(N__28034),
            .I(N__28004));
    Span4Mux_v I__5545 (
            .O(N__28031),
            .I(N__27999));
    Span4Mux_v I__5544 (
            .O(N__28028),
            .I(N__27999));
    InMux I__5543 (
            .O(N__28027),
            .I(N__27996));
    InMux I__5542 (
            .O(N__28026),
            .I(N__27991));
    InMux I__5541 (
            .O(N__28025),
            .I(N__27991));
    Span4Mux_h I__5540 (
            .O(N__28020),
            .I(N__27988));
    Span4Mux_v I__5539 (
            .O(N__28015),
            .I(N__27983));
    Span4Mux_h I__5538 (
            .O(N__28010),
            .I(N__27983));
    LocalMux I__5537 (
            .O(N__28007),
            .I(\ALU.N_225_0 ));
    LocalMux I__5536 (
            .O(N__28004),
            .I(\ALU.N_225_0 ));
    Odrv4 I__5535 (
            .O(N__27999),
            .I(\ALU.N_225_0 ));
    LocalMux I__5534 (
            .O(N__27996),
            .I(\ALU.N_225_0 ));
    LocalMux I__5533 (
            .O(N__27991),
            .I(\ALU.N_225_0 ));
    Odrv4 I__5532 (
            .O(N__27988),
            .I(\ALU.N_225_0 ));
    Odrv4 I__5531 (
            .O(N__27983),
            .I(\ALU.N_225_0 ));
    CascadeMux I__5530 (
            .O(N__27968),
            .I(\ALU.a_15_m2_5_cascade_ ));
    InMux I__5529 (
            .O(N__27965),
            .I(N__27962));
    LocalMux I__5528 (
            .O(N__27962),
            .I(N__27959));
    Span4Mux_h I__5527 (
            .O(N__27959),
            .I(N__27955));
    InMux I__5526 (
            .O(N__27958),
            .I(N__27952));
    Odrv4 I__5525 (
            .O(N__27955),
            .I(\ALU.N_420 ));
    LocalMux I__5524 (
            .O(N__27952),
            .I(\ALU.N_420 ));
    InMux I__5523 (
            .O(N__27947),
            .I(N__27944));
    LocalMux I__5522 (
            .O(N__27944),
            .I(\ALU.a_15_m4_5 ));
    InMux I__5521 (
            .O(N__27941),
            .I(N__27937));
    InMux I__5520 (
            .O(N__27940),
            .I(N__27934));
    LocalMux I__5519 (
            .O(N__27937),
            .I(N__27931));
    LocalMux I__5518 (
            .O(N__27934),
            .I(N__27928));
    Span4Mux_h I__5517 (
            .O(N__27931),
            .I(N__27925));
    Span12Mux_h I__5516 (
            .O(N__27928),
            .I(N__27921));
    Span4Mux_v I__5515 (
            .O(N__27925),
            .I(N__27918));
    InMux I__5514 (
            .O(N__27924),
            .I(N__27915));
    Odrv12 I__5513 (
            .O(N__27921),
            .I(a_4));
    Odrv4 I__5512 (
            .O(N__27918),
            .I(a_4));
    LocalMux I__5511 (
            .O(N__27915),
            .I(a_4));
    InMux I__5510 (
            .O(N__27908),
            .I(N__27905));
    LocalMux I__5509 (
            .O(N__27905),
            .I(N__27902));
    Span4Mux_v I__5508 (
            .O(N__27902),
            .I(N__27899));
    Sp12to4 I__5507 (
            .O(N__27899),
            .I(N__27894));
    InMux I__5506 (
            .O(N__27898),
            .I(N__27891));
    InMux I__5505 (
            .O(N__27897),
            .I(N__27888));
    Span12Mux_s8_h I__5504 (
            .O(N__27894),
            .I(N__27883));
    LocalMux I__5503 (
            .O(N__27891),
            .I(N__27883));
    LocalMux I__5502 (
            .O(N__27888),
            .I(N__27880));
    Odrv12 I__5501 (
            .O(N__27883),
            .I(a_6));
    Odrv4 I__5500 (
            .O(N__27880),
            .I(a_6));
    InMux I__5499 (
            .O(N__27875),
            .I(N__27871));
    InMux I__5498 (
            .O(N__27874),
            .I(N__27867));
    LocalMux I__5497 (
            .O(N__27871),
            .I(N__27864));
    InMux I__5496 (
            .O(N__27870),
            .I(N__27861));
    LocalMux I__5495 (
            .O(N__27867),
            .I(N__27858));
    Span4Mux_h I__5494 (
            .O(N__27864),
            .I(N__27855));
    LocalMux I__5493 (
            .O(N__27861),
            .I(N__27852));
    Span12Mux_v I__5492 (
            .O(N__27858),
            .I(N__27849));
    Span4Mux_h I__5491 (
            .O(N__27855),
            .I(N__27846));
    Span4Mux_h I__5490 (
            .O(N__27852),
            .I(N__27843));
    Odrv12 I__5489 (
            .O(N__27849),
            .I(a_7));
    Odrv4 I__5488 (
            .O(N__27846),
            .I(a_7));
    Odrv4 I__5487 (
            .O(N__27843),
            .I(a_7));
    InMux I__5486 (
            .O(N__27836),
            .I(N__27833));
    LocalMux I__5485 (
            .O(N__27833),
            .I(N__27830));
    Odrv4 I__5484 (
            .O(N__27830),
            .I(\ALU.a_15_m2_12 ));
    InMux I__5483 (
            .O(N__27827),
            .I(N__27824));
    LocalMux I__5482 (
            .O(N__27824),
            .I(\ALU.rshift_15_ns_1_7 ));
    CascadeMux I__5481 (
            .O(N__27821),
            .I(\ALU.rshift_3_ns_1_3_cascade_ ));
    CascadeMux I__5480 (
            .O(N__27818),
            .I(\ALU.N_471_cascade_ ));
    InMux I__5479 (
            .O(N__27815),
            .I(N__27812));
    LocalMux I__5478 (
            .O(N__27812),
            .I(\ALU.N_475 ));
    InMux I__5477 (
            .O(N__27809),
            .I(N__27806));
    LocalMux I__5476 (
            .O(N__27806),
            .I(\ALU.rshift_3_ns_1_7 ));
    InMux I__5475 (
            .O(N__27803),
            .I(N__27797));
    InMux I__5474 (
            .O(N__27802),
            .I(N__27797));
    LocalMux I__5473 (
            .O(N__27797),
            .I(\ALU.N_576 ));
    CascadeMux I__5472 (
            .O(N__27794),
            .I(\ALU.a_15_m5_5_cascade_ ));
    InMux I__5471 (
            .O(N__27791),
            .I(N__27788));
    LocalMux I__5470 (
            .O(N__27788),
            .I(N__27785));
    Span4Mux_h I__5469 (
            .O(N__27785),
            .I(N__27782));
    Span4Mux_v I__5468 (
            .O(N__27782),
            .I(N__27779));
    Odrv4 I__5467 (
            .O(N__27779),
            .I(\ALU.mult_5 ));
    InMux I__5466 (
            .O(N__27776),
            .I(N__27773));
    LocalMux I__5465 (
            .O(N__27773),
            .I(N__27770));
    Odrv4 I__5464 (
            .O(N__27770),
            .I(\ALU.d_RNIPFIBI1Z0Z_9 ));
    CascadeMux I__5463 (
            .O(N__27767),
            .I(\ALU.dout_3_ns_1_6_cascade_ ));
    InMux I__5462 (
            .O(N__27764),
            .I(N__27761));
    LocalMux I__5461 (
            .O(N__27761),
            .I(\ALU.N_705 ));
    InMux I__5460 (
            .O(N__27758),
            .I(N__27755));
    LocalMux I__5459 (
            .O(N__27755),
            .I(N__27752));
    Span4Mux_v I__5458 (
            .O(N__27752),
            .I(N__27749));
    Span4Mux_v I__5457 (
            .O(N__27749),
            .I(N__27746));
    Span4Mux_v I__5456 (
            .O(N__27746),
            .I(N__27742));
    CascadeMux I__5455 (
            .O(N__27745),
            .I(N__27739));
    Sp12to4 I__5454 (
            .O(N__27742),
            .I(N__27736));
    InMux I__5453 (
            .O(N__27739),
            .I(N__27733));
    Odrv12 I__5452 (
            .O(N__27736),
            .I(testWordZ0Z_7));
    LocalMux I__5451 (
            .O(N__27733),
            .I(testWordZ0Z_7));
    CEMux I__5450 (
            .O(N__27728),
            .I(N__27724));
    CEMux I__5449 (
            .O(N__27727),
            .I(N__27720));
    LocalMux I__5448 (
            .O(N__27724),
            .I(N__27716));
    CEMux I__5447 (
            .O(N__27723),
            .I(N__27713));
    LocalMux I__5446 (
            .O(N__27720),
            .I(N__27710));
    CEMux I__5445 (
            .O(N__27719),
            .I(N__27707));
    Span4Mux_h I__5444 (
            .O(N__27716),
            .I(N__27704));
    LocalMux I__5443 (
            .O(N__27713),
            .I(N__27701));
    Span4Mux_v I__5442 (
            .O(N__27710),
            .I(N__27698));
    LocalMux I__5441 (
            .O(N__27707),
            .I(N__27694));
    Span4Mux_h I__5440 (
            .O(N__27704),
            .I(N__27691));
    Span4Mux_h I__5439 (
            .O(N__27701),
            .I(N__27688));
    Span4Mux_h I__5438 (
            .O(N__27698),
            .I(N__27685));
    CEMux I__5437 (
            .O(N__27697),
            .I(N__27682));
    Span4Mux_h I__5436 (
            .O(N__27694),
            .I(N__27679));
    Span4Mux_v I__5435 (
            .O(N__27691),
            .I(N__27674));
    Span4Mux_h I__5434 (
            .O(N__27688),
            .I(N__27674));
    IoSpan4Mux I__5433 (
            .O(N__27685),
            .I(N__27671));
    LocalMux I__5432 (
            .O(N__27682),
            .I(N__27668));
    Span4Mux_h I__5431 (
            .O(N__27679),
            .I(N__27665));
    Span4Mux_v I__5430 (
            .O(N__27674),
            .I(N__27662));
    IoSpan4Mux I__5429 (
            .O(N__27671),
            .I(N__27659));
    Span4Mux_v I__5428 (
            .O(N__27668),
            .I(N__27656));
    Span4Mux_s2_h I__5427 (
            .O(N__27665),
            .I(N__27653));
    Span4Mux_v I__5426 (
            .O(N__27662),
            .I(N__27650));
    IoSpan4Mux I__5425 (
            .O(N__27659),
            .I(N__27645));
    Span4Mux_h I__5424 (
            .O(N__27656),
            .I(N__27645));
    Span4Mux_v I__5423 (
            .O(N__27653),
            .I(N__27642));
    Span4Mux_h I__5422 (
            .O(N__27650),
            .I(N__27639));
    Span4Mux_s3_h I__5421 (
            .O(N__27645),
            .I(N__27636));
    Span4Mux_v I__5420 (
            .O(N__27642),
            .I(N__27633));
    Span4Mux_h I__5419 (
            .O(N__27639),
            .I(N__27630));
    Span4Mux_v I__5418 (
            .O(N__27636),
            .I(N__27627));
    Odrv4 I__5417 (
            .O(N__27633),
            .I(\CONTROL.operand1_cnvZ0Z_0 ));
    Odrv4 I__5416 (
            .O(N__27630),
            .I(\CONTROL.operand1_cnvZ0Z_0 ));
    Odrv4 I__5415 (
            .O(N__27627),
            .I(\CONTROL.operand1_cnvZ0Z_0 ));
    CascadeMux I__5414 (
            .O(N__27620),
            .I(\ALU.c_RNI72MICZ0Z_15_cascade_ ));
    InMux I__5413 (
            .O(N__27617),
            .I(N__27614));
    LocalMux I__5412 (
            .O(N__27614),
            .I(N__27611));
    Odrv4 I__5411 (
            .O(N__27611),
            .I(\ALU.d_RNI4HG101Z0Z_7 ));
    InMux I__5410 (
            .O(N__27608),
            .I(N__27604));
    InMux I__5409 (
            .O(N__27607),
            .I(N__27590));
    LocalMux I__5408 (
            .O(N__27604),
            .I(N__27583));
    InMux I__5407 (
            .O(N__27603),
            .I(N__27580));
    InMux I__5406 (
            .O(N__27602),
            .I(N__27577));
    InMux I__5405 (
            .O(N__27601),
            .I(N__27570));
    InMux I__5404 (
            .O(N__27600),
            .I(N__27570));
    InMux I__5403 (
            .O(N__27599),
            .I(N__27570));
    InMux I__5402 (
            .O(N__27598),
            .I(N__27567));
    InMux I__5401 (
            .O(N__27597),
            .I(N__27559));
    InMux I__5400 (
            .O(N__27596),
            .I(N__27559));
    InMux I__5399 (
            .O(N__27595),
            .I(N__27559));
    CascadeMux I__5398 (
            .O(N__27594),
            .I(N__27555));
    InMux I__5397 (
            .O(N__27593),
            .I(N__27551));
    LocalMux I__5396 (
            .O(N__27590),
            .I(N__27547));
    InMux I__5395 (
            .O(N__27589),
            .I(N__27544));
    InMux I__5394 (
            .O(N__27588),
            .I(N__27541));
    InMux I__5393 (
            .O(N__27587),
            .I(N__27536));
    CascadeMux I__5392 (
            .O(N__27586),
            .I(N__27531));
    Span4Mux_s3_v I__5391 (
            .O(N__27583),
            .I(N__27526));
    LocalMux I__5390 (
            .O(N__27580),
            .I(N__27526));
    LocalMux I__5389 (
            .O(N__27577),
            .I(N__27521));
    LocalMux I__5388 (
            .O(N__27570),
            .I(N__27521));
    LocalMux I__5387 (
            .O(N__27567),
            .I(N__27518));
    InMux I__5386 (
            .O(N__27566),
            .I(N__27515));
    LocalMux I__5385 (
            .O(N__27559),
            .I(N__27512));
    InMux I__5384 (
            .O(N__27558),
            .I(N__27508));
    InMux I__5383 (
            .O(N__27555),
            .I(N__27503));
    InMux I__5382 (
            .O(N__27554),
            .I(N__27503));
    LocalMux I__5381 (
            .O(N__27551),
            .I(N__27500));
    InMux I__5380 (
            .O(N__27550),
            .I(N__27496));
    Span4Mux_v I__5379 (
            .O(N__27547),
            .I(N__27493));
    LocalMux I__5378 (
            .O(N__27544),
            .I(N__27488));
    LocalMux I__5377 (
            .O(N__27541),
            .I(N__27488));
    InMux I__5376 (
            .O(N__27540),
            .I(N__27485));
    InMux I__5375 (
            .O(N__27539),
            .I(N__27482));
    LocalMux I__5374 (
            .O(N__27536),
            .I(N__27479));
    InMux I__5373 (
            .O(N__27535),
            .I(N__27472));
    InMux I__5372 (
            .O(N__27534),
            .I(N__27472));
    InMux I__5371 (
            .O(N__27531),
            .I(N__27472));
    Span4Mux_v I__5370 (
            .O(N__27526),
            .I(N__27469));
    Span4Mux_v I__5369 (
            .O(N__27521),
            .I(N__27466));
    Span4Mux_h I__5368 (
            .O(N__27518),
            .I(N__27463));
    LocalMux I__5367 (
            .O(N__27515),
            .I(N__27460));
    Span4Mux_v I__5366 (
            .O(N__27512),
            .I(N__27457));
    InMux I__5365 (
            .O(N__27511),
            .I(N__27454));
    LocalMux I__5364 (
            .O(N__27508),
            .I(N__27451));
    LocalMux I__5363 (
            .O(N__27503),
            .I(N__27446));
    Span4Mux_v I__5362 (
            .O(N__27500),
            .I(N__27446));
    InMux I__5361 (
            .O(N__27499),
            .I(N__27443));
    LocalMux I__5360 (
            .O(N__27496),
            .I(N__27436));
    Span4Mux_h I__5359 (
            .O(N__27493),
            .I(N__27436));
    Span4Mux_v I__5358 (
            .O(N__27488),
            .I(N__27436));
    LocalMux I__5357 (
            .O(N__27485),
            .I(N__27431));
    LocalMux I__5356 (
            .O(N__27482),
            .I(N__27431));
    Span4Mux_v I__5355 (
            .O(N__27479),
            .I(N__27428));
    LocalMux I__5354 (
            .O(N__27472),
            .I(N__27425));
    Span4Mux_v I__5353 (
            .O(N__27469),
            .I(N__27414));
    Span4Mux_h I__5352 (
            .O(N__27466),
            .I(N__27414));
    Span4Mux_v I__5351 (
            .O(N__27463),
            .I(N__27414));
    Span4Mux_v I__5350 (
            .O(N__27460),
            .I(N__27414));
    Span4Mux_h I__5349 (
            .O(N__27457),
            .I(N__27414));
    LocalMux I__5348 (
            .O(N__27454),
            .I(N__27405));
    Span4Mux_v I__5347 (
            .O(N__27451),
            .I(N__27405));
    Span4Mux_h I__5346 (
            .O(N__27446),
            .I(N__27405));
    LocalMux I__5345 (
            .O(N__27443),
            .I(N__27405));
    Span4Mux_v I__5344 (
            .O(N__27436),
            .I(N__27400));
    Span4Mux_h I__5343 (
            .O(N__27431),
            .I(N__27400));
    Span4Mux_v I__5342 (
            .O(N__27428),
            .I(N__27395));
    Span4Mux_s3_h I__5341 (
            .O(N__27425),
            .I(N__27395));
    Odrv4 I__5340 (
            .O(N__27414),
            .I(\ALU.aluOut_10 ));
    Odrv4 I__5339 (
            .O(N__27405),
            .I(\ALU.aluOut_10 ));
    Odrv4 I__5338 (
            .O(N__27400),
            .I(\ALU.aluOut_10 ));
    Odrv4 I__5337 (
            .O(N__27395),
            .I(\ALU.aluOut_10 ));
    CascadeMux I__5336 (
            .O(N__27386),
            .I(\ALU.N_475_cascade_ ));
    InMux I__5335 (
            .O(N__27383),
            .I(N__27380));
    LocalMux I__5334 (
            .O(N__27380),
            .I(\ALU.rshift_7 ));
    InMux I__5333 (
            .O(N__27377),
            .I(N__27374));
    LocalMux I__5332 (
            .O(N__27374),
            .I(N__27371));
    Span4Mux_h I__5331 (
            .O(N__27371),
            .I(N__27368));
    Odrv4 I__5330 (
            .O(N__27368),
            .I(\ALU.g_RNI0MJNZ0Z_1 ));
    InMux I__5329 (
            .O(N__27365),
            .I(N__27362));
    LocalMux I__5328 (
            .O(N__27362),
            .I(N__27359));
    Span4Mux_h I__5327 (
            .O(N__27359),
            .I(N__27356));
    Odrv4 I__5326 (
            .O(N__27356),
            .I(\ALU.dout_6_ns_1_3 ));
    CascadeMux I__5325 (
            .O(N__27353),
            .I(N__27350));
    InMux I__5324 (
            .O(N__27350),
            .I(N__27345));
    InMux I__5323 (
            .O(N__27349),
            .I(N__27342));
    CascadeMux I__5322 (
            .O(N__27348),
            .I(N__27339));
    LocalMux I__5321 (
            .O(N__27345),
            .I(N__27331));
    LocalMux I__5320 (
            .O(N__27342),
            .I(N__27331));
    InMux I__5319 (
            .O(N__27339),
            .I(N__27326));
    InMux I__5318 (
            .O(N__27338),
            .I(N__27326));
    CascadeMux I__5317 (
            .O(N__27337),
            .I(N__27322));
    InMux I__5316 (
            .O(N__27336),
            .I(N__27318));
    Span4Mux_v I__5315 (
            .O(N__27331),
            .I(N__27315));
    LocalMux I__5314 (
            .O(N__27326),
            .I(N__27312));
    InMux I__5313 (
            .O(N__27325),
            .I(N__27309));
    InMux I__5312 (
            .O(N__27322),
            .I(N__27304));
    InMux I__5311 (
            .O(N__27321),
            .I(N__27304));
    LocalMux I__5310 (
            .O(N__27318),
            .I(N__27299));
    Sp12to4 I__5309 (
            .O(N__27315),
            .I(N__27299));
    Span4Mux_h I__5308 (
            .O(N__27312),
            .I(N__27296));
    LocalMux I__5307 (
            .O(N__27309),
            .I(aluOperand1_2_rep1));
    LocalMux I__5306 (
            .O(N__27304),
            .I(aluOperand1_2_rep1));
    Odrv12 I__5305 (
            .O(N__27299),
            .I(aluOperand1_2_rep1));
    Odrv4 I__5304 (
            .O(N__27296),
            .I(aluOperand1_2_rep1));
    InMux I__5303 (
            .O(N__27287),
            .I(N__27284));
    LocalMux I__5302 (
            .O(N__27284),
            .I(N__27281));
    Span4Mux_h I__5301 (
            .O(N__27281),
            .I(N__27278));
    Odrv4 I__5300 (
            .O(N__27278),
            .I(\ALU.dout_6_ns_1_4 ));
    InMux I__5299 (
            .O(N__27275),
            .I(N__27272));
    LocalMux I__5298 (
            .O(N__27272),
            .I(N__27269));
    Span4Mux_h I__5297 (
            .O(N__27269),
            .I(N__27266));
    Odrv4 I__5296 (
            .O(N__27266),
            .I(\ALU.N_747 ));
    InMux I__5295 (
            .O(N__27263),
            .I(N__27260));
    LocalMux I__5294 (
            .O(N__27260),
            .I(N__27257));
    Span4Mux_v I__5293 (
            .O(N__27257),
            .I(N__27253));
    InMux I__5292 (
            .O(N__27256),
            .I(N__27250));
    Odrv4 I__5291 (
            .O(N__27253),
            .I(\ALU.N_699 ));
    LocalMux I__5290 (
            .O(N__27250),
            .I(\ALU.N_699 ));
    InMux I__5289 (
            .O(N__27245),
            .I(N__27242));
    LocalMux I__5288 (
            .O(N__27242),
            .I(N__27239));
    Span4Mux_v I__5287 (
            .O(N__27239),
            .I(N__27236));
    Span4Mux_v I__5286 (
            .O(N__27236),
            .I(N__27232));
    InMux I__5285 (
            .O(N__27235),
            .I(N__27229));
    Span4Mux_v I__5284 (
            .O(N__27232),
            .I(N__27226));
    LocalMux I__5283 (
            .O(N__27229),
            .I(N__27223));
    Span4Mux_h I__5282 (
            .O(N__27226),
            .I(N__27220));
    Span12Mux_s10_v I__5281 (
            .O(N__27223),
            .I(N__27217));
    Odrv4 I__5280 (
            .O(N__27220),
            .I(\ALU.N_404_1 ));
    Odrv12 I__5279 (
            .O(N__27217),
            .I(\ALU.N_404_1 ));
    CascadeMux I__5278 (
            .O(N__27212),
            .I(N__27209));
    InMux I__5277 (
            .O(N__27209),
            .I(N__27206));
    LocalMux I__5276 (
            .O(N__27206),
            .I(N__27203));
    Odrv4 I__5275 (
            .O(N__27203),
            .I(\ALU.dout_6_ns_1_6 ));
    CascadeMux I__5274 (
            .O(N__27200),
            .I(\ALU.N_753_cascade_ ));
    InMux I__5273 (
            .O(N__27197),
            .I(N__27192));
    InMux I__5272 (
            .O(N__27196),
            .I(N__27189));
    InMux I__5271 (
            .O(N__27195),
            .I(N__27186));
    LocalMux I__5270 (
            .O(N__27192),
            .I(N__27182));
    LocalMux I__5269 (
            .O(N__27189),
            .I(N__27177));
    LocalMux I__5268 (
            .O(N__27186),
            .I(N__27177));
    InMux I__5267 (
            .O(N__27185),
            .I(N__27174));
    Span4Mux_v I__5266 (
            .O(N__27182),
            .I(N__27171));
    Span4Mux_v I__5265 (
            .O(N__27177),
            .I(N__27168));
    LocalMux I__5264 (
            .O(N__27174),
            .I(N__27165));
    Span4Mux_h I__5263 (
            .O(N__27171),
            .I(N__27162));
    Span4Mux_h I__5262 (
            .O(N__27168),
            .I(N__27159));
    Span4Mux_h I__5261 (
            .O(N__27165),
            .I(N__27156));
    Span4Mux_h I__5260 (
            .O(N__27162),
            .I(N__27148));
    Span4Mux_h I__5259 (
            .O(N__27159),
            .I(N__27148));
    Span4Mux_h I__5258 (
            .O(N__27156),
            .I(N__27148));
    InMux I__5257 (
            .O(N__27155),
            .I(N__27145));
    Span4Mux_v I__5256 (
            .O(N__27148),
            .I(N__27142));
    LocalMux I__5255 (
            .O(N__27145),
            .I(N__27139));
    Odrv4 I__5254 (
            .O(N__27142),
            .I(testWordZ0Z_9));
    Odrv4 I__5253 (
            .O(N__27139),
            .I(testWordZ0Z_9));
    InMux I__5252 (
            .O(N__27134),
            .I(N__27121));
    InMux I__5251 (
            .O(N__27133),
            .I(N__27117));
    InMux I__5250 (
            .O(N__27132),
            .I(N__27114));
    InMux I__5249 (
            .O(N__27131),
            .I(N__27109));
    InMux I__5248 (
            .O(N__27130),
            .I(N__27109));
    InMux I__5247 (
            .O(N__27129),
            .I(N__27103));
    InMux I__5246 (
            .O(N__27128),
            .I(N__27103));
    InMux I__5245 (
            .O(N__27127),
            .I(N__27100));
    InMux I__5244 (
            .O(N__27126),
            .I(N__27097));
    InMux I__5243 (
            .O(N__27125),
            .I(N__27092));
    InMux I__5242 (
            .O(N__27124),
            .I(N__27092));
    LocalMux I__5241 (
            .O(N__27121),
            .I(N__27089));
    CascadeMux I__5240 (
            .O(N__27120),
            .I(N__27086));
    LocalMux I__5239 (
            .O(N__27117),
            .I(N__27083));
    LocalMux I__5238 (
            .O(N__27114),
            .I(N__27078));
    LocalMux I__5237 (
            .O(N__27109),
            .I(N__27078));
    InMux I__5236 (
            .O(N__27108),
            .I(N__27075));
    LocalMux I__5235 (
            .O(N__27103),
            .I(N__27072));
    LocalMux I__5234 (
            .O(N__27100),
            .I(N__27069));
    LocalMux I__5233 (
            .O(N__27097),
            .I(N__27062));
    LocalMux I__5232 (
            .O(N__27092),
            .I(N__27062));
    Span4Mux_v I__5231 (
            .O(N__27089),
            .I(N__27062));
    InMux I__5230 (
            .O(N__27086),
            .I(N__27059));
    Span4Mux_v I__5229 (
            .O(N__27083),
            .I(N__27054));
    Span4Mux_h I__5228 (
            .O(N__27078),
            .I(N__27054));
    LocalMux I__5227 (
            .O(N__27075),
            .I(aluOperand1_fast_1));
    Odrv4 I__5226 (
            .O(N__27072),
            .I(aluOperand1_fast_1));
    Odrv12 I__5225 (
            .O(N__27069),
            .I(aluOperand1_fast_1));
    Odrv4 I__5224 (
            .O(N__27062),
            .I(aluOperand1_fast_1));
    LocalMux I__5223 (
            .O(N__27059),
            .I(aluOperand1_fast_1));
    Odrv4 I__5222 (
            .O(N__27054),
            .I(aluOperand1_fast_1));
    CascadeMux I__5221 (
            .O(N__27041),
            .I(N__27036));
    CascadeMux I__5220 (
            .O(N__27040),
            .I(N__27033));
    CascadeMux I__5219 (
            .O(N__27039),
            .I(N__27030));
    InMux I__5218 (
            .O(N__27036),
            .I(N__27021));
    InMux I__5217 (
            .O(N__27033),
            .I(N__27021));
    InMux I__5216 (
            .O(N__27030),
            .I(N__27018));
    InMux I__5215 (
            .O(N__27029),
            .I(N__27015));
    CascadeMux I__5214 (
            .O(N__27028),
            .I(N__27012));
    CascadeMux I__5213 (
            .O(N__27027),
            .I(N__27008));
    CascadeMux I__5212 (
            .O(N__27026),
            .I(N__27005));
    LocalMux I__5211 (
            .O(N__27021),
            .I(N__27002));
    LocalMux I__5210 (
            .O(N__27018),
            .I(N__26997));
    LocalMux I__5209 (
            .O(N__27015),
            .I(N__26997));
    InMux I__5208 (
            .O(N__27012),
            .I(N__26990));
    InMux I__5207 (
            .O(N__27011),
            .I(N__26990));
    InMux I__5206 (
            .O(N__27008),
            .I(N__26990));
    InMux I__5205 (
            .O(N__27005),
            .I(N__26987));
    Span4Mux_h I__5204 (
            .O(N__27002),
            .I(N__26984));
    Odrv4 I__5203 (
            .O(N__26997),
            .I(aluOperand1_fast_2));
    LocalMux I__5202 (
            .O(N__26990),
            .I(aluOperand1_fast_2));
    LocalMux I__5201 (
            .O(N__26987),
            .I(aluOperand1_fast_2));
    Odrv4 I__5200 (
            .O(N__26984),
            .I(aluOperand1_fast_2));
    InMux I__5199 (
            .O(N__26975),
            .I(N__26972));
    LocalMux I__5198 (
            .O(N__26972),
            .I(N__26969));
    Span4Mux_h I__5197 (
            .O(N__26969),
            .I(N__26966));
    Odrv4 I__5196 (
            .O(N__26966),
            .I(\ALU.dout_3_ns_1_4 ));
    InMux I__5195 (
            .O(N__26963),
            .I(N__26960));
    LocalMux I__5194 (
            .O(N__26960),
            .I(N__26956));
    InMux I__5193 (
            .O(N__26959),
            .I(N__26953));
    Span4Mux_h I__5192 (
            .O(N__26956),
            .I(N__26950));
    LocalMux I__5191 (
            .O(N__26953),
            .I(\ALU.eZ0Z_4 ));
    Odrv4 I__5190 (
            .O(N__26950),
            .I(\ALU.eZ0Z_4 ));
    InMux I__5189 (
            .O(N__26945),
            .I(N__26942));
    LocalMux I__5188 (
            .O(N__26942),
            .I(N__26939));
    Span4Mux_h I__5187 (
            .O(N__26939),
            .I(N__26936));
    Odrv4 I__5186 (
            .O(N__26936),
            .I(\ALU.e_RNIS97JZ0Z_1 ));
    InMux I__5185 (
            .O(N__26933),
            .I(N__26929));
    InMux I__5184 (
            .O(N__26932),
            .I(N__26926));
    LocalMux I__5183 (
            .O(N__26929),
            .I(N__26923));
    LocalMux I__5182 (
            .O(N__26926),
            .I(\ALU.eZ0Z_1 ));
    Odrv4 I__5181 (
            .O(N__26923),
            .I(\ALU.eZ0Z_1 ));
    InMux I__5180 (
            .O(N__26918),
            .I(N__26915));
    LocalMux I__5179 (
            .O(N__26915),
            .I(\ALU.N_701 ));
    InMux I__5178 (
            .O(N__26912),
            .I(N__26909));
    LocalMux I__5177 (
            .O(N__26909),
            .I(\ALU.dout_3_ns_1_2 ));
    InMux I__5176 (
            .O(N__26906),
            .I(N__26903));
    LocalMux I__5175 (
            .O(N__26903),
            .I(N__26900));
    Odrv12 I__5174 (
            .O(N__26900),
            .I(\ALU.dout_6_ns_1_7 ));
    InMux I__5173 (
            .O(N__26897),
            .I(N__26894));
    LocalMux I__5172 (
            .O(N__26894),
            .I(N__26891));
    Span4Mux_h I__5171 (
            .O(N__26891),
            .I(N__26888));
    Span4Mux_h I__5170 (
            .O(N__26888),
            .I(N__26885));
    Odrv4 I__5169 (
            .O(N__26885),
            .I(\ALU.f_RNIQQJ01Z0Z_7 ));
    InMux I__5168 (
            .O(N__26882),
            .I(N__26874));
    InMux I__5167 (
            .O(N__26881),
            .I(N__26874));
    InMux I__5166 (
            .O(N__26880),
            .I(N__26869));
    InMux I__5165 (
            .O(N__26879),
            .I(N__26869));
    LocalMux I__5164 (
            .O(N__26874),
            .I(N__26866));
    LocalMux I__5163 (
            .O(N__26869),
            .I(N__26863));
    Span4Mux_h I__5162 (
            .O(N__26866),
            .I(N__26860));
    Span4Mux_h I__5161 (
            .O(N__26863),
            .I(N__26857));
    Span4Mux_h I__5160 (
            .O(N__26860),
            .I(N__26854));
    Sp12to4 I__5159 (
            .O(N__26857),
            .I(N__26851));
    Span4Mux_v I__5158 (
            .O(N__26854),
            .I(N__26848));
    Span12Mux_v I__5157 (
            .O(N__26851),
            .I(N__26845));
    Span4Mux_v I__5156 (
            .O(N__26848),
            .I(N__26841));
    Span12Mux_h I__5155 (
            .O(N__26845),
            .I(N__26838));
    InMux I__5154 (
            .O(N__26844),
            .I(N__26835));
    Odrv4 I__5153 (
            .O(N__26841),
            .I(testWordZ0Z_8));
    Odrv12 I__5152 (
            .O(N__26838),
            .I(testWordZ0Z_8));
    LocalMux I__5151 (
            .O(N__26835),
            .I(testWordZ0Z_8));
    InMux I__5150 (
            .O(N__26828),
            .I(N__26823));
    InMux I__5149 (
            .O(N__26827),
            .I(N__26820));
    InMux I__5148 (
            .O(N__26826),
            .I(N__26817));
    LocalMux I__5147 (
            .O(N__26823),
            .I(N__26812));
    LocalMux I__5146 (
            .O(N__26820),
            .I(N__26812));
    LocalMux I__5145 (
            .O(N__26817),
            .I(N__26809));
    Span4Mux_v I__5144 (
            .O(N__26812),
            .I(N__26806));
    Odrv12 I__5143 (
            .O(N__26809),
            .I(\ALU.fZ0Z_10 ));
    Odrv4 I__5142 (
            .O(N__26806),
            .I(\ALU.fZ0Z_10 ));
    InMux I__5141 (
            .O(N__26801),
            .I(N__26798));
    LocalMux I__5140 (
            .O(N__26798),
            .I(N__26795));
    Span4Mux_h I__5139 (
            .O(N__26795),
            .I(N__26792));
    Span4Mux_h I__5138 (
            .O(N__26792),
            .I(N__26789));
    Odrv4 I__5137 (
            .O(N__26789),
            .I(\ALU.b_RNIEHSD1Z0Z_10 ));
    InMux I__5136 (
            .O(N__26786),
            .I(N__26783));
    LocalMux I__5135 (
            .O(N__26783),
            .I(N__26780));
    Span4Mux_v I__5134 (
            .O(N__26780),
            .I(N__26777));
    Span4Mux_h I__5133 (
            .O(N__26777),
            .I(N__26774));
    Odrv4 I__5132 (
            .O(N__26774),
            .I(\ALU.madd_cry_13_ma ));
    CascadeMux I__5131 (
            .O(N__26771),
            .I(N__26768));
    InMux I__5130 (
            .O(N__26768),
            .I(N__26765));
    LocalMux I__5129 (
            .O(N__26765),
            .I(N__26762));
    Span4Mux_h I__5128 (
            .O(N__26762),
            .I(N__26759));
    Span4Mux_h I__5127 (
            .O(N__26759),
            .I(N__26756));
    Odrv4 I__5126 (
            .O(N__26756),
            .I(\ALU.madd_axb_13_l_ofx ));
    InMux I__5125 (
            .O(N__26753),
            .I(\ALU.madd_cry_12 ));
    InMux I__5124 (
            .O(N__26750),
            .I(N__26747));
    LocalMux I__5123 (
            .O(N__26747),
            .I(N__26744));
    Span4Mux_h I__5122 (
            .O(N__26744),
            .I(N__26741));
    Span4Mux_h I__5121 (
            .O(N__26741),
            .I(N__26738));
    Odrv4 I__5120 (
            .O(N__26738),
            .I(\ALU.madd_axb_14 ));
    InMux I__5119 (
            .O(N__26735),
            .I(\ALU.madd_cry_13 ));
    InMux I__5118 (
            .O(N__26732),
            .I(N__26722));
    InMux I__5117 (
            .O(N__26731),
            .I(N__26722));
    InMux I__5116 (
            .O(N__26730),
            .I(N__26717));
    InMux I__5115 (
            .O(N__26729),
            .I(N__26717));
    InMux I__5114 (
            .O(N__26728),
            .I(N__26712));
    InMux I__5113 (
            .O(N__26727),
            .I(N__26708));
    LocalMux I__5112 (
            .O(N__26722),
            .I(N__26705));
    LocalMux I__5111 (
            .O(N__26717),
            .I(N__26702));
    InMux I__5110 (
            .O(N__26716),
            .I(N__26697));
    InMux I__5109 (
            .O(N__26715),
            .I(N__26697));
    LocalMux I__5108 (
            .O(N__26712),
            .I(N__26694));
    InMux I__5107 (
            .O(N__26711),
            .I(N__26691));
    LocalMux I__5106 (
            .O(N__26708),
            .I(N__26686));
    Span4Mux_h I__5105 (
            .O(N__26705),
            .I(N__26683));
    Span4Mux_v I__5104 (
            .O(N__26702),
            .I(N__26678));
    LocalMux I__5103 (
            .O(N__26697),
            .I(N__26678));
    Span4Mux_v I__5102 (
            .O(N__26694),
            .I(N__26673));
    LocalMux I__5101 (
            .O(N__26691),
            .I(N__26673));
    InMux I__5100 (
            .O(N__26690),
            .I(N__26668));
    InMux I__5099 (
            .O(N__26689),
            .I(N__26668));
    Span12Mux_s6_h I__5098 (
            .O(N__26686),
            .I(N__26665));
    Span4Mux_v I__5097 (
            .O(N__26683),
            .I(N__26660));
    Span4Mux_h I__5096 (
            .O(N__26678),
            .I(N__26660));
    Odrv4 I__5095 (
            .O(N__26673),
            .I(\ALU.operand2_6 ));
    LocalMux I__5094 (
            .O(N__26668),
            .I(\ALU.operand2_6 ));
    Odrv12 I__5093 (
            .O(N__26665),
            .I(\ALU.operand2_6 ));
    Odrv4 I__5092 (
            .O(N__26660),
            .I(\ALU.operand2_6 ));
    CascadeMux I__5091 (
            .O(N__26651),
            .I(N__26646));
    InMux I__5090 (
            .O(N__26650),
            .I(N__26643));
    InMux I__5089 (
            .O(N__26649),
            .I(N__26638));
    InMux I__5088 (
            .O(N__26646),
            .I(N__26634));
    LocalMux I__5087 (
            .O(N__26643),
            .I(N__26631));
    CascadeMux I__5086 (
            .O(N__26642),
            .I(N__26628));
    CascadeMux I__5085 (
            .O(N__26641),
            .I(N__26623));
    LocalMux I__5084 (
            .O(N__26638),
            .I(N__26620));
    InMux I__5083 (
            .O(N__26637),
            .I(N__26617));
    LocalMux I__5082 (
            .O(N__26634),
            .I(N__26612));
    Span4Mux_h I__5081 (
            .O(N__26631),
            .I(N__26612));
    InMux I__5080 (
            .O(N__26628),
            .I(N__26609));
    CascadeMux I__5079 (
            .O(N__26627),
            .I(N__26606));
    CascadeMux I__5078 (
            .O(N__26626),
            .I(N__26592));
    InMux I__5077 (
            .O(N__26623),
            .I(N__26589));
    Span4Mux_s1_v I__5076 (
            .O(N__26620),
            .I(N__26583));
    LocalMux I__5075 (
            .O(N__26617),
            .I(N__26583));
    Span4Mux_h I__5074 (
            .O(N__26612),
            .I(N__26578));
    LocalMux I__5073 (
            .O(N__26609),
            .I(N__26578));
    InMux I__5072 (
            .O(N__26606),
            .I(N__26572));
    InMux I__5071 (
            .O(N__26605),
            .I(N__26569));
    CascadeMux I__5070 (
            .O(N__26604),
            .I(N__26565));
    CascadeMux I__5069 (
            .O(N__26603),
            .I(N__26561));
    CascadeMux I__5068 (
            .O(N__26602),
            .I(N__26558));
    CascadeMux I__5067 (
            .O(N__26601),
            .I(N__26555));
    CascadeMux I__5066 (
            .O(N__26600),
            .I(N__26550));
    CascadeMux I__5065 (
            .O(N__26599),
            .I(N__26546));
    CascadeMux I__5064 (
            .O(N__26598),
            .I(N__26543));
    CascadeMux I__5063 (
            .O(N__26597),
            .I(N__26540));
    CascadeMux I__5062 (
            .O(N__26596),
            .I(N__26537));
    InMux I__5061 (
            .O(N__26595),
            .I(N__26530));
    InMux I__5060 (
            .O(N__26592),
            .I(N__26530));
    LocalMux I__5059 (
            .O(N__26589),
            .I(N__26527));
    CascadeMux I__5058 (
            .O(N__26588),
            .I(N__26524));
    Span4Mux_v I__5057 (
            .O(N__26583),
            .I(N__26518));
    Span4Mux_v I__5056 (
            .O(N__26578),
            .I(N__26518));
    CascadeMux I__5055 (
            .O(N__26577),
            .I(N__26515));
    CascadeMux I__5054 (
            .O(N__26576),
            .I(N__26511));
    InMux I__5053 (
            .O(N__26575),
            .I(N__26508));
    LocalMux I__5052 (
            .O(N__26572),
            .I(N__26503));
    LocalMux I__5051 (
            .O(N__26569),
            .I(N__26503));
    InMux I__5050 (
            .O(N__26568),
            .I(N__26500));
    InMux I__5049 (
            .O(N__26565),
            .I(N__26487));
    InMux I__5048 (
            .O(N__26564),
            .I(N__26487));
    InMux I__5047 (
            .O(N__26561),
            .I(N__26487));
    InMux I__5046 (
            .O(N__26558),
            .I(N__26484));
    InMux I__5045 (
            .O(N__26555),
            .I(N__26477));
    InMux I__5044 (
            .O(N__26554),
            .I(N__26477));
    InMux I__5043 (
            .O(N__26553),
            .I(N__26477));
    InMux I__5042 (
            .O(N__26550),
            .I(N__26468));
    InMux I__5041 (
            .O(N__26549),
            .I(N__26468));
    InMux I__5040 (
            .O(N__26546),
            .I(N__26468));
    InMux I__5039 (
            .O(N__26543),
            .I(N__26468));
    InMux I__5038 (
            .O(N__26540),
            .I(N__26463));
    InMux I__5037 (
            .O(N__26537),
            .I(N__26463));
    CascadeMux I__5036 (
            .O(N__26536),
            .I(N__26460));
    CascadeMux I__5035 (
            .O(N__26535),
            .I(N__26457));
    LocalMux I__5034 (
            .O(N__26530),
            .I(N__26452));
    Span4Mux_v I__5033 (
            .O(N__26527),
            .I(N__26452));
    InMux I__5032 (
            .O(N__26524),
            .I(N__26449));
    InMux I__5031 (
            .O(N__26523),
            .I(N__26446));
    Span4Mux_h I__5030 (
            .O(N__26518),
            .I(N__26442));
    InMux I__5029 (
            .O(N__26515),
            .I(N__26439));
    InMux I__5028 (
            .O(N__26514),
            .I(N__26436));
    InMux I__5027 (
            .O(N__26511),
            .I(N__26433));
    LocalMux I__5026 (
            .O(N__26508),
            .I(N__26428));
    Span4Mux_h I__5025 (
            .O(N__26503),
            .I(N__26428));
    LocalMux I__5024 (
            .O(N__26500),
            .I(N__26425));
    InMux I__5023 (
            .O(N__26499),
            .I(N__26418));
    InMux I__5022 (
            .O(N__26498),
            .I(N__26418));
    InMux I__5021 (
            .O(N__26497),
            .I(N__26418));
    CascadeMux I__5020 (
            .O(N__26496),
            .I(N__26415));
    CascadeMux I__5019 (
            .O(N__26495),
            .I(N__26412));
    CascadeMux I__5018 (
            .O(N__26494),
            .I(N__26409));
    LocalMux I__5017 (
            .O(N__26487),
            .I(N__26404));
    LocalMux I__5016 (
            .O(N__26484),
            .I(N__26404));
    LocalMux I__5015 (
            .O(N__26477),
            .I(N__26401));
    LocalMux I__5014 (
            .O(N__26468),
            .I(N__26398));
    LocalMux I__5013 (
            .O(N__26463),
            .I(N__26395));
    InMux I__5012 (
            .O(N__26460),
            .I(N__26390));
    InMux I__5011 (
            .O(N__26457),
            .I(N__26390));
    Span4Mux_h I__5010 (
            .O(N__26452),
            .I(N__26387));
    LocalMux I__5009 (
            .O(N__26449),
            .I(N__26384));
    LocalMux I__5008 (
            .O(N__26446),
            .I(N__26381));
    CascadeMux I__5007 (
            .O(N__26445),
            .I(N__26376));
    Span4Mux_v I__5006 (
            .O(N__26442),
            .I(N__26370));
    LocalMux I__5005 (
            .O(N__26439),
            .I(N__26370));
    LocalMux I__5004 (
            .O(N__26436),
            .I(N__26363));
    LocalMux I__5003 (
            .O(N__26433),
            .I(N__26363));
    Span4Mux_v I__5002 (
            .O(N__26428),
            .I(N__26363));
    Span4Mux_s1_h I__5001 (
            .O(N__26425),
            .I(N__26358));
    LocalMux I__5000 (
            .O(N__26418),
            .I(N__26358));
    InMux I__4999 (
            .O(N__26415),
            .I(N__26355));
    InMux I__4998 (
            .O(N__26412),
            .I(N__26352));
    InMux I__4997 (
            .O(N__26409),
            .I(N__26349));
    Sp12to4 I__4996 (
            .O(N__26404),
            .I(N__26346));
    Span4Mux_h I__4995 (
            .O(N__26401),
            .I(N__26341));
    Span4Mux_v I__4994 (
            .O(N__26398),
            .I(N__26341));
    Span4Mux_h I__4993 (
            .O(N__26395),
            .I(N__26334));
    LocalMux I__4992 (
            .O(N__26390),
            .I(N__26334));
    Span4Mux_v I__4991 (
            .O(N__26387),
            .I(N__26334));
    Span4Mux_v I__4990 (
            .O(N__26384),
            .I(N__26329));
    Span4Mux_h I__4989 (
            .O(N__26381),
            .I(N__26329));
    InMux I__4988 (
            .O(N__26380),
            .I(N__26320));
    InMux I__4987 (
            .O(N__26379),
            .I(N__26320));
    InMux I__4986 (
            .O(N__26376),
            .I(N__26320));
    InMux I__4985 (
            .O(N__26375),
            .I(N__26320));
    Span4Mux_h I__4984 (
            .O(N__26370),
            .I(N__26317));
    Span4Mux_v I__4983 (
            .O(N__26363),
            .I(N__26314));
    Sp12to4 I__4982 (
            .O(N__26358),
            .I(N__26303));
    LocalMux I__4981 (
            .O(N__26355),
            .I(N__26303));
    LocalMux I__4980 (
            .O(N__26352),
            .I(N__26303));
    LocalMux I__4979 (
            .O(N__26349),
            .I(N__26303));
    Span12Mux_h I__4978 (
            .O(N__26346),
            .I(N__26303));
    Span4Mux_h I__4977 (
            .O(N__26341),
            .I(N__26298));
    Span4Mux_v I__4976 (
            .O(N__26334),
            .I(N__26298));
    Odrv4 I__4975 (
            .O(N__26329),
            .I(aluReadBus));
    LocalMux I__4974 (
            .O(N__26320),
            .I(aluReadBus));
    Odrv4 I__4973 (
            .O(N__26317),
            .I(aluReadBus));
    Odrv4 I__4972 (
            .O(N__26314),
            .I(aluReadBus));
    Odrv12 I__4971 (
            .O(N__26303),
            .I(aluReadBus));
    Odrv4 I__4970 (
            .O(N__26298),
            .I(aluReadBus));
    InMux I__4969 (
            .O(N__26285),
            .I(N__26271));
    InMux I__4968 (
            .O(N__26284),
            .I(N__26271));
    InMux I__4967 (
            .O(N__26283),
            .I(N__26268));
    InMux I__4966 (
            .O(N__26282),
            .I(N__26265));
    InMux I__4965 (
            .O(N__26281),
            .I(N__26262));
    InMux I__4964 (
            .O(N__26280),
            .I(N__26259));
    InMux I__4963 (
            .O(N__26279),
            .I(N__26254));
    InMux I__4962 (
            .O(N__26278),
            .I(N__26254));
    InMux I__4961 (
            .O(N__26277),
            .I(N__26248));
    InMux I__4960 (
            .O(N__26276),
            .I(N__26248));
    LocalMux I__4959 (
            .O(N__26271),
            .I(N__26245));
    LocalMux I__4958 (
            .O(N__26268),
            .I(N__26242));
    LocalMux I__4957 (
            .O(N__26265),
            .I(N__26237));
    LocalMux I__4956 (
            .O(N__26262),
            .I(N__26237));
    LocalMux I__4955 (
            .O(N__26259),
            .I(N__26232));
    LocalMux I__4954 (
            .O(N__26254),
            .I(N__26232));
    InMux I__4953 (
            .O(N__26253),
            .I(N__26229));
    LocalMux I__4952 (
            .O(N__26248),
            .I(N__26226));
    Span4Mux_h I__4951 (
            .O(N__26245),
            .I(N__26223));
    Span4Mux_h I__4950 (
            .O(N__26242),
            .I(N__26220));
    Span4Mux_v I__4949 (
            .O(N__26237),
            .I(N__26215));
    Span4Mux_h I__4948 (
            .O(N__26232),
            .I(N__26215));
    LocalMux I__4947 (
            .O(N__26229),
            .I(N__26212));
    Span4Mux_h I__4946 (
            .O(N__26226),
            .I(N__26209));
    Span4Mux_s0_h I__4945 (
            .O(N__26223),
            .I(N__26206));
    Span4Mux_v I__4944 (
            .O(N__26220),
            .I(N__26201));
    Span4Mux_h I__4943 (
            .O(N__26215),
            .I(N__26201));
    Odrv12 I__4942 (
            .O(N__26212),
            .I(\ALU.N_217_0 ));
    Odrv4 I__4941 (
            .O(N__26209),
            .I(\ALU.N_217_0 ));
    Odrv4 I__4940 (
            .O(N__26206),
            .I(\ALU.N_217_0 ));
    Odrv4 I__4939 (
            .O(N__26201),
            .I(\ALU.N_217_0 ));
    CascadeMux I__4938 (
            .O(N__26192),
            .I(\ALU.dout_3_ns_1_15_cascade_ ));
    CascadeMux I__4937 (
            .O(N__26189),
            .I(\ALU.dout_6_ns_1_2_cascade_ ));
    CascadeMux I__4936 (
            .O(N__26186),
            .I(\ALU.N_749_cascade_ ));
    InMux I__4935 (
            .O(N__26183),
            .I(N__26180));
    LocalMux I__4934 (
            .O(N__26180),
            .I(N__26176));
    InMux I__4933 (
            .O(N__26179),
            .I(N__26173));
    Span4Mux_v I__4932 (
            .O(N__26176),
            .I(N__26170));
    LocalMux I__4931 (
            .O(N__26173),
            .I(N__26167));
    Sp12to4 I__4930 (
            .O(N__26170),
            .I(N__26162));
    Span12Mux_h I__4929 (
            .O(N__26167),
            .I(N__26162));
    Odrv12 I__4928 (
            .O(N__26162),
            .I(\ALU.madd_52 ));
    CascadeMux I__4927 (
            .O(N__26159),
            .I(N__26156));
    InMux I__4926 (
            .O(N__26156),
            .I(N__26153));
    LocalMux I__4925 (
            .O(N__26153),
            .I(N__26150));
    Span4Mux_v I__4924 (
            .O(N__26150),
            .I(N__26147));
    Span4Mux_h I__4923 (
            .O(N__26147),
            .I(N__26144));
    Span4Mux_v I__4922 (
            .O(N__26144),
            .I(N__26141));
    Odrv4 I__4921 (
            .O(N__26141),
            .I(\ALU.madd_axb_5_l_fx ));
    InMux I__4920 (
            .O(N__26138),
            .I(\ALU.madd_cry_4 ));
    InMux I__4919 (
            .O(N__26135),
            .I(\ALU.madd_cry_5 ));
    InMux I__4918 (
            .O(N__26132),
            .I(N__26129));
    LocalMux I__4917 (
            .O(N__26129),
            .I(N__26125));
    InMux I__4916 (
            .O(N__26128),
            .I(N__26122));
    Span4Mux_v I__4915 (
            .O(N__26125),
            .I(N__26117));
    LocalMux I__4914 (
            .O(N__26122),
            .I(N__26117));
    Span4Mux_v I__4913 (
            .O(N__26117),
            .I(N__26114));
    Span4Mux_h I__4912 (
            .O(N__26114),
            .I(N__26111));
    Odrv4 I__4911 (
            .O(N__26111),
            .I(\ALU.madd_axb_7 ));
    InMux I__4910 (
            .O(N__26108),
            .I(N__26105));
    LocalMux I__4909 (
            .O(N__26105),
            .I(N__26102));
    Odrv4 I__4908 (
            .O(N__26102),
            .I(\ALU.madd_cry_6_THRU_CO ));
    InMux I__4907 (
            .O(N__26099),
            .I(\ALU.madd_cry_6 ));
    InMux I__4906 (
            .O(N__26096),
            .I(N__26093));
    LocalMux I__4905 (
            .O(N__26093),
            .I(N__26090));
    Span4Mux_h I__4904 (
            .O(N__26090),
            .I(N__26087));
    Span4Mux_h I__4903 (
            .O(N__26087),
            .I(N__26084));
    Span4Mux_v I__4902 (
            .O(N__26084),
            .I(N__26081));
    Odrv4 I__4901 (
            .O(N__26081),
            .I(\ALU.madd_axb_8_l_fx ));
    CascadeMux I__4900 (
            .O(N__26078),
            .I(N__26075));
    InMux I__4899 (
            .O(N__26075),
            .I(N__26072));
    LocalMux I__4898 (
            .O(N__26072),
            .I(N__26069));
    Span4Mux_v I__4897 (
            .O(N__26069),
            .I(N__26065));
    InMux I__4896 (
            .O(N__26068),
            .I(N__26062));
    Span4Mux_h I__4895 (
            .O(N__26065),
            .I(N__26059));
    LocalMux I__4894 (
            .O(N__26062),
            .I(\ALU.madd_159 ));
    Odrv4 I__4893 (
            .O(N__26059),
            .I(\ALU.madd_159 ));
    InMux I__4892 (
            .O(N__26054),
            .I(bfn_9_10_0_));
    InMux I__4891 (
            .O(N__26051),
            .I(N__26048));
    LocalMux I__4890 (
            .O(N__26048),
            .I(N__26045));
    Span12Mux_h I__4889 (
            .O(N__26045),
            .I(N__26042));
    Odrv12 I__4888 (
            .O(N__26042),
            .I(\ALU.madd_cry_9_ma ));
    CascadeMux I__4887 (
            .O(N__26039),
            .I(N__26036));
    InMux I__4886 (
            .O(N__26036),
            .I(N__26033));
    LocalMux I__4885 (
            .O(N__26033),
            .I(N__26030));
    Span4Mux_h I__4884 (
            .O(N__26030),
            .I(N__26027));
    Span4Mux_v I__4883 (
            .O(N__26027),
            .I(N__26024));
    Span4Mux_h I__4882 (
            .O(N__26024),
            .I(N__26021));
    Odrv4 I__4881 (
            .O(N__26021),
            .I(\ALU.madd_axb_9_l_ofx ));
    InMux I__4880 (
            .O(N__26018),
            .I(\ALU.madd_cry_8 ));
    InMux I__4879 (
            .O(N__26015),
            .I(N__26012));
    LocalMux I__4878 (
            .O(N__26012),
            .I(N__26009));
    Span4Mux_h I__4877 (
            .O(N__26009),
            .I(N__26006));
    Span4Mux_h I__4876 (
            .O(N__26006),
            .I(N__26003));
    Span4Mux_h I__4875 (
            .O(N__26003),
            .I(N__26000));
    Odrv4 I__4874 (
            .O(N__26000),
            .I(\ALU.madd_cry_10_ma ));
    CascadeMux I__4873 (
            .O(N__25997),
            .I(N__25994));
    InMux I__4872 (
            .O(N__25994),
            .I(N__25991));
    LocalMux I__4871 (
            .O(N__25991),
            .I(N__25988));
    Span12Mux_h I__4870 (
            .O(N__25988),
            .I(N__25985));
    Odrv12 I__4869 (
            .O(N__25985),
            .I(\ALU.madd_axb_10_l_ofx ));
    InMux I__4868 (
            .O(N__25982),
            .I(\ALU.madd_cry_9 ));
    CascadeMux I__4867 (
            .O(N__25979),
            .I(N__25976));
    InMux I__4866 (
            .O(N__25976),
            .I(N__25973));
    LocalMux I__4865 (
            .O(N__25973),
            .I(N__25970));
    Span12Mux_h I__4864 (
            .O(N__25970),
            .I(N__25967));
    Odrv12 I__4863 (
            .O(N__25967),
            .I(\ALU.madd_axb_11 ));
    InMux I__4862 (
            .O(N__25964),
            .I(\ALU.madd_cry_10 ));
    InMux I__4861 (
            .O(N__25961),
            .I(N__25958));
    LocalMux I__4860 (
            .O(N__25958),
            .I(N__25955));
    Span4Mux_h I__4859 (
            .O(N__25955),
            .I(N__25952));
    Span4Mux_h I__4858 (
            .O(N__25952),
            .I(N__25949));
    Span4Mux_s1_h I__4857 (
            .O(N__25949),
            .I(N__25946));
    Odrv4 I__4856 (
            .O(N__25946),
            .I(\ALU.madd_axb_12_l_fx ));
    CascadeMux I__4855 (
            .O(N__25943),
            .I(N__25940));
    InMux I__4854 (
            .O(N__25940),
            .I(N__25937));
    LocalMux I__4853 (
            .O(N__25937),
            .I(N__25934));
    Span4Mux_v I__4852 (
            .O(N__25934),
            .I(N__25930));
    InMux I__4851 (
            .O(N__25933),
            .I(N__25927));
    Span4Mux_h I__4850 (
            .O(N__25930),
            .I(N__25924));
    LocalMux I__4849 (
            .O(N__25927),
            .I(\ALU.madd_360 ));
    Odrv4 I__4848 (
            .O(N__25924),
            .I(\ALU.madd_360 ));
    InMux I__4847 (
            .O(N__25919),
            .I(\ALU.madd_cry_11 ));
    CascadeMux I__4846 (
            .O(N__25916),
            .I(N__25913));
    InMux I__4845 (
            .O(N__25913),
            .I(N__25909));
    InMux I__4844 (
            .O(N__25912),
            .I(N__25906));
    LocalMux I__4843 (
            .O(N__25909),
            .I(N__25901));
    LocalMux I__4842 (
            .O(N__25906),
            .I(N__25901));
    Span4Mux_v I__4841 (
            .O(N__25901),
            .I(N__25898));
    Span4Mux_v I__4840 (
            .O(N__25898),
            .I(N__25895));
    Odrv4 I__4839 (
            .O(N__25895),
            .I(\ALU.fZ0Z_15 ));
    InMux I__4838 (
            .O(N__25892),
            .I(N__25889));
    LocalMux I__4837 (
            .O(N__25889),
            .I(N__25886));
    Span4Mux_h I__4836 (
            .O(N__25886),
            .I(N__25883));
    Span4Mux_v I__4835 (
            .O(N__25883),
            .I(N__25880));
    Odrv4 I__4834 (
            .O(N__25880),
            .I(\ALU.madd_cry_0_ma ));
    CascadeMux I__4833 (
            .O(N__25877),
            .I(N__25874));
    InMux I__4832 (
            .O(N__25874),
            .I(N__25871));
    LocalMux I__4831 (
            .O(N__25871),
            .I(N__25868));
    Span4Mux_h I__4830 (
            .O(N__25868),
            .I(N__25865));
    Span4Mux_h I__4829 (
            .O(N__25865),
            .I(N__25862));
    Span4Mux_v I__4828 (
            .O(N__25862),
            .I(N__25859));
    Odrv4 I__4827 (
            .O(N__25859),
            .I(\ALU.madd_cry_1_ma ));
    InMux I__4826 (
            .O(N__25856),
            .I(\ALU.madd_cry_0 ));
    InMux I__4825 (
            .O(N__25853),
            .I(N__25850));
    LocalMux I__4824 (
            .O(N__25850),
            .I(N__25847));
    Span4Mux_h I__4823 (
            .O(N__25847),
            .I(N__25844));
    Span4Mux_v I__4822 (
            .O(N__25844),
            .I(N__25841));
    Odrv4 I__4821 (
            .O(N__25841),
            .I(\ALU.madd_axb_2_l_fx ));
    CascadeMux I__4820 (
            .O(N__25838),
            .I(N__25835));
    InMux I__4819 (
            .O(N__25835),
            .I(N__25832));
    LocalMux I__4818 (
            .O(N__25832),
            .I(N__25828));
    CascadeMux I__4817 (
            .O(N__25831),
            .I(N__25825));
    Span4Mux_v I__4816 (
            .O(N__25828),
            .I(N__25822));
    InMux I__4815 (
            .O(N__25825),
            .I(N__25819));
    Span4Mux_v I__4814 (
            .O(N__25822),
            .I(N__25816));
    LocalMux I__4813 (
            .O(N__25819),
            .I(N__25813));
    Span4Mux_v I__4812 (
            .O(N__25816),
            .I(N__25810));
    Span4Mux_v I__4811 (
            .O(N__25813),
            .I(N__25807));
    Sp12to4 I__4810 (
            .O(N__25810),
            .I(N__25804));
    Span4Mux_h I__4809 (
            .O(N__25807),
            .I(N__25801));
    Odrv12 I__4808 (
            .O(N__25804),
            .I(\ALU.madd_6 ));
    Odrv4 I__4807 (
            .O(N__25801),
            .I(\ALU.madd_6 ));
    InMux I__4806 (
            .O(N__25796),
            .I(\ALU.madd_cry_1 ));
    InMux I__4805 (
            .O(N__25793),
            .I(N__25790));
    LocalMux I__4804 (
            .O(N__25790),
            .I(N__25787));
    Span4Mux_h I__4803 (
            .O(N__25787),
            .I(N__25784));
    Odrv4 I__4802 (
            .O(N__25784),
            .I(\ALU.madd_13 ));
    CascadeMux I__4801 (
            .O(N__25781),
            .I(N__25778));
    InMux I__4800 (
            .O(N__25778),
            .I(N__25775));
    LocalMux I__4799 (
            .O(N__25775),
            .I(N__25772));
    Span4Mux_v I__4798 (
            .O(N__25772),
            .I(N__25769));
    Span4Mux_v I__4797 (
            .O(N__25769),
            .I(N__25766));
    Span4Mux_h I__4796 (
            .O(N__25766),
            .I(N__25763));
    Odrv4 I__4795 (
            .O(N__25763),
            .I(\ALU.madd_18 ));
    InMux I__4794 (
            .O(N__25760),
            .I(\ALU.madd_cry_2 ));
    InMux I__4793 (
            .O(N__25757),
            .I(N__25754));
    LocalMux I__4792 (
            .O(N__25754),
            .I(N__25751));
    Span4Mux_h I__4791 (
            .O(N__25751),
            .I(N__25748));
    Span4Mux_h I__4790 (
            .O(N__25748),
            .I(N__25745));
    Odrv4 I__4789 (
            .O(N__25745),
            .I(\ALU.madd_axb_4_l_fx ));
    CascadeMux I__4788 (
            .O(N__25742),
            .I(N__25738));
    InMux I__4787 (
            .O(N__25741),
            .I(N__25735));
    InMux I__4786 (
            .O(N__25738),
            .I(N__25732));
    LocalMux I__4785 (
            .O(N__25735),
            .I(N__25729));
    LocalMux I__4784 (
            .O(N__25732),
            .I(N__25726));
    Span4Mux_h I__4783 (
            .O(N__25729),
            .I(N__25721));
    Span4Mux_v I__4782 (
            .O(N__25726),
            .I(N__25721));
    Span4Mux_h I__4781 (
            .O(N__25721),
            .I(N__25718));
    Odrv4 I__4780 (
            .O(N__25718),
            .I(\ALU.madd_30 ));
    InMux I__4779 (
            .O(N__25715),
            .I(\ALU.madd_cry_3 ));
    InMux I__4778 (
            .O(N__25712),
            .I(N__25709));
    LocalMux I__4777 (
            .O(N__25709),
            .I(N__25706));
    Span4Mux_h I__4776 (
            .O(N__25706),
            .I(N__25703));
    Span4Mux_h I__4775 (
            .O(N__25703),
            .I(N__25700));
    Odrv4 I__4774 (
            .O(N__25700),
            .I(\ALU.d_RNICJE9BZ0Z_8 ));
    InMux I__4773 (
            .O(N__25697),
            .I(N__25694));
    LocalMux I__4772 (
            .O(N__25694),
            .I(N__25691));
    Span4Mux_h I__4771 (
            .O(N__25691),
            .I(N__25688));
    Odrv4 I__4770 (
            .O(N__25688),
            .I(\ALU.d_RNIEUKR11Z0Z_0 ));
    InMux I__4769 (
            .O(N__25685),
            .I(N__25682));
    LocalMux I__4768 (
            .O(N__25682),
            .I(N__25679));
    Span4Mux_v I__4767 (
            .O(N__25679),
            .I(N__25676));
    Span4Mux_h I__4766 (
            .O(N__25676),
            .I(N__25673));
    Span4Mux_h I__4765 (
            .O(N__25673),
            .I(N__25670));
    Odrv4 I__4764 (
            .O(N__25670),
            .I(\ALU.a_15_m3_8 ));
    CascadeMux I__4763 (
            .O(N__25667),
            .I(\ALU.a_15_m4_8_cascade_ ));
    InMux I__4762 (
            .O(N__25664),
            .I(N__25661));
    LocalMux I__4761 (
            .O(N__25661),
            .I(\ALU.a_15_m5_8 ));
    CascadeMux I__4760 (
            .O(N__25658),
            .I(N__25655));
    InMux I__4759 (
            .O(N__25655),
            .I(N__25651));
    CascadeMux I__4758 (
            .O(N__25654),
            .I(N__25648));
    LocalMux I__4757 (
            .O(N__25651),
            .I(N__25645));
    InMux I__4756 (
            .O(N__25648),
            .I(N__25642));
    Span4Mux_v I__4755 (
            .O(N__25645),
            .I(N__25639));
    LocalMux I__4754 (
            .O(N__25642),
            .I(N__25636));
    Span4Mux_h I__4753 (
            .O(N__25639),
            .I(N__25631));
    Span4Mux_v I__4752 (
            .O(N__25636),
            .I(N__25631));
    Odrv4 I__4751 (
            .O(N__25631),
            .I(\ALU.fZ0Z_8 ));
    InMux I__4750 (
            .O(N__25628),
            .I(N__25624));
    InMux I__4749 (
            .O(N__25627),
            .I(N__25621));
    LocalMux I__4748 (
            .O(N__25624),
            .I(N__25618));
    LocalMux I__4747 (
            .O(N__25621),
            .I(N__25615));
    Span12Mux_v I__4746 (
            .O(N__25618),
            .I(N__25612));
    Odrv12 I__4745 (
            .O(N__25615),
            .I(\ALU.dZ0Z_8 ));
    Odrv12 I__4744 (
            .O(N__25612),
            .I(\ALU.dZ0Z_8 ));
    CascadeMux I__4743 (
            .O(N__25607),
            .I(\ALU.operand2_6_ns_1_8_cascade_ ));
    InMux I__4742 (
            .O(N__25604),
            .I(N__25601));
    LocalMux I__4741 (
            .O(N__25601),
            .I(N__25598));
    Odrv12 I__4740 (
            .O(N__25598),
            .I(\ALU.N_867 ));
    InMux I__4739 (
            .O(N__25595),
            .I(N__25592));
    LocalMux I__4738 (
            .O(N__25592),
            .I(N__25589));
    Span4Mux_h I__4737 (
            .O(N__25589),
            .I(N__25586));
    Span4Mux_h I__4736 (
            .O(N__25586),
            .I(N__25582));
    InMux I__4735 (
            .O(N__25585),
            .I(N__25579));
    Odrv4 I__4734 (
            .O(N__25582),
            .I(\ALU.hZ0Z_8 ));
    LocalMux I__4733 (
            .O(N__25579),
            .I(\ALU.hZ0Z_8 ));
    CascadeMux I__4732 (
            .O(N__25574),
            .I(\ALU.N_186_0_i_cascade_ ));
    InMux I__4731 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__4730 (
            .O(N__25568),
            .I(N__25565));
    Span4Mux_v I__4729 (
            .O(N__25565),
            .I(N__25562));
    Span4Mux_h I__4728 (
            .O(N__25562),
            .I(N__25559));
    Odrv4 I__4727 (
            .O(N__25559),
            .I(\ALU.c_RNIA7OEEZ0Z_11 ));
    CascadeMux I__4726 (
            .O(N__25556),
            .I(N__25553));
    InMux I__4725 (
            .O(N__25553),
            .I(N__25550));
    LocalMux I__4724 (
            .O(N__25550),
            .I(N__25547));
    Span4Mux_v I__4723 (
            .O(N__25547),
            .I(N__25542));
    InMux I__4722 (
            .O(N__25546),
            .I(N__25539));
    CascadeMux I__4721 (
            .O(N__25545),
            .I(N__25535));
    Span4Mux_h I__4720 (
            .O(N__25542),
            .I(N__25531));
    LocalMux I__4719 (
            .O(N__25539),
            .I(N__25528));
    InMux I__4718 (
            .O(N__25538),
            .I(N__25525));
    InMux I__4717 (
            .O(N__25535),
            .I(N__25522));
    InMux I__4716 (
            .O(N__25534),
            .I(N__25519));
    Span4Mux_h I__4715 (
            .O(N__25531),
            .I(N__25516));
    Span4Mux_s1_v I__4714 (
            .O(N__25528),
            .I(N__25513));
    LocalMux I__4713 (
            .O(N__25525),
            .I(N__25506));
    LocalMux I__4712 (
            .O(N__25522),
            .I(N__25506));
    LocalMux I__4711 (
            .O(N__25519),
            .I(N__25506));
    Odrv4 I__4710 (
            .O(N__25516),
            .I(RXbuffer_5));
    Odrv4 I__4709 (
            .O(N__25513),
            .I(RXbuffer_5));
    Odrv12 I__4708 (
            .O(N__25506),
            .I(RXbuffer_5));
    InMux I__4707 (
            .O(N__25499),
            .I(N__25496));
    LocalMux I__4706 (
            .O(N__25496),
            .I(N__25493));
    Span4Mux_h I__4705 (
            .O(N__25493),
            .I(N__25489));
    InMux I__4704 (
            .O(N__25492),
            .I(N__25486));
    Odrv4 I__4703 (
            .O(N__25489),
            .I(\ALU.hZ0Z_12 ));
    LocalMux I__4702 (
            .O(N__25486),
            .I(\ALU.hZ0Z_12 ));
    CascadeMux I__4701 (
            .O(N__25481),
            .I(\ALU.c_RNIJ949Z0Z_12_cascade_ ));
    InMux I__4700 (
            .O(N__25478),
            .I(N__25475));
    LocalMux I__4699 (
            .O(N__25475),
            .I(\ALU.a_RNIFPBOZ0Z_12 ));
    InMux I__4698 (
            .O(N__25472),
            .I(N__25469));
    LocalMux I__4697 (
            .O(N__25469),
            .I(\ALU.d_RNIM5LUZ0Z_12 ));
    CascadeMux I__4696 (
            .O(N__25466),
            .I(\ALU.operand2_7_ns_1_12_cascade_ ));
    InMux I__4695 (
            .O(N__25463),
            .I(N__25454));
    InMux I__4694 (
            .O(N__25462),
            .I(N__25454));
    InMux I__4693 (
            .O(N__25461),
            .I(N__25454));
    LocalMux I__4692 (
            .O(N__25454),
            .I(N__25449));
    InMux I__4691 (
            .O(N__25453),
            .I(N__25446));
    InMux I__4690 (
            .O(N__25452),
            .I(N__25443));
    Span4Mux_h I__4689 (
            .O(N__25449),
            .I(N__25439));
    LocalMux I__4688 (
            .O(N__25446),
            .I(N__25434));
    LocalMux I__4687 (
            .O(N__25443),
            .I(N__25434));
    InMux I__4686 (
            .O(N__25442),
            .I(N__25431));
    Span4Mux_h I__4685 (
            .O(N__25439),
            .I(N__25428));
    Span4Mux_v I__4684 (
            .O(N__25434),
            .I(N__25423));
    LocalMux I__4683 (
            .O(N__25431),
            .I(N__25423));
    Odrv4 I__4682 (
            .O(N__25428),
            .I(\ALU.operand2_12 ));
    Odrv4 I__4681 (
            .O(N__25423),
            .I(\ALU.operand2_12 ));
    CascadeMux I__4680 (
            .O(N__25418),
            .I(\ALU.N_636_cascade_ ));
    InMux I__4679 (
            .O(N__25415),
            .I(N__25412));
    LocalMux I__4678 (
            .O(N__25412),
            .I(N__25409));
    Span4Mux_h I__4677 (
            .O(N__25409),
            .I(N__25406));
    Span4Mux_h I__4676 (
            .O(N__25406),
            .I(N__25403));
    Span4Mux_v I__4675 (
            .O(N__25403),
            .I(N__25400));
    Span4Mux_v I__4674 (
            .O(N__25400),
            .I(N__25397));
    Odrv4 I__4673 (
            .O(N__25397),
            .I(\ALU.N_272_0 ));
    InMux I__4672 (
            .O(N__25394),
            .I(N__25391));
    LocalMux I__4671 (
            .O(N__25391),
            .I(N__25388));
    Span4Mux_h I__4670 (
            .O(N__25388),
            .I(N__25385));
    Span4Mux_h I__4669 (
            .O(N__25385),
            .I(N__25382));
    Odrv4 I__4668 (
            .O(N__25382),
            .I(\ALU.N_264_0 ));
    InMux I__4667 (
            .O(N__25379),
            .I(N__25374));
    InMux I__4666 (
            .O(N__25378),
            .I(N__25367));
    InMux I__4665 (
            .O(N__25377),
            .I(N__25364));
    LocalMux I__4664 (
            .O(N__25374),
            .I(N__25361));
    InMux I__4663 (
            .O(N__25373),
            .I(N__25356));
    InMux I__4662 (
            .O(N__25372),
            .I(N__25356));
    CascadeMux I__4661 (
            .O(N__25371),
            .I(N__25349));
    InMux I__4660 (
            .O(N__25370),
            .I(N__25345));
    LocalMux I__4659 (
            .O(N__25367),
            .I(N__25335));
    LocalMux I__4658 (
            .O(N__25364),
            .I(N__25335));
    Span4Mux_h I__4657 (
            .O(N__25361),
            .I(N__25330));
    LocalMux I__4656 (
            .O(N__25356),
            .I(N__25330));
    InMux I__4655 (
            .O(N__25355),
            .I(N__25327));
    InMux I__4654 (
            .O(N__25354),
            .I(N__25323));
    InMux I__4653 (
            .O(N__25353),
            .I(N__25316));
    InMux I__4652 (
            .O(N__25352),
            .I(N__25316));
    InMux I__4651 (
            .O(N__25349),
            .I(N__25316));
    InMux I__4650 (
            .O(N__25348),
            .I(N__25313));
    LocalMux I__4649 (
            .O(N__25345),
            .I(N__25310));
    InMux I__4648 (
            .O(N__25344),
            .I(N__25301));
    InMux I__4647 (
            .O(N__25343),
            .I(N__25301));
    InMux I__4646 (
            .O(N__25342),
            .I(N__25301));
    InMux I__4645 (
            .O(N__25341),
            .I(N__25301));
    InMux I__4644 (
            .O(N__25340),
            .I(N__25298));
    Span4Mux_v I__4643 (
            .O(N__25335),
            .I(N__25295));
    Span4Mux_h I__4642 (
            .O(N__25330),
            .I(N__25290));
    LocalMux I__4641 (
            .O(N__25327),
            .I(N__25290));
    InMux I__4640 (
            .O(N__25326),
            .I(N__25285));
    LocalMux I__4639 (
            .O(N__25323),
            .I(N__25282));
    LocalMux I__4638 (
            .O(N__25316),
            .I(N__25279));
    LocalMux I__4637 (
            .O(N__25313),
            .I(N__25274));
    Span4Mux_v I__4636 (
            .O(N__25310),
            .I(N__25274));
    LocalMux I__4635 (
            .O(N__25301),
            .I(N__25269));
    LocalMux I__4634 (
            .O(N__25298),
            .I(N__25269));
    Span4Mux_h I__4633 (
            .O(N__25295),
            .I(N__25264));
    Span4Mux_v I__4632 (
            .O(N__25290),
            .I(N__25264));
    InMux I__4631 (
            .O(N__25289),
            .I(N__25259));
    InMux I__4630 (
            .O(N__25288),
            .I(N__25259));
    LocalMux I__4629 (
            .O(N__25285),
            .I(N__25252));
    Span4Mux_v I__4628 (
            .O(N__25282),
            .I(N__25252));
    Span4Mux_s3_h I__4627 (
            .O(N__25279),
            .I(N__25252));
    Odrv4 I__4626 (
            .O(N__25274),
            .I(\ALU.aluOut_12 ));
    Odrv4 I__4625 (
            .O(N__25269),
            .I(\ALU.aluOut_12 ));
    Odrv4 I__4624 (
            .O(N__25264),
            .I(\ALU.aluOut_12 ));
    LocalMux I__4623 (
            .O(N__25259),
            .I(\ALU.aluOut_12 ));
    Odrv4 I__4622 (
            .O(N__25252),
            .I(\ALU.aluOut_12 ));
    InMux I__4621 (
            .O(N__25241),
            .I(N__25238));
    LocalMux I__4620 (
            .O(N__25238),
            .I(\ALU.N_462 ));
    InMux I__4619 (
            .O(N__25235),
            .I(N__25232));
    LocalMux I__4618 (
            .O(N__25232),
            .I(\ALU.N_270_0 ));
    InMux I__4617 (
            .O(N__25229),
            .I(N__25226));
    LocalMux I__4616 (
            .O(N__25226),
            .I(N__25222));
    InMux I__4615 (
            .O(N__25225),
            .I(N__25217));
    Span4Mux_v I__4614 (
            .O(N__25222),
            .I(N__25210));
    InMux I__4613 (
            .O(N__25221),
            .I(N__25207));
    InMux I__4612 (
            .O(N__25220),
            .I(N__25201));
    LocalMux I__4611 (
            .O(N__25217),
            .I(N__25198));
    InMux I__4610 (
            .O(N__25216),
            .I(N__25195));
    InMux I__4609 (
            .O(N__25215),
            .I(N__25192));
    InMux I__4608 (
            .O(N__25214),
            .I(N__25189));
    InMux I__4607 (
            .O(N__25213),
            .I(N__25186));
    Span4Mux_s1_h I__4606 (
            .O(N__25210),
            .I(N__25183));
    LocalMux I__4605 (
            .O(N__25207),
            .I(N__25180));
    InMux I__4604 (
            .O(N__25206),
            .I(N__25177));
    InMux I__4603 (
            .O(N__25205),
            .I(N__25174));
    InMux I__4602 (
            .O(N__25204),
            .I(N__25171));
    LocalMux I__4601 (
            .O(N__25201),
            .I(N__25166));
    Span4Mux_v I__4600 (
            .O(N__25198),
            .I(N__25159));
    LocalMux I__4599 (
            .O(N__25195),
            .I(N__25159));
    LocalMux I__4598 (
            .O(N__25192),
            .I(N__25156));
    LocalMux I__4597 (
            .O(N__25189),
            .I(N__25151));
    LocalMux I__4596 (
            .O(N__25186),
            .I(N__25151));
    Sp12to4 I__4595 (
            .O(N__25183),
            .I(N__25148));
    Span4Mux_h I__4594 (
            .O(N__25180),
            .I(N__25145));
    LocalMux I__4593 (
            .O(N__25177),
            .I(N__25140));
    LocalMux I__4592 (
            .O(N__25174),
            .I(N__25140));
    LocalMux I__4591 (
            .O(N__25171),
            .I(N__25136));
    InMux I__4590 (
            .O(N__25170),
            .I(N__25133));
    InMux I__4589 (
            .O(N__25169),
            .I(N__25130));
    Span4Mux_h I__4588 (
            .O(N__25166),
            .I(N__25127));
    CascadeMux I__4587 (
            .O(N__25165),
            .I(N__25124));
    CascadeMux I__4586 (
            .O(N__25164),
            .I(N__25119));
    Span4Mux_h I__4585 (
            .O(N__25159),
            .I(N__25111));
    Span4Mux_v I__4584 (
            .O(N__25156),
            .I(N__25111));
    Span4Mux_h I__4583 (
            .O(N__25151),
            .I(N__25111));
    Span12Mux_s4_h I__4582 (
            .O(N__25148),
            .I(N__25108));
    Span4Mux_v I__4581 (
            .O(N__25145),
            .I(N__25103));
    Span4Mux_h I__4580 (
            .O(N__25140),
            .I(N__25103));
    InMux I__4579 (
            .O(N__25139),
            .I(N__25100));
    Span12Mux_h I__4578 (
            .O(N__25136),
            .I(N__25091));
    LocalMux I__4577 (
            .O(N__25133),
            .I(N__25091));
    LocalMux I__4576 (
            .O(N__25130),
            .I(N__25091));
    Sp12to4 I__4575 (
            .O(N__25127),
            .I(N__25091));
    InMux I__4574 (
            .O(N__25124),
            .I(N__25084));
    InMux I__4573 (
            .O(N__25123),
            .I(N__25084));
    InMux I__4572 (
            .O(N__25122),
            .I(N__25084));
    InMux I__4571 (
            .O(N__25119),
            .I(N__25079));
    InMux I__4570 (
            .O(N__25118),
            .I(N__25079));
    Span4Mux_v I__4569 (
            .O(N__25111),
            .I(N__25076));
    Odrv12 I__4568 (
            .O(N__25108),
            .I(aluReadBus_fast));
    Odrv4 I__4567 (
            .O(N__25103),
            .I(aluReadBus_fast));
    LocalMux I__4566 (
            .O(N__25100),
            .I(aluReadBus_fast));
    Odrv12 I__4565 (
            .O(N__25091),
            .I(aluReadBus_fast));
    LocalMux I__4564 (
            .O(N__25084),
            .I(aluReadBus_fast));
    LocalMux I__4563 (
            .O(N__25079),
            .I(aluReadBus_fast));
    Odrv4 I__4562 (
            .O(N__25076),
            .I(aluReadBus_fast));
    InMux I__4561 (
            .O(N__25061),
            .I(N__25057));
    InMux I__4560 (
            .O(N__25060),
            .I(N__25054));
    LocalMux I__4559 (
            .O(N__25057),
            .I(N__25049));
    LocalMux I__4558 (
            .O(N__25054),
            .I(N__25046));
    InMux I__4557 (
            .O(N__25053),
            .I(N__25043));
    CascadeMux I__4556 (
            .O(N__25052),
            .I(N__25040));
    Span4Mux_h I__4555 (
            .O(N__25049),
            .I(N__25036));
    Span4Mux_h I__4554 (
            .O(N__25046),
            .I(N__25031));
    LocalMux I__4553 (
            .O(N__25043),
            .I(N__25031));
    InMux I__4552 (
            .O(N__25040),
            .I(N__25026));
    InMux I__4551 (
            .O(N__25039),
            .I(N__25026));
    Span4Mux_v I__4550 (
            .O(N__25036),
            .I(N__25023));
    Span4Mux_h I__4549 (
            .O(N__25031),
            .I(N__25020));
    LocalMux I__4548 (
            .O(N__25026),
            .I(\ALU.N_175_0 ));
    Odrv4 I__4547 (
            .O(N__25023),
            .I(\ALU.N_175_0 ));
    Odrv4 I__4546 (
            .O(N__25020),
            .I(\ALU.N_175_0 ));
    CascadeMux I__4545 (
            .O(N__25013),
            .I(\ALU.N_175_0_cascade_ ));
    InMux I__4544 (
            .O(N__25010),
            .I(N__25003));
    InMux I__4543 (
            .O(N__25009),
            .I(N__25003));
    InMux I__4542 (
            .O(N__25008),
            .I(N__25000));
    LocalMux I__4541 (
            .O(N__25003),
            .I(N__24996));
    LocalMux I__4540 (
            .O(N__25000),
            .I(N__24993));
    InMux I__4539 (
            .O(N__24999),
            .I(N__24990));
    Span4Mux_h I__4538 (
            .O(N__24996),
            .I(N__24985));
    Span4Mux_h I__4537 (
            .O(N__24993),
            .I(N__24985));
    LocalMux I__4536 (
            .O(N__24990),
            .I(\ALU.operand2_13 ));
    Odrv4 I__4535 (
            .O(N__24985),
            .I(\ALU.operand2_13 ));
    CascadeMux I__4534 (
            .O(N__24980),
            .I(\ALU.un2_addsub_axb_13_cascade_ ));
    InMux I__4533 (
            .O(N__24977),
            .I(N__24974));
    LocalMux I__4532 (
            .O(N__24974),
            .I(N__24970));
    InMux I__4531 (
            .O(N__24973),
            .I(N__24966));
    Span4Mux_v I__4530 (
            .O(N__24970),
            .I(N__24963));
    InMux I__4529 (
            .O(N__24969),
            .I(N__24960));
    LocalMux I__4528 (
            .O(N__24966),
            .I(N__24957));
    Span4Mux_h I__4527 (
            .O(N__24963),
            .I(N__24954));
    LocalMux I__4526 (
            .O(N__24960),
            .I(\ALU.N_177_0 ));
    Odrv4 I__4525 (
            .O(N__24957),
            .I(\ALU.N_177_0 ));
    Odrv4 I__4524 (
            .O(N__24954),
            .I(\ALU.N_177_0 ));
    CascadeMux I__4523 (
            .O(N__24947),
            .I(N__24944));
    InMux I__4522 (
            .O(N__24944),
            .I(N__24941));
    LocalMux I__4521 (
            .O(N__24941),
            .I(N__24938));
    Span4Mux_v I__4520 (
            .O(N__24938),
            .I(N__24935));
    Span4Mux_h I__4519 (
            .O(N__24935),
            .I(N__24932));
    Span4Mux_v I__4518 (
            .O(N__24932),
            .I(N__24929));
    Odrv4 I__4517 (
            .O(N__24929),
            .I(\ALU.d_RNI9FOTEZ0Z_13 ));
    InMux I__4516 (
            .O(N__24926),
            .I(N__24923));
    LocalMux I__4515 (
            .O(N__24923),
            .I(N__24919));
    InMux I__4514 (
            .O(N__24922),
            .I(N__24916));
    Span4Mux_v I__4513 (
            .O(N__24919),
            .I(N__24913));
    LocalMux I__4512 (
            .O(N__24916),
            .I(N__24910));
    Span4Mux_v I__4511 (
            .O(N__24913),
            .I(N__24906));
    Span4Mux_v I__4510 (
            .O(N__24910),
            .I(N__24902));
    InMux I__4509 (
            .O(N__24909),
            .I(N__24899));
    Span4Mux_h I__4508 (
            .O(N__24906),
            .I(N__24896));
    InMux I__4507 (
            .O(N__24905),
            .I(N__24893));
    Span4Mux_h I__4506 (
            .O(N__24902),
            .I(N__24889));
    LocalMux I__4505 (
            .O(N__24899),
            .I(N__24886));
    Span4Mux_v I__4504 (
            .O(N__24896),
            .I(N__24883));
    LocalMux I__4503 (
            .O(N__24893),
            .I(N__24880));
    CascadeMux I__4502 (
            .O(N__24892),
            .I(N__24877));
    Span4Mux_v I__4501 (
            .O(N__24889),
            .I(N__24872));
    Span4Mux_h I__4500 (
            .O(N__24886),
            .I(N__24872));
    Span4Mux_s1_h I__4499 (
            .O(N__24883),
            .I(N__24867));
    Span4Mux_h I__4498 (
            .O(N__24880),
            .I(N__24867));
    InMux I__4497 (
            .O(N__24877),
            .I(N__24864));
    Span4Mux_v I__4496 (
            .O(N__24872),
            .I(N__24861));
    Span4Mux_h I__4495 (
            .O(N__24867),
            .I(N__24858));
    LocalMux I__4494 (
            .O(N__24864),
            .I(N__24853));
    Span4Mux_h I__4493 (
            .O(N__24861),
            .I(N__24853));
    Odrv4 I__4492 (
            .O(N__24858),
            .I(ctrlOut_11));
    Odrv4 I__4491 (
            .O(N__24853),
            .I(ctrlOut_11));
    CascadeMux I__4490 (
            .O(N__24848),
            .I(N__24845));
    InMux I__4489 (
            .O(N__24845),
            .I(N__24842));
    LocalMux I__4488 (
            .O(N__24842),
            .I(N__24839));
    Span12Mux_s8_h I__4487 (
            .O(N__24839),
            .I(N__24836));
    Odrv12 I__4486 (
            .O(N__24836),
            .I(\ALU.N_186_0_i ));
    CascadeMux I__4485 (
            .O(N__24833),
            .I(\ALU.a_15_m4_bm_1Z0Z_2_cascade_ ));
    InMux I__4484 (
            .O(N__24830),
            .I(N__24827));
    LocalMux I__4483 (
            .O(N__24827),
            .I(N__24824));
    Odrv4 I__4482 (
            .O(N__24824),
            .I(\ALU.d_RNIII58AZ0Z_2 ));
    CascadeMux I__4481 (
            .O(N__24821),
            .I(\ALU.rshift_3_ns_1_2_cascade_ ));
    InMux I__4480 (
            .O(N__24818),
            .I(N__24815));
    LocalMux I__4479 (
            .O(N__24815),
            .I(N__24812));
    Odrv4 I__4478 (
            .O(N__24812),
            .I(\ALU.N_470 ));
    InMux I__4477 (
            .O(N__24809),
            .I(N__24806));
    LocalMux I__4476 (
            .O(N__24806),
            .I(N__24803));
    Span4Mux_v I__4475 (
            .O(N__24803),
            .I(N__24800));
    Odrv4 I__4474 (
            .O(N__24800),
            .I(\ALU.N_376 ));
    CascadeMux I__4473 (
            .O(N__24797),
            .I(\ALU.N_589_cascade_ ));
    CascadeMux I__4472 (
            .O(N__24794),
            .I(\ALU.rshift_1_13_cascade_ ));
    InMux I__4471 (
            .O(N__24791),
            .I(N__24788));
    LocalMux I__4470 (
            .O(N__24788),
            .I(N__24785));
    Span4Mux_h I__4469 (
            .O(N__24785),
            .I(N__24782));
    Odrv4 I__4468 (
            .O(N__24782),
            .I(\ALU.a_15_m3_13 ));
    CascadeMux I__4467 (
            .O(N__24779),
            .I(\ALU.N_576_cascade_ ));
    InMux I__4466 (
            .O(N__24776),
            .I(N__24773));
    LocalMux I__4465 (
            .O(N__24773),
            .I(N__24769));
    InMux I__4464 (
            .O(N__24772),
            .I(N__24763));
    Span4Mux_h I__4463 (
            .O(N__24769),
            .I(N__24760));
    InMux I__4462 (
            .O(N__24768),
            .I(N__24753));
    InMux I__4461 (
            .O(N__24767),
            .I(N__24753));
    InMux I__4460 (
            .O(N__24766),
            .I(N__24753));
    LocalMux I__4459 (
            .O(N__24763),
            .I(\FTDI.RXstateZ0Z_2 ));
    Odrv4 I__4458 (
            .O(N__24760),
            .I(\FTDI.RXstateZ0Z_2 ));
    LocalMux I__4457 (
            .O(N__24753),
            .I(\FTDI.RXstateZ0Z_2 ));
    CascadeMux I__4456 (
            .O(N__24746),
            .I(\FTDI.N_23_cascade_ ));
    InMux I__4455 (
            .O(N__24743),
            .I(N__24733));
    InMux I__4454 (
            .O(N__24742),
            .I(N__24733));
    InMux I__4453 (
            .O(N__24741),
            .I(N__24733));
    InMux I__4452 (
            .O(N__24740),
            .I(N__24730));
    LocalMux I__4451 (
            .O(N__24733),
            .I(N__24727));
    LocalMux I__4450 (
            .O(N__24730),
            .I(N__24724));
    Span4Mux_s1_v I__4449 (
            .O(N__24727),
            .I(N__24719));
    Span4Mux_s1_v I__4448 (
            .O(N__24724),
            .I(N__24716));
    InMux I__4447 (
            .O(N__24723),
            .I(N__24711));
    InMux I__4446 (
            .O(N__24722),
            .I(N__24711));
    Span4Mux_h I__4445 (
            .O(N__24719),
            .I(N__24708));
    Odrv4 I__4444 (
            .O(N__24716),
            .I(\FTDI.RXstateZ0Z_1 ));
    LocalMux I__4443 (
            .O(N__24711),
            .I(\FTDI.RXstateZ0Z_1 ));
    Odrv4 I__4442 (
            .O(N__24708),
            .I(\FTDI.RXstateZ0Z_1 ));
    InMux I__4441 (
            .O(N__24701),
            .I(N__24698));
    LocalMux I__4440 (
            .O(N__24698),
            .I(N__24695));
    Span4Mux_v I__4439 (
            .O(N__24695),
            .I(N__24692));
    Odrv4 I__4438 (
            .O(N__24692),
            .I(\FTDI.m13_ns_1 ));
    InMux I__4437 (
            .O(N__24689),
            .I(N__24683));
    InMux I__4436 (
            .O(N__24688),
            .I(N__24683));
    LocalMux I__4435 (
            .O(N__24683),
            .I(N__24677));
    InMux I__4434 (
            .O(N__24682),
            .I(N__24670));
    InMux I__4433 (
            .O(N__24681),
            .I(N__24670));
    InMux I__4432 (
            .O(N__24680),
            .I(N__24670));
    Span4Mux_s1_v I__4431 (
            .O(N__24677),
            .I(N__24667));
    LocalMux I__4430 (
            .O(N__24670),
            .I(\FTDI.RXstateZ0Z_0 ));
    Odrv4 I__4429 (
            .O(N__24667),
            .I(\FTDI.RXstateZ0Z_0 ));
    CascadeMux I__4428 (
            .O(N__24662),
            .I(N__24656));
    CascadeMux I__4427 (
            .O(N__24661),
            .I(N__24653));
    CascadeMux I__4426 (
            .O(N__24660),
            .I(N__24649));
    InMux I__4425 (
            .O(N__24659),
            .I(N__24646));
    InMux I__4424 (
            .O(N__24656),
            .I(N__24636));
    InMux I__4423 (
            .O(N__24653),
            .I(N__24636));
    InMux I__4422 (
            .O(N__24652),
            .I(N__24636));
    InMux I__4421 (
            .O(N__24649),
            .I(N__24636));
    LocalMux I__4420 (
            .O(N__24646),
            .I(N__24633));
    CascadeMux I__4419 (
            .O(N__24645),
            .I(N__24628));
    LocalMux I__4418 (
            .O(N__24636),
            .I(N__24624));
    Span4Mux_s1_v I__4417 (
            .O(N__24633),
            .I(N__24621));
    InMux I__4416 (
            .O(N__24632),
            .I(N__24612));
    InMux I__4415 (
            .O(N__24631),
            .I(N__24612));
    InMux I__4414 (
            .O(N__24628),
            .I(N__24612));
    InMux I__4413 (
            .O(N__24627),
            .I(N__24612));
    Span4Mux_s1_v I__4412 (
            .O(N__24624),
            .I(N__24609));
    Odrv4 I__4411 (
            .O(N__24621),
            .I(\FTDI.RXstateZ0Z_3 ));
    LocalMux I__4410 (
            .O(N__24612),
            .I(\FTDI.RXstateZ0Z_3 ));
    Odrv4 I__4409 (
            .O(N__24609),
            .I(\FTDI.RXstateZ0Z_3 ));
    CascadeMux I__4408 (
            .O(N__24602),
            .I(\ALU.a_15_sm0_cascade_ ));
    CascadeMux I__4407 (
            .O(N__24599),
            .I(\ALU.a_15_m2_ns_1Z0Z_12_cascade_ ));
    InMux I__4406 (
            .O(N__24596),
            .I(N__24589));
    InMux I__4405 (
            .O(N__24595),
            .I(N__24589));
    InMux I__4404 (
            .O(N__24594),
            .I(N__24584));
    LocalMux I__4403 (
            .O(N__24589),
            .I(N__24581));
    InMux I__4402 (
            .O(N__24588),
            .I(N__24574));
    InMux I__4401 (
            .O(N__24587),
            .I(N__24574));
    LocalMux I__4400 (
            .O(N__24584),
            .I(N__24571));
    Span4Mux_s2_v I__4399 (
            .O(N__24581),
            .I(N__24568));
    InMux I__4398 (
            .O(N__24580),
            .I(N__24563));
    InMux I__4397 (
            .O(N__24579),
            .I(N__24563));
    LocalMux I__4396 (
            .O(N__24574),
            .I(N__24558));
    Span4Mux_h I__4395 (
            .O(N__24571),
            .I(N__24558));
    Span4Mux_h I__4394 (
            .O(N__24568),
            .I(N__24555));
    LocalMux I__4393 (
            .O(N__24563),
            .I(N__24552));
    Odrv4 I__4392 (
            .O(N__24558),
            .I(\ALU.log_2_sqmuxa ));
    Odrv4 I__4391 (
            .O(N__24555),
            .I(\ALU.log_2_sqmuxa ));
    Odrv12 I__4390 (
            .O(N__24552),
            .I(\ALU.log_2_sqmuxa ));
    InMux I__4389 (
            .O(N__24545),
            .I(N__24542));
    LocalMux I__4388 (
            .O(N__24542),
            .I(N__24539));
    Span4Mux_v I__4387 (
            .O(N__24539),
            .I(N__24536));
    Odrv4 I__4386 (
            .O(N__24536),
            .I(\ALU.a7_b_0 ));
    InMux I__4385 (
            .O(N__24533),
            .I(N__24530));
    LocalMux I__4384 (
            .O(N__24530),
            .I(N__24527));
    Span4Mux_h I__4383 (
            .O(N__24527),
            .I(N__24523));
    InMux I__4382 (
            .O(N__24526),
            .I(N__24520));
    Odrv4 I__4381 (
            .O(N__24523),
            .I(\ALU.a5_b_2 ));
    LocalMux I__4380 (
            .O(N__24520),
            .I(\ALU.a5_b_2 ));
    CascadeMux I__4379 (
            .O(N__24515),
            .I(N__24512));
    InMux I__4378 (
            .O(N__24512),
            .I(N__24506));
    InMux I__4377 (
            .O(N__24511),
            .I(N__24506));
    LocalMux I__4376 (
            .O(N__24506),
            .I(N__24503));
    Odrv4 I__4375 (
            .O(N__24503),
            .I(\ALU.madd_63 ));
    InMux I__4374 (
            .O(N__24500),
            .I(N__24497));
    LocalMux I__4373 (
            .O(N__24497),
            .I(N__24494));
    Span4Mux_h I__4372 (
            .O(N__24494),
            .I(N__24491));
    Odrv4 I__4371 (
            .O(N__24491),
            .I(\ALU.a2_b_1 ));
    InMux I__4370 (
            .O(N__24488),
            .I(N__24485));
    LocalMux I__4369 (
            .O(N__24485),
            .I(N__24482));
    Span4Mux_h I__4368 (
            .O(N__24482),
            .I(N__24478));
    InMux I__4367 (
            .O(N__24481),
            .I(N__24475));
    Odrv4 I__4366 (
            .O(N__24478),
            .I(\ALU.a3_b_0 ));
    LocalMux I__4365 (
            .O(N__24475),
            .I(\ALU.a3_b_0 ));
    InMux I__4364 (
            .O(N__24470),
            .I(N__24467));
    LocalMux I__4363 (
            .O(N__24467),
            .I(N__24464));
    Span4Mux_v I__4362 (
            .O(N__24464),
            .I(N__24461));
    Span4Mux_h I__4361 (
            .O(N__24461),
            .I(N__24457));
    InMux I__4360 (
            .O(N__24460),
            .I(N__24454));
    Odrv4 I__4359 (
            .O(N__24457),
            .I(\ALU.a1_b_2 ));
    LocalMux I__4358 (
            .O(N__24454),
            .I(\ALU.a1_b_2 ));
    CascadeMux I__4357 (
            .O(N__24449),
            .I(N__24446));
    InMux I__4356 (
            .O(N__24446),
            .I(N__24443));
    LocalMux I__4355 (
            .O(N__24443),
            .I(N__24440));
    Span4Mux_v I__4354 (
            .O(N__24440),
            .I(N__24437));
    Span4Mux_v I__4353 (
            .O(N__24437),
            .I(N__24434));
    Odrv4 I__4352 (
            .O(N__24434),
            .I(\ALU.d_RNI2B0LZ0Z_9 ));
    InMux I__4351 (
            .O(N__24431),
            .I(N__24428));
    LocalMux I__4350 (
            .O(N__24428),
            .I(N__24424));
    CascadeMux I__4349 (
            .O(N__24427),
            .I(N__24420));
    Span4Mux_v I__4348 (
            .O(N__24424),
            .I(N__24417));
    InMux I__4347 (
            .O(N__24423),
            .I(N__24414));
    InMux I__4346 (
            .O(N__24420),
            .I(N__24411));
    Odrv4 I__4345 (
            .O(N__24417),
            .I(\ALU.hZ0Z_10 ));
    LocalMux I__4344 (
            .O(N__24414),
            .I(\ALU.hZ0Z_10 ));
    LocalMux I__4343 (
            .O(N__24411),
            .I(\ALU.hZ0Z_10 ));
    InMux I__4342 (
            .O(N__24404),
            .I(N__24401));
    LocalMux I__4341 (
            .O(N__24401),
            .I(N__24398));
    Span4Mux_h I__4340 (
            .O(N__24398),
            .I(N__24395));
    Span4Mux_v I__4339 (
            .O(N__24395),
            .I(N__24392));
    Odrv4 I__4338 (
            .O(N__24392),
            .I(\ALU.d_RNII1LUZ0Z_10 ));
    InMux I__4337 (
            .O(N__24389),
            .I(N__24386));
    LocalMux I__4336 (
            .O(N__24386),
            .I(N__24383));
    Span4Mux_v I__4335 (
            .O(N__24383),
            .I(N__24380));
    Odrv4 I__4334 (
            .O(N__24380),
            .I(\ALU.d_RNIO00LZ0Z_4 ));
    CascadeMux I__4333 (
            .O(N__24377),
            .I(N__24372));
    CascadeMux I__4332 (
            .O(N__24376),
            .I(N__24369));
    CascadeMux I__4331 (
            .O(N__24375),
            .I(N__24366));
    InMux I__4330 (
            .O(N__24372),
            .I(N__24361));
    InMux I__4329 (
            .O(N__24369),
            .I(N__24361));
    InMux I__4328 (
            .O(N__24366),
            .I(N__24358));
    LocalMux I__4327 (
            .O(N__24361),
            .I(N__24355));
    LocalMux I__4326 (
            .O(N__24358),
            .I(N__24352));
    Span4Mux_v I__4325 (
            .O(N__24355),
            .I(N__24349));
    Span4Mux_h I__4324 (
            .O(N__24352),
            .I(N__24346));
    Odrv4 I__4323 (
            .O(N__24349),
            .I(\ALU.a3_b_3 ));
    Odrv4 I__4322 (
            .O(N__24346),
            .I(\ALU.a3_b_3 ));
    CascadeMux I__4321 (
            .O(N__24341),
            .I(N__24337));
    CascadeMux I__4320 (
            .O(N__24340),
            .I(N__24334));
    InMux I__4319 (
            .O(N__24337),
            .I(N__24329));
    InMux I__4318 (
            .O(N__24334),
            .I(N__24329));
    LocalMux I__4317 (
            .O(N__24329),
            .I(N__24326));
    Span4Mux_v I__4316 (
            .O(N__24326),
            .I(N__24322));
    InMux I__4315 (
            .O(N__24325),
            .I(N__24319));
    Span4Mux_v I__4314 (
            .O(N__24322),
            .I(N__24308));
    LocalMux I__4313 (
            .O(N__24319),
            .I(N__24305));
    InMux I__4312 (
            .O(N__24318),
            .I(N__24302));
    CascadeMux I__4311 (
            .O(N__24317),
            .I(N__24299));
    CascadeMux I__4310 (
            .O(N__24316),
            .I(N__24294));
    CascadeMux I__4309 (
            .O(N__24315),
            .I(N__24291));
    CascadeMux I__4308 (
            .O(N__24314),
            .I(N__24287));
    CascadeMux I__4307 (
            .O(N__24313),
            .I(N__24284));
    CascadeMux I__4306 (
            .O(N__24312),
            .I(N__24280));
    InMux I__4305 (
            .O(N__24311),
            .I(N__24277));
    Span4Mux_h I__4304 (
            .O(N__24308),
            .I(N__24270));
    Span4Mux_v I__4303 (
            .O(N__24305),
            .I(N__24270));
    LocalMux I__4302 (
            .O(N__24302),
            .I(N__24270));
    InMux I__4301 (
            .O(N__24299),
            .I(N__24267));
    InMux I__4300 (
            .O(N__24298),
            .I(N__24264));
    InMux I__4299 (
            .O(N__24297),
            .I(N__24260));
    InMux I__4298 (
            .O(N__24294),
            .I(N__24257));
    InMux I__4297 (
            .O(N__24291),
            .I(N__24254));
    CascadeMux I__4296 (
            .O(N__24290),
            .I(N__24250));
    InMux I__4295 (
            .O(N__24287),
            .I(N__24246));
    InMux I__4294 (
            .O(N__24284),
            .I(N__24243));
    CascadeMux I__4293 (
            .O(N__24283),
            .I(N__24239));
    InMux I__4292 (
            .O(N__24280),
            .I(N__24236));
    LocalMux I__4291 (
            .O(N__24277),
            .I(N__24226));
    Span4Mux_v I__4290 (
            .O(N__24270),
            .I(N__24226));
    LocalMux I__4289 (
            .O(N__24267),
            .I(N__24223));
    LocalMux I__4288 (
            .O(N__24264),
            .I(N__24220));
    InMux I__4287 (
            .O(N__24263),
            .I(N__24217));
    LocalMux I__4286 (
            .O(N__24260),
            .I(N__24214));
    LocalMux I__4285 (
            .O(N__24257),
            .I(N__24209));
    LocalMux I__4284 (
            .O(N__24254),
            .I(N__24209));
    InMux I__4283 (
            .O(N__24253),
            .I(N__24202));
    InMux I__4282 (
            .O(N__24250),
            .I(N__24202));
    InMux I__4281 (
            .O(N__24249),
            .I(N__24202));
    LocalMux I__4280 (
            .O(N__24246),
            .I(N__24197));
    LocalMux I__4279 (
            .O(N__24243),
            .I(N__24197));
    CascadeMux I__4278 (
            .O(N__24242),
            .I(N__24194));
    InMux I__4277 (
            .O(N__24239),
            .I(N__24190));
    LocalMux I__4276 (
            .O(N__24236),
            .I(N__24187));
    CascadeMux I__4275 (
            .O(N__24235),
            .I(N__24184));
    InMux I__4274 (
            .O(N__24234),
            .I(N__24181));
    InMux I__4273 (
            .O(N__24233),
            .I(N__24176));
    InMux I__4272 (
            .O(N__24232),
            .I(N__24176));
    InMux I__4271 (
            .O(N__24231),
            .I(N__24173));
    IoSpan4Mux I__4270 (
            .O(N__24226),
            .I(N__24170));
    Span4Mux_v I__4269 (
            .O(N__24223),
            .I(N__24161));
    Span4Mux_s3_h I__4268 (
            .O(N__24220),
            .I(N__24161));
    LocalMux I__4267 (
            .O(N__24217),
            .I(N__24161));
    Span4Mux_s3_h I__4266 (
            .O(N__24214),
            .I(N__24161));
    Span4Mux_v I__4265 (
            .O(N__24209),
            .I(N__24154));
    LocalMux I__4264 (
            .O(N__24202),
            .I(N__24154));
    Span4Mux_v I__4263 (
            .O(N__24197),
            .I(N__24154));
    InMux I__4262 (
            .O(N__24194),
            .I(N__24150));
    CascadeMux I__4261 (
            .O(N__24193),
            .I(N__24145));
    LocalMux I__4260 (
            .O(N__24190),
            .I(N__24141));
    Span4Mux_h I__4259 (
            .O(N__24187),
            .I(N__24138));
    InMux I__4258 (
            .O(N__24184),
            .I(N__24135));
    LocalMux I__4257 (
            .O(N__24181),
            .I(N__24131));
    LocalMux I__4256 (
            .O(N__24176),
            .I(N__24128));
    LocalMux I__4255 (
            .O(N__24173),
            .I(N__24121));
    Span4Mux_s3_h I__4254 (
            .O(N__24170),
            .I(N__24121));
    Span4Mux_v I__4253 (
            .O(N__24161),
            .I(N__24121));
    Span4Mux_v I__4252 (
            .O(N__24154),
            .I(N__24118));
    InMux I__4251 (
            .O(N__24153),
            .I(N__24115));
    LocalMux I__4250 (
            .O(N__24150),
            .I(N__24112));
    InMux I__4249 (
            .O(N__24149),
            .I(N__24107));
    InMux I__4248 (
            .O(N__24148),
            .I(N__24107));
    InMux I__4247 (
            .O(N__24145),
            .I(N__24104));
    InMux I__4246 (
            .O(N__24144),
            .I(N__24101));
    Span12Mux_s4_h I__4245 (
            .O(N__24141),
            .I(N__24094));
    Sp12to4 I__4244 (
            .O(N__24138),
            .I(N__24094));
    LocalMux I__4243 (
            .O(N__24135),
            .I(N__24094));
    InMux I__4242 (
            .O(N__24134),
            .I(N__24091));
    Span4Mux_v I__4241 (
            .O(N__24131),
            .I(N__24082));
    Span4Mux_s3_h I__4240 (
            .O(N__24128),
            .I(N__24082));
    Span4Mux_v I__4239 (
            .O(N__24121),
            .I(N__24082));
    Span4Mux_h I__4238 (
            .O(N__24118),
            .I(N__24082));
    LocalMux I__4237 (
            .O(N__24115),
            .I(aluReadBus_rep1));
    Odrv12 I__4236 (
            .O(N__24112),
            .I(aluReadBus_rep1));
    LocalMux I__4235 (
            .O(N__24107),
            .I(aluReadBus_rep1));
    LocalMux I__4234 (
            .O(N__24104),
            .I(aluReadBus_rep1));
    LocalMux I__4233 (
            .O(N__24101),
            .I(aluReadBus_rep1));
    Odrv12 I__4232 (
            .O(N__24094),
            .I(aluReadBus_rep1));
    LocalMux I__4231 (
            .O(N__24091),
            .I(aluReadBus_rep1));
    Odrv4 I__4230 (
            .O(N__24082),
            .I(aluReadBus_rep1));
    CascadeMux I__4229 (
            .O(N__24065),
            .I(N__24061));
    InMux I__4228 (
            .O(N__24064),
            .I(N__24056));
    InMux I__4227 (
            .O(N__24061),
            .I(N__24056));
    LocalMux I__4226 (
            .O(N__24056),
            .I(N__24053));
    Span4Mux_h I__4225 (
            .O(N__24053),
            .I(N__24050));
    Span4Mux_h I__4224 (
            .O(N__24050),
            .I(N__24047));
    Odrv4 I__4223 (
            .O(N__24047),
            .I(\ALU.a2_b_3 ));
    InMux I__4222 (
            .O(N__24044),
            .I(N__24039));
    InMux I__4221 (
            .O(N__24043),
            .I(N__24034));
    InMux I__4220 (
            .O(N__24042),
            .I(N__24034));
    LocalMux I__4219 (
            .O(N__24039),
            .I(N__24031));
    LocalMux I__4218 (
            .O(N__24034),
            .I(N__24026));
    Span4Mux_v I__4217 (
            .O(N__24031),
            .I(N__24023));
    InMux I__4216 (
            .O(N__24030),
            .I(N__24019));
    InMux I__4215 (
            .O(N__24029),
            .I(N__24016));
    Span4Mux_v I__4214 (
            .O(N__24026),
            .I(N__24010));
    Span4Mux_v I__4213 (
            .O(N__24023),
            .I(N__24007));
    InMux I__4212 (
            .O(N__24022),
            .I(N__24004));
    LocalMux I__4211 (
            .O(N__24019),
            .I(N__24001));
    LocalMux I__4210 (
            .O(N__24016),
            .I(N__23998));
    InMux I__4209 (
            .O(N__24015),
            .I(N__23991));
    InMux I__4208 (
            .O(N__24014),
            .I(N__23991));
    InMux I__4207 (
            .O(N__24013),
            .I(N__23991));
    Span4Mux_v I__4206 (
            .O(N__24010),
            .I(N__23988));
    Sp12to4 I__4205 (
            .O(N__24007),
            .I(N__23983));
    LocalMux I__4204 (
            .O(N__24004),
            .I(N__23983));
    Span4Mux_h I__4203 (
            .O(N__24001),
            .I(N__23980));
    Span4Mux_h I__4202 (
            .O(N__23998),
            .I(N__23975));
    LocalMux I__4201 (
            .O(N__23991),
            .I(N__23975));
    Sp12to4 I__4200 (
            .O(N__23988),
            .I(N__23969));
    Span12Mux_s6_h I__4199 (
            .O(N__23983),
            .I(N__23964));
    Sp12to4 I__4198 (
            .O(N__23980),
            .I(N__23964));
    Span4Mux_v I__4197 (
            .O(N__23975),
            .I(N__23961));
    InMux I__4196 (
            .O(N__23974),
            .I(N__23954));
    InMux I__4195 (
            .O(N__23973),
            .I(N__23954));
    InMux I__4194 (
            .O(N__23972),
            .I(N__23954));
    Odrv12 I__4193 (
            .O(N__23969),
            .I(\ALU.operand2_3 ));
    Odrv12 I__4192 (
            .O(N__23964),
            .I(\ALU.operand2_3 ));
    Odrv4 I__4191 (
            .O(N__23961),
            .I(\ALU.operand2_3 ));
    LocalMux I__4190 (
            .O(N__23954),
            .I(\ALU.operand2_3 ));
    InMux I__4189 (
            .O(N__23945),
            .I(N__23941));
    InMux I__4188 (
            .O(N__23944),
            .I(N__23934));
    LocalMux I__4187 (
            .O(N__23941),
            .I(N__23931));
    InMux I__4186 (
            .O(N__23940),
            .I(N__23922));
    InMux I__4185 (
            .O(N__23939),
            .I(N__23922));
    InMux I__4184 (
            .O(N__23938),
            .I(N__23922));
    InMux I__4183 (
            .O(N__23937),
            .I(N__23922));
    LocalMux I__4182 (
            .O(N__23934),
            .I(N__23913));
    Span4Mux_v I__4181 (
            .O(N__23931),
            .I(N__23910));
    LocalMux I__4180 (
            .O(N__23922),
            .I(N__23907));
    CascadeMux I__4179 (
            .O(N__23921),
            .I(N__23904));
    InMux I__4178 (
            .O(N__23920),
            .I(N__23901));
    InMux I__4177 (
            .O(N__23919),
            .I(N__23894));
    InMux I__4176 (
            .O(N__23918),
            .I(N__23894));
    InMux I__4175 (
            .O(N__23917),
            .I(N__23894));
    InMux I__4174 (
            .O(N__23916),
            .I(N__23891));
    Span4Mux_v I__4173 (
            .O(N__23913),
            .I(N__23888));
    Span4Mux_s3_h I__4172 (
            .O(N__23910),
            .I(N__23885));
    Span4Mux_v I__4171 (
            .O(N__23907),
            .I(N__23882));
    InMux I__4170 (
            .O(N__23904),
            .I(N__23879));
    LocalMux I__4169 (
            .O(N__23901),
            .I(N__23876));
    LocalMux I__4168 (
            .O(N__23894),
            .I(N__23873));
    LocalMux I__4167 (
            .O(N__23891),
            .I(N__23868));
    Span4Mux_v I__4166 (
            .O(N__23888),
            .I(N__23868));
    Span4Mux_v I__4165 (
            .O(N__23885),
            .I(N__23863));
    Span4Mux_h I__4164 (
            .O(N__23882),
            .I(N__23863));
    LocalMux I__4163 (
            .O(N__23879),
            .I(\ALU.N_235_0 ));
    Odrv4 I__4162 (
            .O(N__23876),
            .I(\ALU.N_235_0 ));
    Odrv12 I__4161 (
            .O(N__23873),
            .I(\ALU.N_235_0 ));
    Odrv4 I__4160 (
            .O(N__23868),
            .I(\ALU.N_235_0 ));
    Odrv4 I__4159 (
            .O(N__23863),
            .I(\ALU.N_235_0 ));
    InMux I__4158 (
            .O(N__23852),
            .I(N__23849));
    LocalMux I__4157 (
            .O(N__23849),
            .I(\ALU.un2_addsub_axb_3 ));
    CascadeMux I__4156 (
            .O(N__23846),
            .I(N__23843));
    InMux I__4155 (
            .O(N__23843),
            .I(N__23840));
    LocalMux I__4154 (
            .O(N__23840),
            .I(N__23837));
    Span4Mux_v I__4153 (
            .O(N__23837),
            .I(N__23834));
    Span4Mux_v I__4152 (
            .O(N__23834),
            .I(N__23831));
    Odrv4 I__4151 (
            .O(N__23831),
            .I(\ALU.d_RNIDK21BZ0Z_3 ));
    CascadeMux I__4150 (
            .O(N__23828),
            .I(\ALU.dout_3_ns_1_3_cascade_ ));
    InMux I__4149 (
            .O(N__23825),
            .I(N__23822));
    LocalMux I__4148 (
            .O(N__23822),
            .I(\ALU.N_702 ));
    InMux I__4147 (
            .O(N__23819),
            .I(N__23816));
    LocalMux I__4146 (
            .O(N__23816),
            .I(\ALU.g_RNII4LLZ0Z_3 ));
    CascadeMux I__4145 (
            .O(N__23813),
            .I(\ALU.e_RNITOVJZ0Z_3_cascade_ ));
    InMux I__4144 (
            .O(N__23810),
            .I(N__23807));
    LocalMux I__4143 (
            .O(N__23807),
            .I(\ALU.operand2_7_ns_1_3 ));
    InMux I__4142 (
            .O(N__23804),
            .I(N__23801));
    LocalMux I__4141 (
            .O(N__23801),
            .I(N__23798));
    Span12Mux_v I__4140 (
            .O(N__23798),
            .I(N__23795));
    Odrv12 I__4139 (
            .O(N__23795),
            .I(\ALU.un2_addsub_cry_6_c_RNIL4LMIZ0 ));
    CascadeMux I__4138 (
            .O(N__23792),
            .I(\ALU.operand2_3_ns_1_6_cascade_ ));
    InMux I__4137 (
            .O(N__23789),
            .I(N__23786));
    LocalMux I__4136 (
            .O(N__23786),
            .I(\ALU.N_817 ));
    InMux I__4135 (
            .O(N__23783),
            .I(N__23780));
    LocalMux I__4134 (
            .O(N__23780),
            .I(N__23776));
    InMux I__4133 (
            .O(N__23779),
            .I(N__23772));
    Span4Mux_s2_h I__4132 (
            .O(N__23776),
            .I(N__23769));
    InMux I__4131 (
            .O(N__23775),
            .I(N__23766));
    LocalMux I__4130 (
            .O(N__23772),
            .I(N__23761));
    Span4Mux_v I__4129 (
            .O(N__23769),
            .I(N__23761));
    LocalMux I__4128 (
            .O(N__23766),
            .I(N__23758));
    Span4Mux_h I__4127 (
            .O(N__23761),
            .I(N__23755));
    Odrv12 I__4126 (
            .O(N__23758),
            .I(\ALU.a6_b_6 ));
    Odrv4 I__4125 (
            .O(N__23755),
            .I(\ALU.a6_b_6 ));
    InMux I__4124 (
            .O(N__23750),
            .I(N__23746));
    InMux I__4123 (
            .O(N__23749),
            .I(N__23743));
    LocalMux I__4122 (
            .O(N__23746),
            .I(N__23740));
    LocalMux I__4121 (
            .O(N__23743),
            .I(N__23737));
    Span4Mux_s3_h I__4120 (
            .O(N__23740),
            .I(N__23734));
    Span4Mux_s3_h I__4119 (
            .O(N__23737),
            .I(N__23731));
    Span4Mux_v I__4118 (
            .O(N__23734),
            .I(N__23728));
    Span4Mux_h I__4117 (
            .O(N__23731),
            .I(N__23723));
    Span4Mux_h I__4116 (
            .O(N__23728),
            .I(N__23723));
    Odrv4 I__4115 (
            .O(N__23723),
            .I(\ALU.a3_b_6 ));
    InMux I__4114 (
            .O(N__23720),
            .I(N__23717));
    LocalMux I__4113 (
            .O(N__23717),
            .I(\ALU.operand2_6_ns_1_6 ));
    CascadeMux I__4112 (
            .O(N__23714),
            .I(\ALU.N_750_cascade_ ));
    CascadeMux I__4111 (
            .O(N__23711),
            .I(\ALU.operand2_3_cascade_ ));
    InMux I__4110 (
            .O(N__23708),
            .I(N__23703));
    InMux I__4109 (
            .O(N__23707),
            .I(N__23700));
    InMux I__4108 (
            .O(N__23706),
            .I(N__23697));
    LocalMux I__4107 (
            .O(N__23703),
            .I(N__23694));
    LocalMux I__4106 (
            .O(N__23700),
            .I(N__23691));
    LocalMux I__4105 (
            .O(N__23697),
            .I(N__23688));
    Span4Mux_h I__4104 (
            .O(N__23694),
            .I(N__23685));
    Odrv4 I__4103 (
            .O(N__23691),
            .I(\ALU.aZ0Z_10 ));
    Odrv12 I__4102 (
            .O(N__23688),
            .I(\ALU.aZ0Z_10 ));
    Odrv4 I__4101 (
            .O(N__23685),
            .I(\ALU.aZ0Z_10 ));
    CascadeMux I__4100 (
            .O(N__23678),
            .I(\ALU.dout_3_ns_1_10_cascade_ ));
    CascadeMux I__4099 (
            .O(N__23675),
            .I(\ALU.dout_6_ns_1_10_cascade_ ));
    CascadeMux I__4098 (
            .O(N__23672),
            .I(\ALU.N_757_cascade_ ));
    InMux I__4097 (
            .O(N__23669),
            .I(N__23666));
    LocalMux I__4096 (
            .O(N__23666),
            .I(\ALU.N_709 ));
    InMux I__4095 (
            .O(N__23663),
            .I(N__23660));
    LocalMux I__4094 (
            .O(N__23660),
            .I(N__23657));
    Span4Mux_h I__4093 (
            .O(N__23657),
            .I(N__23654));
    Odrv4 I__4092 (
            .O(N__23654),
            .I(\ALU.dout_6_ns_1_5 ));
    CascadeMux I__4091 (
            .O(N__23651),
            .I(\ALU.N_865_cascade_ ));
    CascadeMux I__4090 (
            .O(N__23648),
            .I(\ALU.d_RNI61SHAZ0Z_1_cascade_ ));
    InMux I__4089 (
            .O(N__23645),
            .I(N__23642));
    LocalMux I__4088 (
            .O(N__23642),
            .I(\ALU.d_RNIJM067Z0Z_1 ));
    InMux I__4087 (
            .O(N__23639),
            .I(N__23636));
    LocalMux I__4086 (
            .O(N__23636),
            .I(N__23633));
    Span12Mux_s4_v I__4085 (
            .O(N__23633),
            .I(N__23630));
    Odrv12 I__4084 (
            .O(N__23630),
            .I(\ALU.a_15_m2_1 ));
    CascadeMux I__4083 (
            .O(N__23627),
            .I(\ALU.g_RNIK6LLZ0Z_4_cascade_ ));
    InMux I__4082 (
            .O(N__23624),
            .I(N__23621));
    LocalMux I__4081 (
            .O(N__23621),
            .I(\ALU.e_RNIGQ8HZ0Z_4 ));
    InMux I__4080 (
            .O(N__23618),
            .I(N__23612));
    InMux I__4079 (
            .O(N__23617),
            .I(N__23612));
    LocalMux I__4078 (
            .O(N__23612),
            .I(N__23609));
    Odrv12 I__4077 (
            .O(N__23609),
            .I(\ALU.a1_b_4 ));
    InMux I__4076 (
            .O(N__23606),
            .I(N__23602));
    InMux I__4075 (
            .O(N__23605),
            .I(N__23599));
    LocalMux I__4074 (
            .O(N__23602),
            .I(N__23596));
    LocalMux I__4073 (
            .O(N__23599),
            .I(N__23593));
    Span4Mux_v I__4072 (
            .O(N__23596),
            .I(N__23590));
    Span4Mux_h I__4071 (
            .O(N__23593),
            .I(N__23587));
    Span4Mux_h I__4070 (
            .O(N__23590),
            .I(N__23584));
    Odrv4 I__4069 (
            .O(N__23587),
            .I(\ALU.a2_b_4 ));
    Odrv4 I__4068 (
            .O(N__23584),
            .I(\ALU.a2_b_4 ));
    InMux I__4067 (
            .O(N__23579),
            .I(N__23576));
    LocalMux I__4066 (
            .O(N__23576),
            .I(\ALU.operand2_7_ns_1_4 ));
    InMux I__4065 (
            .O(N__23573),
            .I(N__23570));
    LocalMux I__4064 (
            .O(N__23570),
            .I(N__23563));
    InMux I__4063 (
            .O(N__23569),
            .I(N__23560));
    InMux I__4062 (
            .O(N__23568),
            .I(N__23555));
    InMux I__4061 (
            .O(N__23567),
            .I(N__23552));
    InMux I__4060 (
            .O(N__23566),
            .I(N__23549));
    Span4Mux_v I__4059 (
            .O(N__23563),
            .I(N__23544));
    LocalMux I__4058 (
            .O(N__23560),
            .I(N__23544));
    InMux I__4057 (
            .O(N__23559),
            .I(N__23539));
    InMux I__4056 (
            .O(N__23558),
            .I(N__23539));
    LocalMux I__4055 (
            .O(N__23555),
            .I(N__23534));
    LocalMux I__4054 (
            .O(N__23552),
            .I(N__23534));
    LocalMux I__4053 (
            .O(N__23549),
            .I(N__23531));
    Span4Mux_v I__4052 (
            .O(N__23544),
            .I(N__23528));
    LocalMux I__4051 (
            .O(N__23539),
            .I(N__23525));
    Span4Mux_h I__4050 (
            .O(N__23534),
            .I(N__23520));
    Span4Mux_h I__4049 (
            .O(N__23531),
            .I(N__23513));
    Span4Mux_h I__4048 (
            .O(N__23528),
            .I(N__23513));
    Span4Mux_v I__4047 (
            .O(N__23525),
            .I(N__23513));
    InMux I__4046 (
            .O(N__23524),
            .I(N__23508));
    InMux I__4045 (
            .O(N__23523),
            .I(N__23508));
    Odrv4 I__4044 (
            .O(N__23520),
            .I(\ALU.operand2_4 ));
    Odrv4 I__4043 (
            .O(N__23513),
            .I(\ALU.operand2_4 ));
    LocalMux I__4042 (
            .O(N__23508),
            .I(\ALU.operand2_4 ));
    InMux I__4041 (
            .O(N__23501),
            .I(N__23497));
    CascadeMux I__4040 (
            .O(N__23500),
            .I(N__23494));
    LocalMux I__4039 (
            .O(N__23497),
            .I(N__23490));
    InMux I__4038 (
            .O(N__23494),
            .I(N__23480));
    InMux I__4037 (
            .O(N__23493),
            .I(N__23480));
    Span4Mux_s2_h I__4036 (
            .O(N__23490),
            .I(N__23477));
    CascadeMux I__4035 (
            .O(N__23489),
            .I(N__23474));
    InMux I__4034 (
            .O(N__23488),
            .I(N__23469));
    InMux I__4033 (
            .O(N__23487),
            .I(N__23469));
    InMux I__4032 (
            .O(N__23486),
            .I(N__23465));
    InMux I__4031 (
            .O(N__23485),
            .I(N__23462));
    LocalMux I__4030 (
            .O(N__23480),
            .I(N__23457));
    Span4Mux_h I__4029 (
            .O(N__23477),
            .I(N__23457));
    InMux I__4028 (
            .O(N__23474),
            .I(N__23453));
    LocalMux I__4027 (
            .O(N__23469),
            .I(N__23450));
    InMux I__4026 (
            .O(N__23468),
            .I(N__23447));
    LocalMux I__4025 (
            .O(N__23465),
            .I(N__23443));
    LocalMux I__4024 (
            .O(N__23462),
            .I(N__23440));
    Sp12to4 I__4023 (
            .O(N__23457),
            .I(N__23437));
    InMux I__4022 (
            .O(N__23456),
            .I(N__23434));
    LocalMux I__4021 (
            .O(N__23453),
            .I(N__23429));
    Span4Mux_h I__4020 (
            .O(N__23450),
            .I(N__23429));
    LocalMux I__4019 (
            .O(N__23447),
            .I(N__23426));
    InMux I__4018 (
            .O(N__23446),
            .I(N__23423));
    Span12Mux_s3_h I__4017 (
            .O(N__23443),
            .I(N__23420));
    Span4Mux_v I__4016 (
            .O(N__23440),
            .I(N__23417));
    Span12Mux_v I__4015 (
            .O(N__23437),
            .I(N__23414));
    LocalMux I__4014 (
            .O(N__23434),
            .I(N__23409));
    Span4Mux_v I__4013 (
            .O(N__23429),
            .I(N__23409));
    Odrv4 I__4012 (
            .O(N__23426),
            .I(\ALU.N_229_0 ));
    LocalMux I__4011 (
            .O(N__23423),
            .I(\ALU.N_229_0 ));
    Odrv12 I__4010 (
            .O(N__23420),
            .I(\ALU.N_229_0 ));
    Odrv4 I__4009 (
            .O(N__23417),
            .I(\ALU.N_229_0 ));
    Odrv12 I__4008 (
            .O(N__23414),
            .I(\ALU.N_229_0 ));
    Odrv4 I__4007 (
            .O(N__23409),
            .I(\ALU.N_229_0 ));
    CascadeMux I__4006 (
            .O(N__23396),
            .I(\ALU.operand2_4_cascade_ ));
    CascadeMux I__4005 (
            .O(N__23393),
            .I(\ALU.N_231_0_cascade_ ));
    InMux I__4004 (
            .O(N__23390),
            .I(N__23387));
    LocalMux I__4003 (
            .O(N__23387),
            .I(N__23384));
    Span4Mux_h I__4002 (
            .O(N__23384),
            .I(N__23381));
    Odrv4 I__4001 (
            .O(N__23381),
            .I(\ALU.madd_93_0 ));
    InMux I__4000 (
            .O(N__23378),
            .I(N__23375));
    LocalMux I__3999 (
            .O(N__23375),
            .I(\ALU.N_758 ));
    CascadeMux I__3998 (
            .O(N__23372),
            .I(\ALU.N_710_cascade_ ));
    CascadeMux I__3997 (
            .O(N__23369),
            .I(\ALU.aluOut_11_cascade_ ));
    InMux I__3996 (
            .O(N__23366),
            .I(N__23363));
    LocalMux I__3995 (
            .O(N__23363),
            .I(N__23360));
    Span4Mux_h I__3994 (
            .O(N__23360),
            .I(N__23357));
    Odrv4 I__3993 (
            .O(N__23357),
            .I(\ALU.madd_484_6 ));
    CascadeMux I__3992 (
            .O(N__23354),
            .I(\ALU.un2_addsub_axb_1_cascade_ ));
    InMux I__3991 (
            .O(N__23351),
            .I(N__23348));
    LocalMux I__3990 (
            .O(N__23348),
            .I(\ALU.d_RNIC4AT9Z0Z_1 ));
    CascadeMux I__3989 (
            .O(N__23345),
            .I(\ALU.dout_7_ns_1_1_cascade_ ));
    InMux I__3988 (
            .O(N__23342),
            .I(N__23339));
    LocalMux I__3987 (
            .O(N__23339),
            .I(N__23333));
    InMux I__3986 (
            .O(N__23338),
            .I(N__23330));
    InMux I__3985 (
            .O(N__23337),
            .I(N__23327));
    InMux I__3984 (
            .O(N__23336),
            .I(N__23324));
    Span4Mux_h I__3983 (
            .O(N__23333),
            .I(N__23321));
    LocalMux I__3982 (
            .O(N__23330),
            .I(N__23316));
    LocalMux I__3981 (
            .O(N__23327),
            .I(N__23316));
    LocalMux I__3980 (
            .O(N__23324),
            .I(N__23313));
    Sp12to4 I__3979 (
            .O(N__23321),
            .I(N__23308));
    Span12Mux_h I__3978 (
            .O(N__23316),
            .I(N__23308));
    Sp12to4 I__3977 (
            .O(N__23313),
            .I(N__23305));
    Odrv12 I__3976 (
            .O(N__23308),
            .I(\ALU.N_247_0 ));
    Odrv12 I__3975 (
            .O(N__23305),
            .I(\ALU.N_247_0 ));
    InMux I__3974 (
            .O(N__23300),
            .I(N__23294));
    InMux I__3973 (
            .O(N__23299),
            .I(N__23294));
    LocalMux I__3972 (
            .O(N__23294),
            .I(N__23291));
    Span4Mux_h I__3971 (
            .O(N__23291),
            .I(N__23287));
    InMux I__3970 (
            .O(N__23290),
            .I(N__23284));
    Odrv4 I__3969 (
            .O(N__23287),
            .I(\ALU.operand2_1 ));
    LocalMux I__3968 (
            .O(N__23284),
            .I(\ALU.operand2_1 ));
    CascadeMux I__3967 (
            .O(N__23279),
            .I(N__23275));
    InMux I__3966 (
            .O(N__23278),
            .I(N__23272));
    InMux I__3965 (
            .O(N__23275),
            .I(N__23269));
    LocalMux I__3964 (
            .O(N__23272),
            .I(N__23266));
    LocalMux I__3963 (
            .O(N__23269),
            .I(\ALU.N_249_0 ));
    Odrv4 I__3962 (
            .O(N__23266),
            .I(\ALU.N_249_0 ));
    CascadeMux I__3961 (
            .O(N__23261),
            .I(\ALU.N_249_0_cascade_ ));
    InMux I__3960 (
            .O(N__23258),
            .I(N__23255));
    LocalMux I__3959 (
            .O(N__23255),
            .I(\ALU.a_15_m2_10 ));
    InMux I__3958 (
            .O(N__23252),
            .I(N__23249));
    LocalMux I__3957 (
            .O(N__23249),
            .I(\ALU.a_15_m2_ns_1Z0Z_10 ));
    InMux I__3956 (
            .O(N__23246),
            .I(N__23243));
    LocalMux I__3955 (
            .O(N__23243),
            .I(N__23240));
    Odrv4 I__3954 (
            .O(N__23240),
            .I(\ALU.un2_addsub_cry_9_c_RNIVCOFAZ0 ));
    CascadeMux I__3953 (
            .O(N__23237),
            .I(un9_addsub_cry_9_c_RNI8H83V_cascade_));
    InMux I__3952 (
            .O(N__23234),
            .I(N__23231));
    LocalMux I__3951 (
            .O(N__23231),
            .I(c_RNI5V90O2_10));
    CascadeMux I__3950 (
            .O(N__23228),
            .I(aluOperation_RNINNN4N3_0_cascade_));
    CascadeMux I__3949 (
            .O(N__23225),
            .I(\ALU.dout_6_ns_1_11_cascade_ ));
    CascadeMux I__3948 (
            .O(N__23222),
            .I(\ALU.dout_3_ns_1_11_cascade_ ));
    InMux I__3947 (
            .O(N__23219),
            .I(N__23216));
    LocalMux I__3946 (
            .O(N__23216),
            .I(N__23213));
    Span4Mux_v I__3945 (
            .O(N__23213),
            .I(N__23210));
    Span4Mux_v I__3944 (
            .O(N__23210),
            .I(N__23206));
    CascadeMux I__3943 (
            .O(N__23209),
            .I(N__23203));
    Sp12to4 I__3942 (
            .O(N__23206),
            .I(N__23200));
    InMux I__3941 (
            .O(N__23203),
            .I(N__23197));
    Odrv12 I__3940 (
            .O(N__23200),
            .I(\ALU.a0_b_4 ));
    LocalMux I__3939 (
            .O(N__23197),
            .I(\ALU.a0_b_4 ));
    CascadeMux I__3938 (
            .O(N__23192),
            .I(\ALU.a1_b_3_cascade_ ));
    InMux I__3937 (
            .O(N__23189),
            .I(N__23185));
    InMux I__3936 (
            .O(N__23188),
            .I(N__23182));
    LocalMux I__3935 (
            .O(N__23185),
            .I(N__23179));
    LocalMux I__3934 (
            .O(N__23182),
            .I(N__23176));
    Span4Mux_h I__3933 (
            .O(N__23179),
            .I(N__23173));
    Span4Mux_v I__3932 (
            .O(N__23176),
            .I(N__23170));
    Odrv4 I__3931 (
            .O(N__23173),
            .I(\ALU.madd_0 ));
    Odrv4 I__3930 (
            .O(N__23170),
            .I(\ALU.madd_0 ));
    InMux I__3929 (
            .O(N__23165),
            .I(N__23162));
    LocalMux I__3928 (
            .O(N__23162),
            .I(N__23159));
    Span4Mux_v I__3927 (
            .O(N__23159),
            .I(N__23155));
    InMux I__3926 (
            .O(N__23158),
            .I(N__23152));
    Span4Mux_h I__3925 (
            .O(N__23155),
            .I(N__23149));
    LocalMux I__3924 (
            .O(N__23152),
            .I(\ALU.a0_b_3 ));
    Odrv4 I__3923 (
            .O(N__23149),
            .I(\ALU.a0_b_3 ));
    InMux I__3922 (
            .O(N__23144),
            .I(N__23138));
    InMux I__3921 (
            .O(N__23143),
            .I(N__23134));
    InMux I__3920 (
            .O(N__23142),
            .I(N__23129));
    InMux I__3919 (
            .O(N__23141),
            .I(N__23129));
    LocalMux I__3918 (
            .O(N__23138),
            .I(N__23126));
    InMux I__3917 (
            .O(N__23137),
            .I(N__23123));
    LocalMux I__3916 (
            .O(N__23134),
            .I(N__23118));
    LocalMux I__3915 (
            .O(N__23129),
            .I(N__23118));
    Odrv12 I__3914 (
            .O(N__23126),
            .I(\ALU.N_375 ));
    LocalMux I__3913 (
            .O(N__23123),
            .I(\ALU.N_375 ));
    Odrv4 I__3912 (
            .O(N__23118),
            .I(\ALU.N_375 ));
    InMux I__3911 (
            .O(N__23111),
            .I(N__23108));
    LocalMux I__3910 (
            .O(N__23108),
            .I(\ALU.rshift_3_ns_1_0 ));
    InMux I__3909 (
            .O(N__23105),
            .I(N__23101));
    InMux I__3908 (
            .O(N__23104),
            .I(N__23098));
    LocalMux I__3907 (
            .O(N__23101),
            .I(N__23093));
    LocalMux I__3906 (
            .O(N__23098),
            .I(N__23093));
    Odrv4 I__3905 (
            .O(N__23093),
            .I(\ALU.N_249 ));
    InMux I__3904 (
            .O(N__23090),
            .I(N__23086));
    InMux I__3903 (
            .O(N__23089),
            .I(N__23083));
    LocalMux I__3902 (
            .O(N__23086),
            .I(\ALU.N_245 ));
    LocalMux I__3901 (
            .O(N__23083),
            .I(\ALU.N_245 ));
    InMux I__3900 (
            .O(N__23078),
            .I(N__23075));
    LocalMux I__3899 (
            .O(N__23075),
            .I(N__23072));
    Odrv4 I__3898 (
            .O(N__23072),
            .I(\ALU.lshift_10 ));
    InMux I__3897 (
            .O(N__23069),
            .I(N__23066));
    LocalMux I__3896 (
            .O(N__23066),
            .I(N__23063));
    Span4Mux_v I__3895 (
            .O(N__23063),
            .I(N__23060));
    Odrv4 I__3894 (
            .O(N__23060),
            .I(\ALU.a_15_m3_10 ));
    CascadeMux I__3893 (
            .O(N__23057),
            .I(\ALU.a_15_m4_10_cascade_ ));
    InMux I__3892 (
            .O(N__23054),
            .I(N__23049));
    InMux I__3891 (
            .O(N__23053),
            .I(N__23044));
    InMux I__3890 (
            .O(N__23052),
            .I(N__23044));
    LocalMux I__3889 (
            .O(N__23049),
            .I(N__23040));
    LocalMux I__3888 (
            .O(N__23044),
            .I(N__23037));
    InMux I__3887 (
            .O(N__23043),
            .I(N__23034));
    Odrv12 I__3886 (
            .O(N__23040),
            .I(\ALU.N_377 ));
    Odrv4 I__3885 (
            .O(N__23037),
            .I(\ALU.N_377 ));
    LocalMux I__3884 (
            .O(N__23034),
            .I(\ALU.N_377 ));
    CascadeMux I__3883 (
            .O(N__23027),
            .I(\ALU.N_377_cascade_ ));
    InMux I__3882 (
            .O(N__23024),
            .I(N__23021));
    LocalMux I__3881 (
            .O(N__23021),
            .I(\ALU.N_216 ));
    InMux I__3880 (
            .O(N__23018),
            .I(N__23015));
    LocalMux I__3879 (
            .O(N__23015),
            .I(\ALU.N_404 ));
    InMux I__3878 (
            .O(N__23012),
            .I(N__23009));
    LocalMux I__3877 (
            .O(N__23009),
            .I(N__23005));
    InMux I__3876 (
            .O(N__23008),
            .I(N__23002));
    Odrv4 I__3875 (
            .O(N__23005),
            .I(\ALU.N_246 ));
    LocalMux I__3874 (
            .O(N__23002),
            .I(\ALU.N_246 ));
    CascadeMux I__3873 (
            .O(N__22997),
            .I(\ALU.N_376_cascade_ ));
    CascadeMux I__3872 (
            .O(N__22994),
            .I(\ALU.d_RNIEBMRAZ0Z_0_cascade_ ));
    InMux I__3871 (
            .O(N__22991),
            .I(N__22988));
    LocalMux I__3870 (
            .O(N__22988),
            .I(\ALU.d_RNI1GH4VZ0Z_7 ));
    InMux I__3869 (
            .O(N__22985),
            .I(N__22982));
    LocalMux I__3868 (
            .O(N__22982),
            .I(N__22979));
    Span4Mux_h I__3867 (
            .O(N__22979),
            .I(N__22976));
    Span4Mux_v I__3866 (
            .O(N__22976),
            .I(N__22973));
    Odrv4 I__3865 (
            .O(N__22973),
            .I(\ALU.N_468 ));
    InMux I__3864 (
            .O(N__22970),
            .I(N__22967));
    LocalMux I__3863 (
            .O(N__22967),
            .I(N__22964));
    Span4Mux_v I__3862 (
            .O(N__22964),
            .I(N__22961));
    Span4Mux_h I__3861 (
            .O(N__22961),
            .I(N__22958));
    Odrv4 I__3860 (
            .O(N__22958),
            .I(\ALU.a1_b_3 ));
    CascadeMux I__3859 (
            .O(N__22955),
            .I(\ALU.d_RNIA28GU1Z0Z_1_cascade_ ));
    InMux I__3858 (
            .O(N__22952),
            .I(N__22949));
    LocalMux I__3857 (
            .O(N__22949),
            .I(\ALU.d_RNIJ1PCQZ0Z_1 ));
    InMux I__3856 (
            .O(N__22946),
            .I(N__22943));
    LocalMux I__3855 (
            .O(N__22943),
            .I(N__22940));
    Span4Mux_v I__3854 (
            .O(N__22940),
            .I(N__22937));
    Odrv4 I__3853 (
            .O(N__22937),
            .I(\ALU.N_225 ));
    InMux I__3852 (
            .O(N__22934),
            .I(N__22930));
    InMux I__3851 (
            .O(N__22933),
            .I(N__22927));
    LocalMux I__3850 (
            .O(N__22930),
            .I(N__22924));
    LocalMux I__3849 (
            .O(N__22927),
            .I(\ALU.N_223 ));
    Odrv4 I__3848 (
            .O(N__22924),
            .I(\ALU.N_223 ));
    InMux I__3847 (
            .O(N__22919),
            .I(N__22916));
    LocalMux I__3846 (
            .O(N__22916),
            .I(N__22912));
    InMux I__3845 (
            .O(N__22915),
            .I(N__22909));
    Span4Mux_h I__3844 (
            .O(N__22912),
            .I(N__22906));
    LocalMux I__3843 (
            .O(N__22909),
            .I(N__22903));
    Odrv4 I__3842 (
            .O(N__22906),
            .I(\ALU.N_221 ));
    Odrv4 I__3841 (
            .O(N__22903),
            .I(\ALU.N_221 ));
    CascadeMux I__3840 (
            .O(N__22898),
            .I(\ALU.lshift_7_ns_1_13_cascade_ ));
    InMux I__3839 (
            .O(N__22895),
            .I(N__22888));
    InMux I__3838 (
            .O(N__22894),
            .I(N__22888));
    InMux I__3837 (
            .O(N__22893),
            .I(N__22885));
    LocalMux I__3836 (
            .O(N__22888),
            .I(N__22882));
    LocalMux I__3835 (
            .O(N__22885),
            .I(N__22879));
    Span4Mux_h I__3834 (
            .O(N__22882),
            .I(N__22876));
    Odrv12 I__3833 (
            .O(N__22879),
            .I(\ALU.N_219 ));
    Odrv4 I__3832 (
            .O(N__22876),
            .I(\ALU.N_219 ));
    CascadeMux I__3831 (
            .O(N__22871),
            .I(\ALU.N_315_cascade_ ));
    CascadeMux I__3830 (
            .O(N__22868),
            .I(\ALU.lshift_13_cascade_ ));
    InMux I__3829 (
            .O(N__22865),
            .I(N__22862));
    LocalMux I__3828 (
            .O(N__22862),
            .I(N__22859));
    Odrv4 I__3827 (
            .O(N__22859),
            .I(\ALU.a_15_m2_13 ));
    CascadeMux I__3826 (
            .O(N__22856),
            .I(\ALU.a_15_m4_13_cascade_ ));
    InMux I__3825 (
            .O(N__22853),
            .I(N__22850));
    LocalMux I__3824 (
            .O(N__22850),
            .I(\ALU.N_247 ));
    InMux I__3823 (
            .O(N__22847),
            .I(N__22844));
    LocalMux I__3822 (
            .O(N__22844),
            .I(\ALU.lshift_15_ns_1_15 ));
    InMux I__3821 (
            .O(N__22841),
            .I(N__22835));
    InMux I__3820 (
            .O(N__22840),
            .I(N__22835));
    LocalMux I__3819 (
            .O(N__22835),
            .I(\ALU.N_416 ));
    CascadeMux I__3818 (
            .O(N__22832),
            .I(\ALU.rshift_3_ns_1_9_cascade_ ));
    InMux I__3817 (
            .O(N__22829),
            .I(N__22826));
    LocalMux I__3816 (
            .O(N__22826),
            .I(\ALU.rshift_3_ns_1_1 ));
    InMux I__3815 (
            .O(N__22823),
            .I(N__22820));
    LocalMux I__3814 (
            .O(N__22820),
            .I(N__22817));
    Odrv4 I__3813 (
            .O(N__22817),
            .I(\ALU.d_RNINEO9E_0Z0Z_1 ));
    InMux I__3812 (
            .O(N__22814),
            .I(N__22811));
    LocalMux I__3811 (
            .O(N__22811),
            .I(N__22807));
    InMux I__3810 (
            .O(N__22810),
            .I(N__22804));
    Span4Mux_v I__3809 (
            .O(N__22807),
            .I(N__22800));
    LocalMux I__3808 (
            .O(N__22804),
            .I(N__22797));
    InMux I__3807 (
            .O(N__22803),
            .I(N__22794));
    Odrv4 I__3806 (
            .O(N__22800),
            .I(\ALU.N_217 ));
    Odrv4 I__3805 (
            .O(N__22797),
            .I(\ALU.N_217 ));
    LocalMux I__3804 (
            .O(N__22794),
            .I(\ALU.N_217 ));
    InMux I__3803 (
            .O(N__22787),
            .I(N__22784));
    LocalMux I__3802 (
            .O(N__22784),
            .I(\ALU.lshift_7_ns_1_9 ));
    CascadeMux I__3801 (
            .O(N__22781),
            .I(\ALU.N_311_cascade_ ));
    CascadeMux I__3800 (
            .O(N__22778),
            .I(\ALU.lshift_9_cascade_ ));
    InMux I__3799 (
            .O(N__22775),
            .I(N__22772));
    LocalMux I__3798 (
            .O(N__22772),
            .I(N__22769));
    Span4Mux_h I__3797 (
            .O(N__22769),
            .I(N__22766));
    Odrv4 I__3796 (
            .O(N__22766),
            .I(\ALU.a_15_m2_9 ));
    InMux I__3795 (
            .O(N__22763),
            .I(N__22760));
    LocalMux I__3794 (
            .O(N__22760),
            .I(N__22757));
    Span4Mux_h I__3793 (
            .O(N__22757),
            .I(N__22754));
    Odrv4 I__3792 (
            .O(N__22754),
            .I(\ALU.N_292_0 ));
    InMux I__3791 (
            .O(N__22751),
            .I(N__22748));
    LocalMux I__3790 (
            .O(N__22748),
            .I(\ALU.rshift_1 ));
    CascadeMux I__3789 (
            .O(N__22745),
            .I(\ALU.N_473_cascade_ ));
    InMux I__3788 (
            .O(N__22742),
            .I(N__22739));
    LocalMux I__3787 (
            .O(N__22739),
            .I(\ALU.m42_nsZ0Z_1 ));
    CascadeMux I__3786 (
            .O(N__22736),
            .I(N__22733));
    InMux I__3785 (
            .O(N__22733),
            .I(N__22730));
    LocalMux I__3784 (
            .O(N__22730),
            .I(N__22726));
    InMux I__3783 (
            .O(N__22729),
            .I(N__22716));
    Span4Mux_v I__3782 (
            .O(N__22726),
            .I(N__22712));
    InMux I__3781 (
            .O(N__22725),
            .I(N__22707));
    InMux I__3780 (
            .O(N__22724),
            .I(N__22707));
    InMux I__3779 (
            .O(N__22723),
            .I(N__22700));
    InMux I__3778 (
            .O(N__22722),
            .I(N__22700));
    InMux I__3777 (
            .O(N__22721),
            .I(N__22700));
    InMux I__3776 (
            .O(N__22720),
            .I(N__22693));
    CascadeMux I__3775 (
            .O(N__22719),
            .I(N__22688));
    LocalMux I__3774 (
            .O(N__22716),
            .I(N__22681));
    InMux I__3773 (
            .O(N__22715),
            .I(N__22678));
    Span4Mux_v I__3772 (
            .O(N__22712),
            .I(N__22669));
    LocalMux I__3771 (
            .O(N__22707),
            .I(N__22669));
    LocalMux I__3770 (
            .O(N__22700),
            .I(N__22666));
    InMux I__3769 (
            .O(N__22699),
            .I(N__22657));
    InMux I__3768 (
            .O(N__22698),
            .I(N__22657));
    InMux I__3767 (
            .O(N__22697),
            .I(N__22657));
    InMux I__3766 (
            .O(N__22696),
            .I(N__22657));
    LocalMux I__3765 (
            .O(N__22693),
            .I(N__22654));
    InMux I__3764 (
            .O(N__22692),
            .I(N__22645));
    InMux I__3763 (
            .O(N__22691),
            .I(N__22645));
    InMux I__3762 (
            .O(N__22688),
            .I(N__22645));
    InMux I__3761 (
            .O(N__22687),
            .I(N__22645));
    InMux I__3760 (
            .O(N__22686),
            .I(N__22638));
    InMux I__3759 (
            .O(N__22685),
            .I(N__22638));
    InMux I__3758 (
            .O(N__22684),
            .I(N__22638));
    Span4Mux_s1_v I__3757 (
            .O(N__22681),
            .I(N__22635));
    LocalMux I__3756 (
            .O(N__22678),
            .I(N__22632));
    InMux I__3755 (
            .O(N__22677),
            .I(N__22623));
    InMux I__3754 (
            .O(N__22676),
            .I(N__22623));
    InMux I__3753 (
            .O(N__22675),
            .I(N__22623));
    InMux I__3752 (
            .O(N__22674),
            .I(N__22623));
    Span4Mux_s1_v I__3751 (
            .O(N__22669),
            .I(N__22618));
    Span4Mux_h I__3750 (
            .O(N__22666),
            .I(N__22618));
    LocalMux I__3749 (
            .O(N__22657),
            .I(testWordZ0Z_1));
    Odrv4 I__3748 (
            .O(N__22654),
            .I(testWordZ0Z_1));
    LocalMux I__3747 (
            .O(N__22645),
            .I(testWordZ0Z_1));
    LocalMux I__3746 (
            .O(N__22638),
            .I(testWordZ0Z_1));
    Odrv4 I__3745 (
            .O(N__22635),
            .I(testWordZ0Z_1));
    Odrv4 I__3744 (
            .O(N__22632),
            .I(testWordZ0Z_1));
    LocalMux I__3743 (
            .O(N__22623),
            .I(testWordZ0Z_1));
    Odrv4 I__3742 (
            .O(N__22618),
            .I(testWordZ0Z_1));
    CascadeMux I__3741 (
            .O(N__22601),
            .I(N__22591));
    CascadeMux I__3740 (
            .O(N__22600),
            .I(N__22588));
    CascadeMux I__3739 (
            .O(N__22599),
            .I(N__22585));
    CascadeMux I__3738 (
            .O(N__22598),
            .I(N__22578));
    CascadeMux I__3737 (
            .O(N__22597),
            .I(N__22575));
    CascadeMux I__3736 (
            .O(N__22596),
            .I(N__22570));
    CascadeMux I__3735 (
            .O(N__22595),
            .I(N__22566));
    InMux I__3734 (
            .O(N__22594),
            .I(N__22559));
    InMux I__3733 (
            .O(N__22591),
            .I(N__22559));
    InMux I__3732 (
            .O(N__22588),
            .I(N__22559));
    InMux I__3731 (
            .O(N__22585),
            .I(N__22556));
    CascadeMux I__3730 (
            .O(N__22584),
            .I(N__22552));
    CascadeMux I__3729 (
            .O(N__22583),
            .I(N__22549));
    CascadeMux I__3728 (
            .O(N__22582),
            .I(N__22546));
    InMux I__3727 (
            .O(N__22581),
            .I(N__22537));
    InMux I__3726 (
            .O(N__22578),
            .I(N__22537));
    InMux I__3725 (
            .O(N__22575),
            .I(N__22537));
    InMux I__3724 (
            .O(N__22574),
            .I(N__22537));
    InMux I__3723 (
            .O(N__22573),
            .I(N__22530));
    InMux I__3722 (
            .O(N__22570),
            .I(N__22530));
    InMux I__3721 (
            .O(N__22569),
            .I(N__22530));
    InMux I__3720 (
            .O(N__22566),
            .I(N__22527));
    LocalMux I__3719 (
            .O(N__22559),
            .I(N__22520));
    LocalMux I__3718 (
            .O(N__22556),
            .I(N__22520));
    InMux I__3717 (
            .O(N__22555),
            .I(N__22511));
    InMux I__3716 (
            .O(N__22552),
            .I(N__22511));
    InMux I__3715 (
            .O(N__22549),
            .I(N__22511));
    InMux I__3714 (
            .O(N__22546),
            .I(N__22511));
    LocalMux I__3713 (
            .O(N__22537),
            .I(N__22508));
    LocalMux I__3712 (
            .O(N__22530),
            .I(N__22505));
    LocalMux I__3711 (
            .O(N__22527),
            .I(N__22501));
    CascadeMux I__3710 (
            .O(N__22526),
            .I(N__22498));
    CascadeMux I__3709 (
            .O(N__22525),
            .I(N__22494));
    Span4Mux_s3_v I__3708 (
            .O(N__22520),
            .I(N__22489));
    LocalMux I__3707 (
            .O(N__22511),
            .I(N__22482));
    Span4Mux_h I__3706 (
            .O(N__22508),
            .I(N__22482));
    Span4Mux_s1_v I__3705 (
            .O(N__22505),
            .I(N__22482));
    InMux I__3704 (
            .O(N__22504),
            .I(N__22479));
    Span4Mux_h I__3703 (
            .O(N__22501),
            .I(N__22476));
    InMux I__3702 (
            .O(N__22498),
            .I(N__22473));
    InMux I__3701 (
            .O(N__22497),
            .I(N__22468));
    InMux I__3700 (
            .O(N__22494),
            .I(N__22468));
    InMux I__3699 (
            .O(N__22493),
            .I(N__22463));
    InMux I__3698 (
            .O(N__22492),
            .I(N__22463));
    Span4Mux_h I__3697 (
            .O(N__22489),
            .I(N__22460));
    Span4Mux_h I__3696 (
            .O(N__22482),
            .I(N__22457));
    LocalMux I__3695 (
            .O(N__22479),
            .I(testWordZ0Z_4));
    Odrv4 I__3694 (
            .O(N__22476),
            .I(testWordZ0Z_4));
    LocalMux I__3693 (
            .O(N__22473),
            .I(testWordZ0Z_4));
    LocalMux I__3692 (
            .O(N__22468),
            .I(testWordZ0Z_4));
    LocalMux I__3691 (
            .O(N__22463),
            .I(testWordZ0Z_4));
    Odrv4 I__3690 (
            .O(N__22460),
            .I(testWordZ0Z_4));
    Odrv4 I__3689 (
            .O(N__22457),
            .I(testWordZ0Z_4));
    CascadeMux I__3688 (
            .O(N__22442),
            .I(N__22433));
    InMux I__3687 (
            .O(N__22441),
            .I(N__22423));
    InMux I__3686 (
            .O(N__22440),
            .I(N__22423));
    InMux I__3685 (
            .O(N__22439),
            .I(N__22423));
    InMux I__3684 (
            .O(N__22438),
            .I(N__22420));
    InMux I__3683 (
            .O(N__22437),
            .I(N__22410));
    InMux I__3682 (
            .O(N__22436),
            .I(N__22410));
    InMux I__3681 (
            .O(N__22433),
            .I(N__22410));
    InMux I__3680 (
            .O(N__22432),
            .I(N__22410));
    InMux I__3679 (
            .O(N__22431),
            .I(N__22397));
    InMux I__3678 (
            .O(N__22430),
            .I(N__22397));
    LocalMux I__3677 (
            .O(N__22423),
            .I(N__22392));
    LocalMux I__3676 (
            .O(N__22420),
            .I(N__22392));
    InMux I__3675 (
            .O(N__22419),
            .I(N__22389));
    LocalMux I__3674 (
            .O(N__22410),
            .I(N__22382));
    InMux I__3673 (
            .O(N__22409),
            .I(N__22379));
    InMux I__3672 (
            .O(N__22408),
            .I(N__22376));
    InMux I__3671 (
            .O(N__22407),
            .I(N__22373));
    InMux I__3670 (
            .O(N__22406),
            .I(N__22366));
    InMux I__3669 (
            .O(N__22405),
            .I(N__22366));
    InMux I__3668 (
            .O(N__22404),
            .I(N__22366));
    InMux I__3667 (
            .O(N__22403),
            .I(N__22361));
    InMux I__3666 (
            .O(N__22402),
            .I(N__22361));
    LocalMux I__3665 (
            .O(N__22397),
            .I(N__22354));
    Span4Mux_h I__3664 (
            .O(N__22392),
            .I(N__22354));
    LocalMux I__3663 (
            .O(N__22389),
            .I(N__22354));
    InMux I__3662 (
            .O(N__22388),
            .I(N__22345));
    InMux I__3661 (
            .O(N__22387),
            .I(N__22345));
    InMux I__3660 (
            .O(N__22386),
            .I(N__22345));
    InMux I__3659 (
            .O(N__22385),
            .I(N__22345));
    Span12Mux_s1_v I__3658 (
            .O(N__22382),
            .I(N__22342));
    LocalMux I__3657 (
            .O(N__22379),
            .I(testWordZ0Z_2));
    LocalMux I__3656 (
            .O(N__22376),
            .I(testWordZ0Z_2));
    LocalMux I__3655 (
            .O(N__22373),
            .I(testWordZ0Z_2));
    LocalMux I__3654 (
            .O(N__22366),
            .I(testWordZ0Z_2));
    LocalMux I__3653 (
            .O(N__22361),
            .I(testWordZ0Z_2));
    Odrv4 I__3652 (
            .O(N__22354),
            .I(testWordZ0Z_2));
    LocalMux I__3651 (
            .O(N__22345),
            .I(testWordZ0Z_2));
    Odrv12 I__3650 (
            .O(N__22342),
            .I(testWordZ0Z_2));
    CascadeMux I__3649 (
            .O(N__22325),
            .I(N__22316));
    InMux I__3648 (
            .O(N__22324),
            .I(N__22307));
    InMux I__3647 (
            .O(N__22323),
            .I(N__22307));
    InMux I__3646 (
            .O(N__22322),
            .I(N__22307));
    InMux I__3645 (
            .O(N__22321),
            .I(N__22307));
    InMux I__3644 (
            .O(N__22320),
            .I(N__22300));
    InMux I__3643 (
            .O(N__22319),
            .I(N__22300));
    InMux I__3642 (
            .O(N__22316),
            .I(N__22300));
    LocalMux I__3641 (
            .O(N__22307),
            .I(N__22286));
    LocalMux I__3640 (
            .O(N__22300),
            .I(N__22286));
    InMux I__3639 (
            .O(N__22299),
            .I(N__22282));
    CascadeMux I__3638 (
            .O(N__22298),
            .I(N__22277));
    InMux I__3637 (
            .O(N__22297),
            .I(N__22267));
    InMux I__3636 (
            .O(N__22296),
            .I(N__22267));
    InMux I__3635 (
            .O(N__22295),
            .I(N__22267));
    InMux I__3634 (
            .O(N__22294),
            .I(N__22258));
    InMux I__3633 (
            .O(N__22293),
            .I(N__22258));
    InMux I__3632 (
            .O(N__22292),
            .I(N__22258));
    InMux I__3631 (
            .O(N__22291),
            .I(N__22258));
    Span4Mux_s3_v I__3630 (
            .O(N__22286),
            .I(N__22252));
    InMux I__3629 (
            .O(N__22285),
            .I(N__22249));
    LocalMux I__3628 (
            .O(N__22282),
            .I(N__22246));
    InMux I__3627 (
            .O(N__22281),
            .I(N__22241));
    InMux I__3626 (
            .O(N__22280),
            .I(N__22241));
    InMux I__3625 (
            .O(N__22277),
            .I(N__22232));
    InMux I__3624 (
            .O(N__22276),
            .I(N__22232));
    InMux I__3623 (
            .O(N__22275),
            .I(N__22232));
    InMux I__3622 (
            .O(N__22274),
            .I(N__22232));
    LocalMux I__3621 (
            .O(N__22267),
            .I(N__22229));
    LocalMux I__3620 (
            .O(N__22258),
            .I(N__22226));
    InMux I__3619 (
            .O(N__22257),
            .I(N__22219));
    InMux I__3618 (
            .O(N__22256),
            .I(N__22219));
    InMux I__3617 (
            .O(N__22255),
            .I(N__22219));
    IoSpan4Mux I__3616 (
            .O(N__22252),
            .I(N__22216));
    LocalMux I__3615 (
            .O(N__22249),
            .I(N__22213));
    Span4Mux_s1_v I__3614 (
            .O(N__22246),
            .I(N__22204));
    LocalMux I__3613 (
            .O(N__22241),
            .I(N__22204));
    LocalMux I__3612 (
            .O(N__22232),
            .I(N__22204));
    Span4Mux_h I__3611 (
            .O(N__22229),
            .I(N__22204));
    Span4Mux_v I__3610 (
            .O(N__22226),
            .I(N__22200));
    LocalMux I__3609 (
            .O(N__22219),
            .I(N__22197));
    Span4Mux_s0_h I__3608 (
            .O(N__22216),
            .I(N__22192));
    Span4Mux_h I__3607 (
            .O(N__22213),
            .I(N__22192));
    Span4Mux_h I__3606 (
            .O(N__22204),
            .I(N__22189));
    InMux I__3605 (
            .O(N__22203),
            .I(N__22186));
    Span4Mux_h I__3604 (
            .O(N__22200),
            .I(N__22181));
    Span4Mux_v I__3603 (
            .O(N__22197),
            .I(N__22181));
    Span4Mux_v I__3602 (
            .O(N__22192),
            .I(N__22178));
    Span4Mux_v I__3601 (
            .O(N__22189),
            .I(N__22175));
    LocalMux I__3600 (
            .O(N__22186),
            .I(testWordZ0Z_3));
    Odrv4 I__3599 (
            .O(N__22181),
            .I(testWordZ0Z_3));
    Odrv4 I__3598 (
            .O(N__22178),
            .I(testWordZ0Z_3));
    Odrv4 I__3597 (
            .O(N__22175),
            .I(testWordZ0Z_3));
    CascadeMux I__3596 (
            .O(N__22166),
            .I(\ALU.N_469_cascade_ ));
    InMux I__3595 (
            .O(N__22163),
            .I(N__22160));
    LocalMux I__3594 (
            .O(N__22160),
            .I(\ALU.N_473 ));
    CascadeMux I__3593 (
            .O(N__22157),
            .I(\ALU.rshift_15_ns_1_1_cascade_ ));
    InMux I__3592 (
            .O(N__22154),
            .I(N__22151));
    LocalMux I__3591 (
            .O(N__22151),
            .I(N__22148));
    Span4Mux_h I__3590 (
            .O(N__22148),
            .I(N__22145));
    Span4Mux_h I__3589 (
            .O(N__22145),
            .I(N__22142));
    Odrv4 I__3588 (
            .O(N__22142),
            .I(N_305_0));
    CEMux I__3587 (
            .O(N__22139),
            .I(N__22134));
    InMux I__3586 (
            .O(N__22138),
            .I(N__22131));
    InMux I__3585 (
            .O(N__22137),
            .I(N__22128));
    LocalMux I__3584 (
            .O(N__22134),
            .I(N__22125));
    LocalMux I__3583 (
            .O(N__22131),
            .I(N__22121));
    LocalMux I__3582 (
            .O(N__22128),
            .I(N__22118));
    Span4Mux_h I__3581 (
            .O(N__22125),
            .I(N__22115));
    InMux I__3580 (
            .O(N__22124),
            .I(N__22112));
    Span4Mux_h I__3579 (
            .O(N__22121),
            .I(N__22107));
    Span4Mux_s2_v I__3578 (
            .O(N__22118),
            .I(N__22107));
    Odrv4 I__3577 (
            .O(N__22115),
            .I(\CONTROL.aluParams_cnvZ0Z_0 ));
    LocalMux I__3576 (
            .O(N__22112),
            .I(\CONTROL.aluParams_cnvZ0Z_0 ));
    Odrv4 I__3575 (
            .O(N__22107),
            .I(\CONTROL.aluParams_cnvZ0Z_0 ));
    InMux I__3574 (
            .O(N__22100),
            .I(N__22097));
    LocalMux I__3573 (
            .O(N__22097),
            .I(\ALU.a4_b_4 ));
    InMux I__3572 (
            .O(N__22094),
            .I(N__22091));
    LocalMux I__3571 (
            .O(N__22091),
            .I(\ALU.a3_b_5 ));
    CascadeMux I__3570 (
            .O(N__22088),
            .I(\ALU.a4_b_4_cascade_ ));
    InMux I__3569 (
            .O(N__22085),
            .I(N__22082));
    LocalMux I__3568 (
            .O(N__22082),
            .I(N__22079));
    Span4Mux_h I__3567 (
            .O(N__22079),
            .I(N__22076));
    Odrv4 I__3566 (
            .O(N__22076),
            .I(\ALU.madd_98 ));
    CascadeMux I__3565 (
            .O(N__22073),
            .I(N__22069));
    InMux I__3564 (
            .O(N__22072),
            .I(N__22061));
    InMux I__3563 (
            .O(N__22069),
            .I(N__22058));
    InMux I__3562 (
            .O(N__22068),
            .I(N__22054));
    InMux I__3561 (
            .O(N__22067),
            .I(N__22049));
    InMux I__3560 (
            .O(N__22066),
            .I(N__22049));
    InMux I__3559 (
            .O(N__22065),
            .I(N__22044));
    InMux I__3558 (
            .O(N__22064),
            .I(N__22041));
    LocalMux I__3557 (
            .O(N__22061),
            .I(N__22036));
    LocalMux I__3556 (
            .O(N__22058),
            .I(N__22036));
    InMux I__3555 (
            .O(N__22057),
            .I(N__22033));
    LocalMux I__3554 (
            .O(N__22054),
            .I(N__22030));
    LocalMux I__3553 (
            .O(N__22049),
            .I(N__22027));
    InMux I__3552 (
            .O(N__22048),
            .I(N__22022));
    InMux I__3551 (
            .O(N__22047),
            .I(N__22022));
    LocalMux I__3550 (
            .O(N__22044),
            .I(N__22019));
    LocalMux I__3549 (
            .O(N__22041),
            .I(N__22014));
    Span4Mux_v I__3548 (
            .O(N__22036),
            .I(N__22014));
    LocalMux I__3547 (
            .O(N__22033),
            .I(N__22007));
    Span4Mux_v I__3546 (
            .O(N__22030),
            .I(N__22007));
    Span4Mux_h I__3545 (
            .O(N__22027),
            .I(N__22007));
    LocalMux I__3544 (
            .O(N__22022),
            .I(N__22004));
    Span4Mux_v I__3543 (
            .O(N__22019),
            .I(N__21997));
    Span4Mux_v I__3542 (
            .O(N__22014),
            .I(N__21997));
    Span4Mux_v I__3541 (
            .O(N__22007),
            .I(N__21992));
    Span4Mux_h I__3540 (
            .O(N__22004),
            .I(N__21992));
    InMux I__3539 (
            .O(N__22003),
            .I(N__21987));
    InMux I__3538 (
            .O(N__22002),
            .I(N__21987));
    Odrv4 I__3537 (
            .O(N__21997),
            .I(\ALU.N_207_0 ));
    Odrv4 I__3536 (
            .O(N__21992),
            .I(\ALU.N_207_0 ));
    LocalMux I__3535 (
            .O(N__21987),
            .I(\ALU.N_207_0 ));
    CascadeMux I__3534 (
            .O(N__21980),
            .I(\ALU.madd_98_cascade_ ));
    InMux I__3533 (
            .O(N__21977),
            .I(N__21974));
    LocalMux I__3532 (
            .O(N__21974),
            .I(N__21970));
    InMux I__3531 (
            .O(N__21973),
            .I(N__21967));
    Span4Mux_s3_h I__3530 (
            .O(N__21970),
            .I(N__21964));
    LocalMux I__3529 (
            .O(N__21967),
            .I(N__21961));
    Sp12to4 I__3528 (
            .O(N__21964),
            .I(N__21958));
    Span4Mux_h I__3527 (
            .O(N__21961),
            .I(N__21955));
    Odrv12 I__3526 (
            .O(N__21958),
            .I(\ALU.madd_93 ));
    Odrv4 I__3525 (
            .O(N__21955),
            .I(\ALU.madd_93 ));
    InMux I__3524 (
            .O(N__21950),
            .I(N__21941));
    InMux I__3523 (
            .O(N__21949),
            .I(N__21941));
    InMux I__3522 (
            .O(N__21948),
            .I(N__21941));
    LocalMux I__3521 (
            .O(N__21941),
            .I(\ALU.madd_139 ));
    InMux I__3520 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__3519 (
            .O(N__21935),
            .I(N__21931));
    CascadeMux I__3518 (
            .O(N__21934),
            .I(N__21928));
    Span4Mux_v I__3517 (
            .O(N__21931),
            .I(N__21925));
    InMux I__3516 (
            .O(N__21928),
            .I(N__21922));
    Span4Mux_h I__3515 (
            .O(N__21925),
            .I(N__21917));
    LocalMux I__3514 (
            .O(N__21922),
            .I(N__21917));
    Span4Mux_h I__3513 (
            .O(N__21917),
            .I(N__21914));
    Span4Mux_h I__3512 (
            .O(N__21914),
            .I(N__21911));
    Span4Mux_h I__3511 (
            .O(N__21911),
            .I(N__21908));
    Span4Mux_h I__3510 (
            .O(N__21908),
            .I(N__21905));
    Odrv4 I__3509 (
            .O(N__21905),
            .I(RX_c));
    InMux I__3508 (
            .O(N__21902),
            .I(N__21899));
    LocalMux I__3507 (
            .O(N__21899),
            .I(N__21896));
    Span4Mux_v I__3506 (
            .O(N__21896),
            .I(N__21892));
    InMux I__3505 (
            .O(N__21895),
            .I(N__21889));
    Span4Mux_v I__3504 (
            .O(N__21892),
            .I(N__21884));
    LocalMux I__3503 (
            .O(N__21889),
            .I(N__21880));
    InMux I__3502 (
            .O(N__21888),
            .I(N__21875));
    InMux I__3501 (
            .O(N__21887),
            .I(N__21875));
    Span4Mux_h I__3500 (
            .O(N__21884),
            .I(N__21872));
    InMux I__3499 (
            .O(N__21883),
            .I(N__21869));
    Odrv4 I__3498 (
            .O(N__21880),
            .I(RXready));
    LocalMux I__3497 (
            .O(N__21875),
            .I(RXready));
    Odrv4 I__3496 (
            .O(N__21872),
            .I(RXready));
    LocalMux I__3495 (
            .O(N__21869),
            .I(RXready));
    CascadeMux I__3494 (
            .O(N__21860),
            .I(N__21856));
    CascadeMux I__3493 (
            .O(N__21859),
            .I(N__21853));
    InMux I__3492 (
            .O(N__21856),
            .I(N__21850));
    InMux I__3491 (
            .O(N__21853),
            .I(N__21847));
    LocalMux I__3490 (
            .O(N__21850),
            .I(N__21843));
    LocalMux I__3489 (
            .O(N__21847),
            .I(N__21840));
    InMux I__3488 (
            .O(N__21846),
            .I(N__21837));
    Span12Mux_s3_v I__3487 (
            .O(N__21843),
            .I(N__21834));
    Span4Mux_h I__3486 (
            .O(N__21840),
            .I(N__21831));
    LocalMux I__3485 (
            .O(N__21837),
            .I(ctrlOut_1));
    Odrv12 I__3484 (
            .O(N__21834),
            .I(ctrlOut_1));
    Odrv4 I__3483 (
            .O(N__21831),
            .I(ctrlOut_1));
    CascadeMux I__3482 (
            .O(N__21824),
            .I(\ALU.N_41_0_0_cascade_ ));
    InMux I__3481 (
            .O(N__21821),
            .I(N__21818));
    LocalMux I__3480 (
            .O(N__21818),
            .I(\ALU.rshift_3_ns_1_5 ));
    CascadeMux I__3479 (
            .O(N__21815),
            .I(\ALU.N_752_cascade_ ));
    CascadeMux I__3478 (
            .O(N__21812),
            .I(\ALU.dout_3_ns_1_5_cascade_ ));
    InMux I__3477 (
            .O(N__21809),
            .I(N__21806));
    LocalMux I__3476 (
            .O(N__21806),
            .I(\ALU.N_704 ));
    CascadeMux I__3475 (
            .O(N__21803),
            .I(\ALU.un2_addsub_axb_4_cascade_ ));
    CascadeMux I__3474 (
            .O(N__21800),
            .I(N__21797));
    InMux I__3473 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__3472 (
            .O(N__21794),
            .I(N__21791));
    Odrv12 I__3471 (
            .O(N__21791),
            .I(\ALU.d_RNI312TBZ0Z_4 ));
    InMux I__3470 (
            .O(N__21788),
            .I(N__21781));
    InMux I__3469 (
            .O(N__21787),
            .I(N__21776));
    InMux I__3468 (
            .O(N__21786),
            .I(N__21776));
    InMux I__3467 (
            .O(N__21785),
            .I(N__21773));
    InMux I__3466 (
            .O(N__21784),
            .I(N__21770));
    LocalMux I__3465 (
            .O(N__21781),
            .I(N__21767));
    LocalMux I__3464 (
            .O(N__21776),
            .I(N__21762));
    LocalMux I__3463 (
            .O(N__21773),
            .I(N__21759));
    LocalMux I__3462 (
            .O(N__21770),
            .I(N__21754));
    Span4Mux_v I__3461 (
            .O(N__21767),
            .I(N__21754));
    InMux I__3460 (
            .O(N__21766),
            .I(N__21749));
    InMux I__3459 (
            .O(N__21765),
            .I(N__21749));
    Span4Mux_v I__3458 (
            .O(N__21762),
            .I(N__21746));
    Span4Mux_h I__3457 (
            .O(N__21759),
            .I(N__21739));
    Span4Mux_h I__3456 (
            .O(N__21754),
            .I(N__21739));
    LocalMux I__3455 (
            .O(N__21749),
            .I(N__21739));
    Span4Mux_v I__3454 (
            .O(N__21746),
            .I(N__21736));
    Span4Mux_v I__3453 (
            .O(N__21739),
            .I(N__21733));
    Odrv4 I__3452 (
            .O(N__21736),
            .I(\ALU.N_223_0 ));
    Odrv4 I__3451 (
            .O(N__21733),
            .I(\ALU.N_223_0 ));
    InMux I__3450 (
            .O(N__21728),
            .I(N__21725));
    LocalMux I__3449 (
            .O(N__21725),
            .I(N__21718));
    InMux I__3448 (
            .O(N__21724),
            .I(N__21715));
    InMux I__3447 (
            .O(N__21723),
            .I(N__21710));
    InMux I__3446 (
            .O(N__21722),
            .I(N__21710));
    InMux I__3445 (
            .O(N__21721),
            .I(N__21707));
    Span4Mux_v I__3444 (
            .O(N__21718),
            .I(N__21704));
    LocalMux I__3443 (
            .O(N__21715),
            .I(N__21701));
    LocalMux I__3442 (
            .O(N__21710),
            .I(N__21696));
    LocalMux I__3441 (
            .O(N__21707),
            .I(N__21693));
    Span4Mux_v I__3440 (
            .O(N__21704),
            .I(N__21688));
    Span4Mux_v I__3439 (
            .O(N__21701),
            .I(N__21688));
    InMux I__3438 (
            .O(N__21700),
            .I(N__21683));
    InMux I__3437 (
            .O(N__21699),
            .I(N__21683));
    Odrv4 I__3436 (
            .O(N__21696),
            .I(\ALU.operand2_5 ));
    Odrv12 I__3435 (
            .O(N__21693),
            .I(\ALU.operand2_5 ));
    Odrv4 I__3434 (
            .O(N__21688),
            .I(\ALU.operand2_5 ));
    LocalMux I__3433 (
            .O(N__21683),
            .I(\ALU.operand2_5 ));
    CascadeMux I__3432 (
            .O(N__21674),
            .I(\ALU.a3_b_5_cascade_ ));
    InMux I__3431 (
            .O(N__21671),
            .I(N__21665));
    InMux I__3430 (
            .O(N__21670),
            .I(N__21665));
    LocalMux I__3429 (
            .O(N__21665),
            .I(N__21662));
    Odrv12 I__3428 (
            .O(N__21662),
            .I(\ALU.madd_94 ));
    CascadeMux I__3427 (
            .O(N__21659),
            .I(\ALU.g_RNIT0COZ0Z_1_cascade_ ));
    CascadeMux I__3426 (
            .O(N__21656),
            .I(\ALU.operand2_7_ns_1_1_cascade_ ));
    InMux I__3425 (
            .O(N__21653),
            .I(N__21650));
    LocalMux I__3424 (
            .O(N__21650),
            .I(N__21647));
    Odrv4 I__3423 (
            .O(N__21647),
            .I(\ALU.e_RNIPKVJZ0Z_1 ));
    InMux I__3422 (
            .O(N__21644),
            .I(N__21641));
    LocalMux I__3421 (
            .O(N__21641),
            .I(N__21638));
    Odrv4 I__3420 (
            .O(N__21638),
            .I(\ALU.madd_4 ));
    InMux I__3419 (
            .O(N__21635),
            .I(N__21632));
    LocalMux I__3418 (
            .O(N__21632),
            .I(N__21629));
    Odrv4 I__3417 (
            .O(N__21629),
            .I(\ALU.madd_12_0_tz ));
    CascadeMux I__3416 (
            .O(N__21626),
            .I(\ALU.dout_6_ns_1_15_cascade_ ));
    CascadeMux I__3415 (
            .O(N__21623),
            .I(\ALU.N_747_cascade_ ));
    CascadeMux I__3414 (
            .O(N__21620),
            .I(\ALU.aluOut_0_cascade_ ));
    InMux I__3413 (
            .O(N__21617),
            .I(N__21614));
    LocalMux I__3412 (
            .O(N__21614),
            .I(N__21611));
    Span4Mux_s2_h I__3411 (
            .O(N__21611),
            .I(N__21608));
    Span4Mux_v I__3410 (
            .O(N__21608),
            .I(N__21605));
    Span4Mux_h I__3409 (
            .O(N__21605),
            .I(N__21602));
    Odrv4 I__3408 (
            .O(N__21602),
            .I(\ALU.g0_0_0_N_2L1 ));
    InMux I__3407 (
            .O(N__21599),
            .I(N__21596));
    LocalMux I__3406 (
            .O(N__21596),
            .I(\ALU.dout_3_ns_1_7 ));
    CascadeMux I__3405 (
            .O(N__21593),
            .I(N__21590));
    InMux I__3404 (
            .O(N__21590),
            .I(N__21587));
    LocalMux I__3403 (
            .O(N__21587),
            .I(N__21584));
    Odrv12 I__3402 (
            .O(N__21584),
            .I(\ALU.a_15_m5_0 ));
    CascadeMux I__3401 (
            .O(N__21581),
            .I(\ALU.d_RNI9BO713Z0Z_0_cascade_ ));
    CascadeMux I__3400 (
            .O(N__21578),
            .I(\ALU.operand2_7_ns_1_0_cascade_ ));
    InMux I__3399 (
            .O(N__21575),
            .I(N__21572));
    LocalMux I__3398 (
            .O(N__21572),
            .I(N__21569));
    Span4Mux_h I__3397 (
            .O(N__21569),
            .I(N__21565));
    InMux I__3396 (
            .O(N__21568),
            .I(N__21560));
    Span4Mux_v I__3395 (
            .O(N__21565),
            .I(N__21557));
    InMux I__3394 (
            .O(N__21564),
            .I(N__21554));
    InMux I__3393 (
            .O(N__21563),
            .I(N__21551));
    LocalMux I__3392 (
            .O(N__21560),
            .I(N__21546));
    Span4Mux_v I__3391 (
            .O(N__21557),
            .I(N__21546));
    LocalMux I__3390 (
            .O(N__21554),
            .I(ctrlOut_0));
    LocalMux I__3389 (
            .O(N__21551),
            .I(ctrlOut_0));
    Odrv4 I__3388 (
            .O(N__21546),
            .I(ctrlOut_0));
    CascadeMux I__3387 (
            .O(N__21539),
            .I(\ALU.operand2_0_cascade_ ));
    InMux I__3386 (
            .O(N__21536),
            .I(N__21532));
    InMux I__3385 (
            .O(N__21535),
            .I(N__21529));
    LocalMux I__3384 (
            .O(N__21532),
            .I(\ALU.hZ0Z_0 ));
    LocalMux I__3383 (
            .O(N__21529),
            .I(\ALU.hZ0Z_0 ));
    InMux I__3382 (
            .O(N__21524),
            .I(N__21521));
    LocalMux I__3381 (
            .O(N__21521),
            .I(\ALU.d_RNIE4R7Z0Z_0 ));
    InMux I__3380 (
            .O(N__21518),
            .I(N__21515));
    LocalMux I__3379 (
            .O(N__21515),
            .I(\ALU.g0_7_a3_0Z0Z_0 ));
    CascadeMux I__3378 (
            .O(N__21512),
            .I(\ALU.N_8_1_cascade_ ));
    InMux I__3377 (
            .O(N__21509),
            .I(N__21506));
    LocalMux I__3376 (
            .O(N__21506),
            .I(\ALU.g0_2Z0Z_1 ));
    CascadeMux I__3375 (
            .O(N__21503),
            .I(\ALU.g0_7_m4_0_1_cascade_ ));
    InMux I__3374 (
            .O(N__21500),
            .I(N__21497));
    LocalMux I__3373 (
            .O(N__21497),
            .I(\ALU.N_9_2 ));
    CascadeMux I__3372 (
            .O(N__21494),
            .I(\ALU.dout_3_ns_1_0_cascade_ ));
    CascadeMux I__3371 (
            .O(N__21491),
            .I(\ALU.dout_6_ns_1_0_cascade_ ));
    InMux I__3370 (
            .O(N__21488),
            .I(N__21481));
    CascadeMux I__3369 (
            .O(N__21487),
            .I(N__21478));
    CascadeMux I__3368 (
            .O(N__21486),
            .I(N__21475));
    CascadeMux I__3367 (
            .O(N__21485),
            .I(N__21472));
    InMux I__3366 (
            .O(N__21484),
            .I(N__21466));
    LocalMux I__3365 (
            .O(N__21481),
            .I(N__21463));
    InMux I__3364 (
            .O(N__21478),
            .I(N__21460));
    InMux I__3363 (
            .O(N__21475),
            .I(N__21457));
    InMux I__3362 (
            .O(N__21472),
            .I(N__21454));
    InMux I__3361 (
            .O(N__21471),
            .I(N__21451));
    CascadeMux I__3360 (
            .O(N__21470),
            .I(N__21448));
    CascadeMux I__3359 (
            .O(N__21469),
            .I(N__21445));
    LocalMux I__3358 (
            .O(N__21466),
            .I(N__21441));
    Span4Mux_v I__3357 (
            .O(N__21463),
            .I(N__21438));
    LocalMux I__3356 (
            .O(N__21460),
            .I(N__21431));
    LocalMux I__3355 (
            .O(N__21457),
            .I(N__21431));
    LocalMux I__3354 (
            .O(N__21454),
            .I(N__21431));
    LocalMux I__3353 (
            .O(N__21451),
            .I(N__21428));
    InMux I__3352 (
            .O(N__21448),
            .I(N__21421));
    InMux I__3351 (
            .O(N__21445),
            .I(N__21421));
    InMux I__3350 (
            .O(N__21444),
            .I(N__21421));
    Span4Mux_v I__3349 (
            .O(N__21441),
            .I(N__21416));
    Span4Mux_h I__3348 (
            .O(N__21438),
            .I(N__21416));
    Span4Mux_v I__3347 (
            .O(N__21431),
            .I(N__21413));
    Odrv12 I__3346 (
            .O(N__21428),
            .I(\ALU.N_201_0 ));
    LocalMux I__3345 (
            .O(N__21421),
            .I(\ALU.N_201_0 ));
    Odrv4 I__3344 (
            .O(N__21416),
            .I(\ALU.N_201_0 ));
    Odrv4 I__3343 (
            .O(N__21413),
            .I(\ALU.N_201_0 ));
    CascadeMux I__3342 (
            .O(N__21404),
            .I(N__21401));
    InMux I__3341 (
            .O(N__21401),
            .I(N__21398));
    LocalMux I__3340 (
            .O(N__21398),
            .I(N__21395));
    Span4Mux_h I__3339 (
            .O(N__21395),
            .I(N__21392));
    Span4Mux_v I__3338 (
            .O(N__21392),
            .I(N__21389));
    Odrv4 I__3337 (
            .O(N__21389),
            .I(\ALU.d_RNIQ74VBZ0Z_8 ));
    InMux I__3336 (
            .O(N__21386),
            .I(bfn_6_10_0_));
    CascadeMux I__3335 (
            .O(N__21383),
            .I(N__21380));
    InMux I__3334 (
            .O(N__21380),
            .I(N__21377));
    LocalMux I__3333 (
            .O(N__21377),
            .I(N__21374));
    Span12Mux_h I__3332 (
            .O(N__21374),
            .I(N__21371));
    Odrv12 I__3331 (
            .O(N__21371),
            .I(\ALU.d_RNI6B7KDZ0Z_9 ));
    InMux I__3330 (
            .O(N__21368),
            .I(\ALU.un2_addsub_cry_8 ));
    CascadeMux I__3329 (
            .O(N__21365),
            .I(N__21362));
    InMux I__3328 (
            .O(N__21362),
            .I(N__21359));
    LocalMux I__3327 (
            .O(N__21359),
            .I(N__21356));
    Span4Mux_h I__3326 (
            .O(N__21356),
            .I(N__21353));
    Span4Mux_h I__3325 (
            .O(N__21353),
            .I(N__21350));
    Odrv4 I__3324 (
            .O(N__21350),
            .I(\ALU.N_192_0_i ));
    InMux I__3323 (
            .O(N__21347),
            .I(\ALU.un2_addsub_cry_9 ));
    InMux I__3322 (
            .O(N__21344),
            .I(\ALU.un2_addsub_cry_10 ));
    CascadeMux I__3321 (
            .O(N__21341),
            .I(N__21338));
    InMux I__3320 (
            .O(N__21338),
            .I(N__21335));
    LocalMux I__3319 (
            .O(N__21335),
            .I(N__21332));
    Span4Mux_h I__3318 (
            .O(N__21332),
            .I(N__21329));
    Span4Mux_h I__3317 (
            .O(N__21329),
            .I(N__21326));
    Span4Mux_v I__3316 (
            .O(N__21326),
            .I(N__21323));
    Odrv4 I__3315 (
            .O(N__21323),
            .I(\ALU.N_180_0_i ));
    InMux I__3314 (
            .O(N__21320),
            .I(\ALU.un2_addsub_cry_11 ));
    InMux I__3313 (
            .O(N__21317),
            .I(\ALU.un2_addsub_cry_12 ));
    InMux I__3312 (
            .O(N__21314),
            .I(N__21308));
    InMux I__3311 (
            .O(N__21313),
            .I(N__21305));
    InMux I__3310 (
            .O(N__21312),
            .I(N__21301));
    InMux I__3309 (
            .O(N__21311),
            .I(N__21298));
    LocalMux I__3308 (
            .O(N__21308),
            .I(N__21291));
    LocalMux I__3307 (
            .O(N__21305),
            .I(N__21291));
    InMux I__3306 (
            .O(N__21304),
            .I(N__21288));
    LocalMux I__3305 (
            .O(N__21301),
            .I(N__21285));
    LocalMux I__3304 (
            .O(N__21298),
            .I(N__21282));
    InMux I__3303 (
            .O(N__21297),
            .I(N__21277));
    InMux I__3302 (
            .O(N__21296),
            .I(N__21277));
    Span4Mux_v I__3301 (
            .O(N__21291),
            .I(N__21274));
    LocalMux I__3300 (
            .O(N__21288),
            .I(\ALU.N_171_0 ));
    Odrv4 I__3299 (
            .O(N__21285),
            .I(\ALU.N_171_0 ));
    Odrv4 I__3298 (
            .O(N__21282),
            .I(\ALU.N_171_0 ));
    LocalMux I__3297 (
            .O(N__21277),
            .I(\ALU.N_171_0 ));
    Odrv4 I__3296 (
            .O(N__21274),
            .I(\ALU.N_171_0 ));
    CascadeMux I__3295 (
            .O(N__21263),
            .I(N__21260));
    InMux I__3294 (
            .O(N__21260),
            .I(N__21257));
    LocalMux I__3293 (
            .O(N__21257),
            .I(N__21254));
    Span4Mux_h I__3292 (
            .O(N__21254),
            .I(N__21251));
    Span4Mux_v I__3291 (
            .O(N__21251),
            .I(N__21248));
    Odrv4 I__3290 (
            .O(N__21248),
            .I(\ALU.d_RNI1M3JEZ0Z_14 ));
    InMux I__3289 (
            .O(N__21245),
            .I(\ALU.un2_addsub_cry_13 ));
    InMux I__3288 (
            .O(N__21242),
            .I(\ALU.un2_addsub_cry_14 ));
    CascadeMux I__3287 (
            .O(N__21239),
            .I(N__21236));
    InMux I__3286 (
            .O(N__21236),
            .I(N__21227));
    InMux I__3285 (
            .O(N__21235),
            .I(N__21227));
    InMux I__3284 (
            .O(N__21234),
            .I(N__21227));
    LocalMux I__3283 (
            .O(N__21227),
            .I(N__21224));
    Span4Mux_v I__3282 (
            .O(N__21224),
            .I(N__21221));
    Span4Mux_h I__3281 (
            .O(N__21221),
            .I(N__21218));
    Odrv4 I__3280 (
            .O(N__21218),
            .I(\ALU.a0_b_11 ));
    InMux I__3279 (
            .O(N__21215),
            .I(\ALU.un2_addsub_cry_0 ));
    InMux I__3278 (
            .O(N__21212),
            .I(N__21209));
    LocalMux I__3277 (
            .O(N__21209),
            .I(N__21206));
    Sp12to4 I__3276 (
            .O(N__21206),
            .I(N__21203));
    Span12Mux_s4_h I__3275 (
            .O(N__21203),
            .I(N__21200));
    Odrv12 I__3274 (
            .O(N__21200),
            .I(\ALU.d_RNIEDJEAZ0Z_2 ));
    CascadeMux I__3273 (
            .O(N__21197),
            .I(N__21194));
    InMux I__3272 (
            .O(N__21194),
            .I(N__21191));
    LocalMux I__3271 (
            .O(N__21191),
            .I(N__21188));
    Span4Mux_h I__3270 (
            .O(N__21188),
            .I(N__21185));
    Span4Mux_h I__3269 (
            .O(N__21185),
            .I(N__21182));
    Odrv4 I__3268 (
            .O(N__21182),
            .I(\ALU.N_240_0_i ));
    InMux I__3267 (
            .O(N__21179),
            .I(\ALU.un2_addsub_cry_1 ));
    InMux I__3266 (
            .O(N__21176),
            .I(\ALU.un2_addsub_cry_2 ));
    InMux I__3265 (
            .O(N__21173),
            .I(\ALU.un2_addsub_cry_3 ));
    CascadeMux I__3264 (
            .O(N__21170),
            .I(N__21167));
    InMux I__3263 (
            .O(N__21167),
            .I(N__21164));
    LocalMux I__3262 (
            .O(N__21164),
            .I(N__21161));
    Span4Mux_h I__3261 (
            .O(N__21161),
            .I(N__21158));
    Span4Mux_v I__3260 (
            .O(N__21158),
            .I(N__21155));
    Odrv4 I__3259 (
            .O(N__21155),
            .I(\ALU.d_RNIVR3QAZ0Z_5 ));
    InMux I__3258 (
            .O(N__21152),
            .I(\ALU.un2_addsub_cry_4 ));
    CascadeMux I__3257 (
            .O(N__21149),
            .I(N__21146));
    InMux I__3256 (
            .O(N__21146),
            .I(N__21143));
    LocalMux I__3255 (
            .O(N__21143),
            .I(N__21140));
    Span4Mux_v I__3254 (
            .O(N__21140),
            .I(N__21137));
    Span4Mux_v I__3253 (
            .O(N__21137),
            .I(N__21134));
    Span4Mux_h I__3252 (
            .O(N__21134),
            .I(N__21131));
    Odrv4 I__3251 (
            .O(N__21131),
            .I(\ALU.d_RNIGLK5BZ0Z_6 ));
    InMux I__3250 (
            .O(N__21128),
            .I(\ALU.un2_addsub_cry_5 ));
    CascadeMux I__3249 (
            .O(N__21125),
            .I(N__21122));
    InMux I__3248 (
            .O(N__21122),
            .I(N__21119));
    LocalMux I__3247 (
            .O(N__21119),
            .I(N__21116));
    Span4Mux_h I__3246 (
            .O(N__21116),
            .I(N__21113));
    Span4Mux_h I__3245 (
            .O(N__21113),
            .I(N__21110));
    Span4Mux_s1_h I__3244 (
            .O(N__21110),
            .I(N__21107));
    Span4Mux_v I__3243 (
            .O(N__21107),
            .I(N__21104));
    Odrv4 I__3242 (
            .O(N__21104),
            .I(\ALU.d_RNITAM9DZ0Z_7 ));
    InMux I__3241 (
            .O(N__21101),
            .I(\ALU.un2_addsub_cry_6 ));
    InMux I__3240 (
            .O(N__21098),
            .I(N__21090));
    InMux I__3239 (
            .O(N__21097),
            .I(N__21086));
    InMux I__3238 (
            .O(N__21096),
            .I(N__21083));
    InMux I__3237 (
            .O(N__21095),
            .I(N__21076));
    InMux I__3236 (
            .O(N__21094),
            .I(N__21076));
    InMux I__3235 (
            .O(N__21093),
            .I(N__21076));
    LocalMux I__3234 (
            .O(N__21090),
            .I(N__21073));
    InMux I__3233 (
            .O(N__21089),
            .I(N__21070));
    LocalMux I__3232 (
            .O(N__21086),
            .I(N__21067));
    LocalMux I__3231 (
            .O(N__21083),
            .I(N__21064));
    LocalMux I__3230 (
            .O(N__21076),
            .I(N__21061));
    Span4Mux_v I__3229 (
            .O(N__21073),
            .I(N__21058));
    LocalMux I__3228 (
            .O(N__21070),
            .I(N__21054));
    Span4Mux_v I__3227 (
            .O(N__21067),
            .I(N__21049));
    Span4Mux_v I__3226 (
            .O(N__21064),
            .I(N__21049));
    Span4Mux_h I__3225 (
            .O(N__21061),
            .I(N__21044));
    Span4Mux_h I__3224 (
            .O(N__21058),
            .I(N__21044));
    InMux I__3223 (
            .O(N__21057),
            .I(N__21041));
    Odrv12 I__3222 (
            .O(N__21054),
            .I(\ALU.N_205_0 ));
    Odrv4 I__3221 (
            .O(N__21049),
            .I(\ALU.N_205_0 ));
    Odrv4 I__3220 (
            .O(N__21044),
            .I(\ALU.N_205_0 ));
    LocalMux I__3219 (
            .O(N__21041),
            .I(\ALU.N_205_0 ));
    CascadeMux I__3218 (
            .O(N__21032),
            .I(\ALU.operand2_9_cascade_ ));
    CascadeMux I__3217 (
            .O(N__21029),
            .I(\ALU.a_15_m2_ns_1Z0Z_9_cascade_ ));
    CascadeMux I__3216 (
            .O(N__21026),
            .I(\ALU.d_RNIO7LUZ0Z_13_cascade_ ));
    CascadeMux I__3215 (
            .O(N__21023),
            .I(\ALU.operand2_13_cascade_ ));
    CascadeMux I__3214 (
            .O(N__21020),
            .I(\ALU.N_177_0_cascade_ ));
    InMux I__3213 (
            .O(N__21017),
            .I(N__21014));
    LocalMux I__3212 (
            .O(N__21014),
            .I(N__21011));
    Odrv12 I__3211 (
            .O(N__21011),
            .I(\ALU.madd_484_3 ));
    InMux I__3210 (
            .O(N__21008),
            .I(N__21005));
    LocalMux I__3209 (
            .O(N__21005),
            .I(N__21002));
    Span4Mux_v I__3208 (
            .O(N__21002),
            .I(N__20999));
    Odrv4 I__3207 (
            .O(N__20999),
            .I(\ALU.madd_484_1 ));
    CascadeMux I__3206 (
            .O(N__20996),
            .I(\ALU.madd_484_2_cascade_ ));
    InMux I__3205 (
            .O(N__20993),
            .I(N__20990));
    LocalMux I__3204 (
            .O(N__20990),
            .I(N__20987));
    Odrv4 I__3203 (
            .O(N__20987),
            .I(\ALU.madd_484_0 ));
    InMux I__3202 (
            .O(N__20984),
            .I(N__20981));
    LocalMux I__3201 (
            .O(N__20981),
            .I(N__20978));
    Odrv4 I__3200 (
            .O(N__20978),
            .I(\ALU.madd_484_12 ));
    CascadeMux I__3199 (
            .O(N__20975),
            .I(\ALU.m270_nsZ0Z_1_cascade_ ));
    CascadeMux I__3198 (
            .O(N__20972),
            .I(N__20967));
    CascadeMux I__3197 (
            .O(N__20971),
            .I(N__20963));
    CascadeMux I__3196 (
            .O(N__20970),
            .I(N__20960));
    InMux I__3195 (
            .O(N__20967),
            .I(N__20957));
    InMux I__3194 (
            .O(N__20966),
            .I(N__20950));
    InMux I__3193 (
            .O(N__20963),
            .I(N__20950));
    InMux I__3192 (
            .O(N__20960),
            .I(N__20950));
    LocalMux I__3191 (
            .O(N__20957),
            .I(ctrlOut_12));
    LocalMux I__3190 (
            .O(N__20950),
            .I(ctrlOut_12));
    CascadeMux I__3189 (
            .O(N__20945),
            .I(N__20941));
    InMux I__3188 (
            .O(N__20944),
            .I(N__20937));
    InMux I__3187 (
            .O(N__20941),
            .I(N__20934));
    InMux I__3186 (
            .O(N__20940),
            .I(N__20931));
    LocalMux I__3185 (
            .O(N__20937),
            .I(N__20926));
    LocalMux I__3184 (
            .O(N__20934),
            .I(N__20926));
    LocalMux I__3183 (
            .O(N__20931),
            .I(ctrlOut_15));
    Odrv12 I__3182 (
            .O(N__20926),
            .I(ctrlOut_15));
    CascadeMux I__3181 (
            .O(N__20921),
            .I(\ALU.N_7_0_cascade_ ));
    InMux I__3180 (
            .O(N__20918),
            .I(N__20908));
    InMux I__3179 (
            .O(N__20917),
            .I(N__20908));
    InMux I__3178 (
            .O(N__20916),
            .I(N__20908));
    InMux I__3177 (
            .O(N__20915),
            .I(N__20905));
    LocalMux I__3176 (
            .O(N__20908),
            .I(N__20902));
    LocalMux I__3175 (
            .O(N__20905),
            .I(N__20899));
    Sp12to4 I__3174 (
            .O(N__20902),
            .I(N__20896));
    Span4Mux_v I__3173 (
            .O(N__20899),
            .I(N__20891));
    Span12Mux_s5_h I__3172 (
            .O(N__20896),
            .I(N__20888));
    InMux I__3171 (
            .O(N__20895),
            .I(N__20885));
    InMux I__3170 (
            .O(N__20894),
            .I(N__20882));
    Odrv4 I__3169 (
            .O(N__20891),
            .I(\ALU.N_179_0 ));
    Odrv12 I__3168 (
            .O(N__20888),
            .I(\ALU.N_179_0 ));
    LocalMux I__3167 (
            .O(N__20885),
            .I(\ALU.N_179_0 ));
    LocalMux I__3166 (
            .O(N__20882),
            .I(\ALU.N_179_0 ));
    CascadeMux I__3165 (
            .O(N__20873),
            .I(\ALU.a_15_m2_ns_1Z0Z_13_cascade_ ));
    InMux I__3164 (
            .O(N__20870),
            .I(N__20861));
    InMux I__3163 (
            .O(N__20869),
            .I(N__20861));
    InMux I__3162 (
            .O(N__20868),
            .I(N__20858));
    InMux I__3161 (
            .O(N__20867),
            .I(N__20855));
    InMux I__3160 (
            .O(N__20866),
            .I(N__20852));
    LocalMux I__3159 (
            .O(N__20861),
            .I(N__20849));
    LocalMux I__3158 (
            .O(N__20858),
            .I(N__20846));
    LocalMux I__3157 (
            .O(N__20855),
            .I(N__20843));
    LocalMux I__3156 (
            .O(N__20852),
            .I(N__20840));
    Span4Mux_v I__3155 (
            .O(N__20849),
            .I(N__20833));
    Span4Mux_s2_h I__3154 (
            .O(N__20846),
            .I(N__20833));
    Span4Mux_v I__3153 (
            .O(N__20843),
            .I(N__20833));
    Span4Mux_h I__3152 (
            .O(N__20840),
            .I(N__20830));
    Odrv4 I__3151 (
            .O(N__20833),
            .I(\ALU.operand2_9 ));
    Odrv4 I__3150 (
            .O(N__20830),
            .I(\ALU.operand2_9 ));
    InMux I__3149 (
            .O(N__20825),
            .I(N__20822));
    LocalMux I__3148 (
            .O(N__20822),
            .I(\ALU.N_220 ));
    CascadeMux I__3147 (
            .O(N__20819),
            .I(N__20816));
    InMux I__3146 (
            .O(N__20816),
            .I(N__20813));
    LocalMux I__3145 (
            .O(N__20813),
            .I(\ALU.N_250 ));
    CascadeMux I__3144 (
            .O(N__20810),
            .I(\ALU.N_250_cascade_ ));
    InMux I__3143 (
            .O(N__20807),
            .I(N__20804));
    LocalMux I__3142 (
            .O(N__20804),
            .I(\ALU.N_254 ));
    InMux I__3141 (
            .O(N__20801),
            .I(N__20798));
    LocalMux I__3140 (
            .O(N__20798),
            .I(\ALU.N_218 ));
    CascadeMux I__3139 (
            .O(N__20795),
            .I(\ALU.N_218_cascade_ ));
    CascadeMux I__3138 (
            .O(N__20792),
            .I(\ALU.N_361_cascade_ ));
    InMux I__3137 (
            .O(N__20789),
            .I(N__20785));
    InMux I__3136 (
            .O(N__20788),
            .I(N__20782));
    LocalMux I__3135 (
            .O(N__20785),
            .I(\ALU.N_252 ));
    LocalMux I__3134 (
            .O(N__20782),
            .I(\ALU.N_252 ));
    InMux I__3133 (
            .O(N__20777),
            .I(N__20774));
    LocalMux I__3132 (
            .O(N__20774),
            .I(\ALU.N_257 ));
    CascadeMux I__3131 (
            .O(N__20771),
            .I(\ALU.N_249_cascade_ ));
    InMux I__3130 (
            .O(N__20768),
            .I(N__20762));
    InMux I__3129 (
            .O(N__20767),
            .I(N__20762));
    LocalMux I__3128 (
            .O(N__20762),
            .I(\ALU.N_253 ));
    CascadeMux I__3127 (
            .O(N__20759),
            .I(\ALU.c_RNIUGCLVZ0Z_11_cascade_ ));
    InMux I__3126 (
            .O(N__20756),
            .I(N__20752));
    InMux I__3125 (
            .O(N__20755),
            .I(N__20749));
    LocalMux I__3124 (
            .O(N__20752),
            .I(\ALU.N_415 ));
    LocalMux I__3123 (
            .O(N__20749),
            .I(\ALU.N_415 ));
    InMux I__3122 (
            .O(N__20744),
            .I(N__20741));
    LocalMux I__3121 (
            .O(N__20741),
            .I(\ALU.N_310 ));
    CascadeMux I__3120 (
            .O(N__20738),
            .I(\ALU.lshift_3_ns_1_4_cascade_ ));
    InMux I__3119 (
            .O(N__20735),
            .I(N__20732));
    LocalMux I__3118 (
            .O(N__20732),
            .I(N__20729));
    Span4Mux_h I__3117 (
            .O(N__20729),
            .I(N__20726));
    Span4Mux_v I__3116 (
            .O(N__20726),
            .I(N__20723));
    Odrv4 I__3115 (
            .O(N__20723),
            .I(\ALU.N_273_0 ));
    InMux I__3114 (
            .O(N__20720),
            .I(N__20717));
    LocalMux I__3113 (
            .O(N__20717),
            .I(\ALU.N_461 ));
    InMux I__3112 (
            .O(N__20714),
            .I(N__20711));
    LocalMux I__3111 (
            .O(N__20711),
            .I(N__20708));
    Odrv4 I__3110 (
            .O(N__20708),
            .I(\ALU.N_474 ));
    CascadeMux I__3109 (
            .O(N__20705),
            .I(\ALU.N_530_cascade_ ));
    InMux I__3108 (
            .O(N__20702),
            .I(N__20696));
    InMux I__3107 (
            .O(N__20701),
            .I(N__20696));
    LocalMux I__3106 (
            .O(N__20696),
            .I(\ALU.N_635 ));
    CascadeMux I__3105 (
            .O(N__20693),
            .I(\ALU.d_RNIP8ITN1Z0Z_5_cascade_ ));
    InMux I__3104 (
            .O(N__20690),
            .I(N__20687));
    LocalMux I__3103 (
            .O(N__20687),
            .I(N__20684));
    Odrv4 I__3102 (
            .O(N__20684),
            .I(\ALU.d_RNILBFG4Z0Z_2 ));
    CascadeMux I__3101 (
            .O(N__20681),
            .I(\ALU.a_15_m3_2_cascade_ ));
    CascadeMux I__3100 (
            .O(N__20678),
            .I(\ALU.d_RNIE937BZ0Z_0_cascade_ ));
    InMux I__3099 (
            .O(N__20675),
            .I(N__20672));
    LocalMux I__3098 (
            .O(N__20672),
            .I(\ALU.a_15_m4_2 ));
    InMux I__3097 (
            .O(N__20669),
            .I(N__20663));
    InMux I__3096 (
            .O(N__20668),
            .I(N__20663));
    LocalMux I__3095 (
            .O(N__20663),
            .I(\FTDI.N_28 ));
    InMux I__3094 (
            .O(N__20660),
            .I(N__20657));
    LocalMux I__3093 (
            .O(N__20657),
            .I(\ALU.a_15_m1_0 ));
    CascadeMux I__3092 (
            .O(N__20654),
            .I(\ALU.a_15_m4_ns_1_0_cascade_ ));
    CascadeMux I__3091 (
            .O(N__20651),
            .I(\ALU.a_15_m4_0_cascade_ ));
    InMux I__3090 (
            .O(N__20648),
            .I(N__20645));
    LocalMux I__3089 (
            .O(N__20645),
            .I(\ALU.a_15_m3_0 ));
    InMux I__3088 (
            .O(N__20642),
            .I(N__20639));
    LocalMux I__3087 (
            .O(N__20639),
            .I(N__20636));
    Span4Mux_v I__3086 (
            .O(N__20636),
            .I(N__20633));
    Span4Mux_v I__3085 (
            .O(N__20633),
            .I(N__20630));
    Span4Mux_s1_v I__3084 (
            .O(N__20630),
            .I(N__20627));
    Odrv4 I__3083 (
            .O(N__20627),
            .I(\ALU.a_15_m4_bm_1Z0Z_8 ));
    InMux I__3082 (
            .O(N__20624),
            .I(N__20621));
    LocalMux I__3081 (
            .O(N__20621),
            .I(\ALU.a_15_m0_0 ));
    InMux I__3080 (
            .O(N__20618),
            .I(N__20615));
    LocalMux I__3079 (
            .O(N__20615),
            .I(N__20612));
    Span4Mux_h I__3078 (
            .O(N__20612),
            .I(N__20609));
    Odrv4 I__3077 (
            .O(N__20609),
            .I(i53_mux_0));
    InMux I__3076 (
            .O(N__20606),
            .I(N__20603));
    LocalMux I__3075 (
            .O(N__20603),
            .I(\ALU.madd_33 ));
    InMux I__3074 (
            .O(N__20600),
            .I(N__20597));
    LocalMux I__3073 (
            .O(N__20597),
            .I(\ALU.madd_68_0_tz ));
    InMux I__3072 (
            .O(N__20594),
            .I(N__20591));
    LocalMux I__3071 (
            .O(N__20591),
            .I(\ALU.madd_68 ));
    InMux I__3070 (
            .O(N__20588),
            .I(N__20582));
    InMux I__3069 (
            .O(N__20587),
            .I(N__20582));
    LocalMux I__3068 (
            .O(N__20582),
            .I(N__20579));
    Odrv4 I__3067 (
            .O(N__20579),
            .I(\ALU.madd_89_0 ));
    CascadeMux I__3066 (
            .O(N__20576),
            .I(\ALU.madd_68_cascade_ ));
    InMux I__3065 (
            .O(N__20573),
            .I(N__20567));
    InMux I__3064 (
            .O(N__20572),
            .I(N__20567));
    LocalMux I__3063 (
            .O(N__20567),
            .I(N__20563));
    InMux I__3062 (
            .O(N__20566),
            .I(N__20560));
    Odrv4 I__3061 (
            .O(N__20563),
            .I(\ALU.a7_b_1 ));
    LocalMux I__3060 (
            .O(N__20560),
            .I(\ALU.a7_b_1 ));
    InMux I__3059 (
            .O(N__20555),
            .I(N__20549));
    InMux I__3058 (
            .O(N__20554),
            .I(N__20549));
    LocalMux I__3057 (
            .O(N__20549),
            .I(\ALU.madd_108 ));
    CascadeMux I__3056 (
            .O(N__20546),
            .I(\ALU.madd_108_cascade_ ));
    InMux I__3055 (
            .O(N__20543),
            .I(N__20534));
    InMux I__3054 (
            .O(N__20542),
            .I(N__20534));
    InMux I__3053 (
            .O(N__20541),
            .I(N__20534));
    LocalMux I__3052 (
            .O(N__20534),
            .I(N__20531));
    Span4Mux_h I__3051 (
            .O(N__20531),
            .I(N__20528));
    Odrv4 I__3050 (
            .O(N__20528),
            .I(\ALU.madd_134 ));
    InMux I__3049 (
            .O(N__20525),
            .I(N__20519));
    InMux I__3048 (
            .O(N__20524),
            .I(N__20519));
    LocalMux I__3047 (
            .O(N__20519),
            .I(N__20516));
    Span4Mux_h I__3046 (
            .O(N__20516),
            .I(N__20513));
    Odrv4 I__3045 (
            .O(N__20513),
            .I(\ALU.madd_153 ));
    CEMux I__3044 (
            .O(N__20510),
            .I(N__20506));
    CEMux I__3043 (
            .O(N__20509),
            .I(N__20503));
    LocalMux I__3042 (
            .O(N__20506),
            .I(N__20500));
    LocalMux I__3041 (
            .O(N__20503),
            .I(N__20497));
    Span4Mux_s1_h I__3040 (
            .O(N__20500),
            .I(N__20494));
    Span12Mux_v I__3039 (
            .O(N__20497),
            .I(N__20491));
    Span4Mux_h I__3038 (
            .O(N__20494),
            .I(N__20488));
    Odrv12 I__3037 (
            .O(N__20491),
            .I(\FTDI.N_201_2 ));
    Odrv4 I__3036 (
            .O(N__20488),
            .I(\FTDI.N_201_2 ));
    InMux I__3035 (
            .O(N__20483),
            .I(N__20480));
    LocalMux I__3034 (
            .O(N__20480),
            .I(N__20475));
    InMux I__3033 (
            .O(N__20479),
            .I(N__20472));
    InMux I__3032 (
            .O(N__20478),
            .I(N__20469));
    Odrv4 I__3031 (
            .O(N__20475),
            .I(aluOperation_3));
    LocalMux I__3030 (
            .O(N__20472),
            .I(aluOperation_3));
    LocalMux I__3029 (
            .O(N__20469),
            .I(aluOperation_3));
    CascadeMux I__3028 (
            .O(N__20462),
            .I(\ALU.m681Z0Z_1_cascade_ ));
    InMux I__3027 (
            .O(N__20459),
            .I(N__20450));
    InMux I__3026 (
            .O(N__20458),
            .I(N__20445));
    InMux I__3025 (
            .O(N__20457),
            .I(N__20445));
    InMux I__3024 (
            .O(N__20456),
            .I(N__20436));
    InMux I__3023 (
            .O(N__20455),
            .I(N__20436));
    InMux I__3022 (
            .O(N__20454),
            .I(N__20436));
    InMux I__3021 (
            .O(N__20453),
            .I(N__20436));
    LocalMux I__3020 (
            .O(N__20450),
            .I(N__20428));
    LocalMux I__3019 (
            .O(N__20445),
            .I(N__20428));
    LocalMux I__3018 (
            .O(N__20436),
            .I(N__20428));
    InMux I__3017 (
            .O(N__20435),
            .I(N__20425));
    Span4Mux_v I__3016 (
            .O(N__20428),
            .I(N__20420));
    LocalMux I__3015 (
            .O(N__20425),
            .I(N__20420));
    Odrv4 I__3014 (
            .O(N__20420),
            .I(\ALU.N_730_mux ));
    CascadeMux I__3013 (
            .O(N__20417),
            .I(\ALU.a7_b_0_cascade_ ));
    InMux I__3012 (
            .O(N__20414),
            .I(N__20411));
    LocalMux I__3011 (
            .O(N__20411),
            .I(N__20408));
    Span4Mux_h I__3010 (
            .O(N__20408),
            .I(N__20404));
    InMux I__3009 (
            .O(N__20407),
            .I(N__20401));
    Odrv4 I__3008 (
            .O(N__20404),
            .I(\ALU.madd_59 ));
    LocalMux I__3007 (
            .O(N__20401),
            .I(\ALU.madd_59 ));
    CascadeMux I__3006 (
            .O(N__20396),
            .I(N__20393));
    InMux I__3005 (
            .O(N__20393),
            .I(N__20390));
    LocalMux I__3004 (
            .O(N__20390),
            .I(N__20387));
    Span4Mux_h I__3003 (
            .O(N__20387),
            .I(N__20384));
    Span4Mux_v I__3002 (
            .O(N__20384),
            .I(N__20381));
    Span4Mux_h I__3001 (
            .O(N__20381),
            .I(N__20378));
    Odrv4 I__3000 (
            .O(N__20378),
            .I(\ALU.madd_484_5 ));
    InMux I__2999 (
            .O(N__20375),
            .I(N__20372));
    LocalMux I__2998 (
            .O(N__20372),
            .I(N__20369));
    Odrv12 I__2997 (
            .O(N__20369),
            .I(\ALU.madd_128_0_tz_0 ));
    InMux I__2996 (
            .O(N__20366),
            .I(N__20360));
    InMux I__2995 (
            .O(N__20365),
            .I(N__20360));
    LocalMux I__2994 (
            .O(N__20360),
            .I(N__20357));
    Odrv12 I__2993 (
            .O(N__20357),
            .I(\ALU.madd_104 ));
    InMux I__2992 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__2991 (
            .O(N__20351),
            .I(N__20348));
    Span12Mux_s4_h I__2990 (
            .O(N__20348),
            .I(N__20344));
    InMux I__2989 (
            .O(N__20347),
            .I(N__20341));
    Odrv12 I__2988 (
            .O(N__20344),
            .I(\ALU.madd_149 ));
    LocalMux I__2987 (
            .O(N__20341),
            .I(\ALU.madd_149 ));
    InMux I__2986 (
            .O(N__20336),
            .I(N__20333));
    LocalMux I__2985 (
            .O(N__20333),
            .I(\ALU.madd_128_0_tz ));
    InMux I__2984 (
            .O(N__20330),
            .I(N__20324));
    InMux I__2983 (
            .O(N__20329),
            .I(N__20324));
    LocalMux I__2982 (
            .O(N__20324),
            .I(N__20321));
    Odrv4 I__2981 (
            .O(N__20321),
            .I(\ALU.madd_128_0 ));
    InMux I__2980 (
            .O(N__20318),
            .I(N__20315));
    LocalMux I__2979 (
            .O(N__20315),
            .I(N__20312));
    Span4Mux_h I__2978 (
            .O(N__20312),
            .I(N__20309));
    Odrv4 I__2977 (
            .O(N__20309),
            .I(\ALU.madd_N_1_i ));
    CascadeMux I__2976 (
            .O(N__20306),
            .I(\ALU.madd_20_0_cascade_ ));
    InMux I__2975 (
            .O(N__20303),
            .I(N__20294));
    InMux I__2974 (
            .O(N__20302),
            .I(N__20294));
    InMux I__2973 (
            .O(N__20301),
            .I(N__20294));
    LocalMux I__2972 (
            .O(N__20294),
            .I(\ALU.madd_20 ));
    InMux I__2971 (
            .O(N__20291),
            .I(N__20286));
    InMux I__2970 (
            .O(N__20290),
            .I(N__20281));
    InMux I__2969 (
            .O(N__20289),
            .I(N__20281));
    LocalMux I__2968 (
            .O(N__20286),
            .I(N__20278));
    LocalMux I__2967 (
            .O(N__20281),
            .I(N__20273));
    Span12Mux_s9_h I__2966 (
            .O(N__20278),
            .I(N__20270));
    InMux I__2965 (
            .O(N__20277),
            .I(N__20265));
    InMux I__2964 (
            .O(N__20276),
            .I(N__20265));
    Span4Mux_v I__2963 (
            .O(N__20273),
            .I(N__20262));
    Span12Mux_v I__2962 (
            .O(N__20270),
            .I(N__20259));
    LocalMux I__2961 (
            .O(N__20265),
            .I(ctrlOut_2));
    Odrv4 I__2960 (
            .O(N__20262),
            .I(ctrlOut_2));
    Odrv12 I__2959 (
            .O(N__20259),
            .I(ctrlOut_2));
    CascadeMux I__2958 (
            .O(N__20252),
            .I(\ALU.N_5_0_cascade_ ));
    CascadeMux I__2957 (
            .O(N__20249),
            .I(\ALU.N_240_0_cascade_ ));
    InMux I__2956 (
            .O(N__20246),
            .I(N__20243));
    LocalMux I__2955 (
            .O(N__20243),
            .I(\ALU.madd_24_0_tz ));
    InMux I__2954 (
            .O(N__20240),
            .I(N__20237));
    LocalMux I__2953 (
            .O(N__20237),
            .I(N__20234));
    Span4Mux_h I__2952 (
            .O(N__20234),
            .I(N__20231));
    Odrv4 I__2951 (
            .O(N__20231),
            .I(\ALU.madd_8_0 ));
    InMux I__2950 (
            .O(N__20228),
            .I(N__20225));
    LocalMux I__2949 (
            .O(N__20225),
            .I(N__20222));
    Span4Mux_h I__2948 (
            .O(N__20222),
            .I(N__20219));
    Odrv4 I__2947 (
            .O(N__20219),
            .I(\ALU.madd_5 ));
    CascadeMux I__2946 (
            .O(N__20216),
            .I(\ALU.madd_8_0_cascade_ ));
    CascadeMux I__2945 (
            .O(N__20213),
            .I(\ALU.N_706_cascade_ ));
    InMux I__2944 (
            .O(N__20210),
            .I(N__20207));
    LocalMux I__2943 (
            .O(N__20207),
            .I(\ALU.N_754 ));
    CascadeMux I__2942 (
            .O(N__20204),
            .I(\ALU.aluOut_7_cascade_ ));
    InMux I__2941 (
            .O(N__20201),
            .I(N__20198));
    LocalMux I__2940 (
            .O(N__20198),
            .I(N__20195));
    Span4Mux_h I__2939 (
            .O(N__20195),
            .I(N__20192));
    Span4Mux_v I__2938 (
            .O(N__20192),
            .I(N__20189));
    Odrv4 I__2937 (
            .O(N__20189),
            .I(\ALU.a7_b_0_6 ));
    CascadeMux I__2936 (
            .O(N__20186),
            .I(N__20183));
    InMux I__2935 (
            .O(N__20183),
            .I(N__20180));
    LocalMux I__2934 (
            .O(N__20180),
            .I(N__20177));
    Span4Mux_h I__2933 (
            .O(N__20177),
            .I(N__20174));
    Odrv4 I__2932 (
            .O(N__20174),
            .I(\ALU.m271_nsZ0Z_1 ));
    CascadeMux I__2931 (
            .O(N__20171),
            .I(\ALU.N_708_cascade_ ));
    CascadeMux I__2930 (
            .O(N__20168),
            .I(\ALU.dout_6_ns_1_9_cascade_ ));
    InMux I__2929 (
            .O(N__20165),
            .I(N__20162));
    LocalMux I__2928 (
            .O(N__20162),
            .I(\ALU.N_756 ));
    CascadeMux I__2927 (
            .O(N__20159),
            .I(\ALU.N_751_cascade_ ));
    InMux I__2926 (
            .O(N__20156),
            .I(N__20153));
    LocalMux I__2925 (
            .O(N__20153),
            .I(\ALU.N_703 ));
    CascadeMux I__2924 (
            .O(N__20150),
            .I(\ALU.rshift_3_ns_1_4_cascade_ ));
    InMux I__2923 (
            .O(N__20147),
            .I(N__20144));
    LocalMux I__2922 (
            .O(N__20144),
            .I(N__20141));
    Span12Mux_s11_v I__2921 (
            .O(N__20141),
            .I(N__20138));
    Odrv12 I__2920 (
            .O(N__20138),
            .I(\ALU.N_472 ));
    CascadeMux I__2919 (
            .O(N__20135),
            .I(\ALU.N_472_cascade_ ));
    InMux I__2918 (
            .O(N__20132),
            .I(N__20129));
    LocalMux I__2917 (
            .O(N__20129),
            .I(N__20126));
    Span4Mux_v I__2916 (
            .O(N__20126),
            .I(N__20123));
    Span4Mux_v I__2915 (
            .O(N__20123),
            .I(N__20119));
    InMux I__2914 (
            .O(N__20122),
            .I(N__20116));
    Odrv4 I__2913 (
            .O(N__20119),
            .I(\ALU.N_476 ));
    LocalMux I__2912 (
            .O(N__20116),
            .I(\ALU.N_476 ));
    CascadeMux I__2911 (
            .O(N__20111),
            .I(\ALU.m272_nsZ0Z_1_cascade_ ));
    CascadeMux I__2910 (
            .O(N__20108),
            .I(N__20105));
    InMux I__2909 (
            .O(N__20105),
            .I(N__20102));
    LocalMux I__2908 (
            .O(N__20102),
            .I(N__20099));
    Span4Mux_v I__2907 (
            .O(N__20099),
            .I(N__20096));
    Span4Mux_h I__2906 (
            .O(N__20096),
            .I(N__20093));
    Odrv4 I__2905 (
            .O(N__20093),
            .I(\ALU.N_191_0_0 ));
    CascadeMux I__2904 (
            .O(N__20090),
            .I(N__20084));
    InMux I__2903 (
            .O(N__20089),
            .I(N__20069));
    InMux I__2902 (
            .O(N__20088),
            .I(N__20069));
    InMux I__2901 (
            .O(N__20087),
            .I(N__20069));
    InMux I__2900 (
            .O(N__20084),
            .I(N__20069));
    InMux I__2899 (
            .O(N__20083),
            .I(N__20069));
    InMux I__2898 (
            .O(N__20082),
            .I(N__20069));
    LocalMux I__2897 (
            .O(N__20069),
            .I(ctrlOut_10));
    CascadeMux I__2896 (
            .O(N__20066),
            .I(N__20062));
    CascadeMux I__2895 (
            .O(N__20065),
            .I(N__20059));
    InMux I__2894 (
            .O(N__20062),
            .I(N__20054));
    InMux I__2893 (
            .O(N__20059),
            .I(N__20054));
    LocalMux I__2892 (
            .O(N__20054),
            .I(N__20051));
    Span4Mux_v I__2891 (
            .O(N__20051),
            .I(N__20048));
    IoSpan4Mux I__2890 (
            .O(N__20048),
            .I(N__20045));
    Span4Mux_s2_h I__2889 (
            .O(N__20045),
            .I(N__20042));
    Span4Mux_v I__2888 (
            .O(N__20042),
            .I(N__20037));
    InMux I__2887 (
            .O(N__20041),
            .I(N__20032));
    InMux I__2886 (
            .O(N__20040),
            .I(N__20032));
    Odrv4 I__2885 (
            .O(N__20037),
            .I(\ALU.N_191_0 ));
    LocalMux I__2884 (
            .O(N__20032),
            .I(\ALU.N_191_0 ));
    CascadeMux I__2883 (
            .O(N__20027),
            .I(\ALU.N_191_0_cascade_ ));
    InMux I__2882 (
            .O(N__20024),
            .I(N__20015));
    InMux I__2881 (
            .O(N__20023),
            .I(N__20015));
    InMux I__2880 (
            .O(N__20022),
            .I(N__20015));
    LocalMux I__2879 (
            .O(N__20015),
            .I(N__20010));
    InMux I__2878 (
            .O(N__20014),
            .I(N__20007));
    InMux I__2877 (
            .O(N__20013),
            .I(N__20004));
    Odrv4 I__2876 (
            .O(N__20010),
            .I(\ALU.operand2_10 ));
    LocalMux I__2875 (
            .O(N__20007),
            .I(\ALU.operand2_10 ));
    LocalMux I__2874 (
            .O(N__20004),
            .I(\ALU.operand2_10 ));
    InMux I__2873 (
            .O(N__19997),
            .I(N__19994));
    LocalMux I__2872 (
            .O(N__19994),
            .I(N__19991));
    Span4Mux_s3_h I__2871 (
            .O(N__19991),
            .I(N__19988));
    Odrv4 I__2870 (
            .O(N__19988),
            .I(\ALU.a1_b_10 ));
    CascadeMux I__2869 (
            .O(N__19985),
            .I(\ALU.a1_b_10_cascade_ ));
    InMux I__2868 (
            .O(N__19982),
            .I(N__19975));
    InMux I__2867 (
            .O(N__19981),
            .I(N__19975));
    InMux I__2866 (
            .O(N__19980),
            .I(N__19972));
    LocalMux I__2865 (
            .O(N__19975),
            .I(N__19969));
    LocalMux I__2864 (
            .O(N__19972),
            .I(N__19964));
    Span12Mux_v I__2863 (
            .O(N__19969),
            .I(N__19964));
    Odrv12 I__2862 (
            .O(N__19964),
            .I(\ALU.madd_203 ));
    InMux I__2861 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__2860 (
            .O(N__19958),
            .I(N__19955));
    Span4Mux_v I__2859 (
            .O(N__19955),
            .I(N__19951));
    InMux I__2858 (
            .O(N__19954),
            .I(N__19948));
    Odrv4 I__2857 (
            .O(N__19951),
            .I(\ALU.a9_b_2 ));
    LocalMux I__2856 (
            .O(N__19948),
            .I(\ALU.a9_b_2 ));
    CascadeMux I__2855 (
            .O(N__19943),
            .I(\ALU.dout_3_ns_1_9_cascade_ ));
    CascadeMux I__2854 (
            .O(N__19940),
            .I(\ALU.N_186_0_cascade_ ));
    InMux I__2853 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__2852 (
            .O(N__19934),
            .I(\ALU.a1_b_11 ));
    InMux I__2851 (
            .O(N__19931),
            .I(N__19925));
    InMux I__2850 (
            .O(N__19930),
            .I(N__19925));
    LocalMux I__2849 (
            .O(N__19925),
            .I(\ALU.a0_b_12 ));
    CascadeMux I__2848 (
            .O(N__19922),
            .I(\ALU.a1_b_11_cascade_ ));
    InMux I__2847 (
            .O(N__19919),
            .I(N__19916));
    LocalMux I__2846 (
            .O(N__19916),
            .I(N__19912));
    InMux I__2845 (
            .O(N__19915),
            .I(N__19909));
    Span4Mux_v I__2844 (
            .O(N__19912),
            .I(N__19904));
    LocalMux I__2843 (
            .O(N__19909),
            .I(N__19904));
    Span4Mux_h I__2842 (
            .O(N__19904),
            .I(N__19901));
    Odrv4 I__2841 (
            .O(N__19901),
            .I(\ALU.madd_255 ));
    CascadeMux I__2840 (
            .O(N__19898),
            .I(\ALU.dout_6_ns_1_8_cascade_ ));
    InMux I__2839 (
            .O(N__19895),
            .I(N__19892));
    LocalMux I__2838 (
            .O(N__19892),
            .I(\ALU.dout_3_ns_1_8 ));
    CascadeMux I__2837 (
            .O(N__19889),
            .I(\ALU.N_707_cascade_ ));
    InMux I__2836 (
            .O(N__19886),
            .I(N__19883));
    LocalMux I__2835 (
            .O(N__19883),
            .I(\ALU.N_755 ));
    InMux I__2834 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__2833 (
            .O(N__19877),
            .I(N__19874));
    Odrv12 I__2832 (
            .O(N__19874),
            .I(\ALU.N_283_0 ));
    InMux I__2831 (
            .O(N__19871),
            .I(N__19868));
    LocalMux I__2830 (
            .O(N__19868),
            .I(N__19864));
    InMux I__2829 (
            .O(N__19867),
            .I(N__19861));
    Span4Mux_v I__2828 (
            .O(N__19864),
            .I(N__19858));
    LocalMux I__2827 (
            .O(N__19861),
            .I(ctrlOut_7));
    Odrv4 I__2826 (
            .O(N__19858),
            .I(ctrlOut_7));
    InMux I__2825 (
            .O(N__19853),
            .I(N__19850));
    LocalMux I__2824 (
            .O(N__19850),
            .I(N__19846));
    InMux I__2823 (
            .O(N__19849),
            .I(N__19843));
    Span4Mux_v I__2822 (
            .O(N__19846),
            .I(N__19839));
    LocalMux I__2821 (
            .O(N__19843),
            .I(N__19834));
    InMux I__2820 (
            .O(N__19842),
            .I(N__19831));
    IoSpan4Mux I__2819 (
            .O(N__19839),
            .I(N__19828));
    InMux I__2818 (
            .O(N__19838),
            .I(N__19823));
    InMux I__2817 (
            .O(N__19837),
            .I(N__19823));
    Span4Mux_v I__2816 (
            .O(N__19834),
            .I(N__19816));
    LocalMux I__2815 (
            .O(N__19831),
            .I(N__19813));
    Span4Mux_s1_h I__2814 (
            .O(N__19828),
            .I(N__19808));
    LocalMux I__2813 (
            .O(N__19823),
            .I(N__19808));
    InMux I__2812 (
            .O(N__19822),
            .I(N__19805));
    InMux I__2811 (
            .O(N__19821),
            .I(N__19802));
    InMux I__2810 (
            .O(N__19820),
            .I(N__19799));
    InMux I__2809 (
            .O(N__19819),
            .I(N__19796));
    Span4Mux_s1_h I__2808 (
            .O(N__19816),
            .I(N__19789));
    Span4Mux_h I__2807 (
            .O(N__19813),
            .I(N__19789));
    Span4Mux_v I__2806 (
            .O(N__19808),
            .I(N__19789));
    LocalMux I__2805 (
            .O(N__19805),
            .I(N__19785));
    LocalMux I__2804 (
            .O(N__19802),
            .I(N__19778));
    LocalMux I__2803 (
            .O(N__19799),
            .I(N__19778));
    LocalMux I__2802 (
            .O(N__19796),
            .I(N__19778));
    Span4Mux_v I__2801 (
            .O(N__19789),
            .I(N__19775));
    InMux I__2800 (
            .O(N__19788),
            .I(N__19772));
    Span12Mux_s6_v I__2799 (
            .O(N__19785),
            .I(N__19767));
    Span12Mux_v I__2798 (
            .O(N__19778),
            .I(N__19767));
    Span4Mux_s1_h I__2797 (
            .O(N__19775),
            .I(N__19764));
    LocalMux I__2796 (
            .O(N__19772),
            .I(\ALU.N_211_0 ));
    Odrv12 I__2795 (
            .O(N__19767),
            .I(\ALU.N_211_0 ));
    Odrv4 I__2794 (
            .O(N__19764),
            .I(\ALU.N_211_0 ));
    CascadeMux I__2793 (
            .O(N__19757),
            .I(N__19754));
    InMux I__2792 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__2791 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_h I__2790 (
            .O(N__19748),
            .I(N__19744));
    InMux I__2789 (
            .O(N__19747),
            .I(N__19741));
    Span4Mux_h I__2788 (
            .O(N__19744),
            .I(N__19738));
    LocalMux I__2787 (
            .O(N__19741),
            .I(ctrlOut_9));
    Odrv4 I__2786 (
            .O(N__19738),
            .I(ctrlOut_9));
    InMux I__2785 (
            .O(N__19733),
            .I(N__19727));
    InMux I__2784 (
            .O(N__19732),
            .I(N__19727));
    LocalMux I__2783 (
            .O(N__19727),
            .I(N__19724));
    Span4Mux_v I__2782 (
            .O(N__19724),
            .I(N__19721));
    Odrv4 I__2781 (
            .O(N__19721),
            .I(\ALU.madd_367 ));
    CascadeMux I__2780 (
            .O(N__19718),
            .I(N__19715));
    InMux I__2779 (
            .O(N__19715),
            .I(N__19712));
    LocalMux I__2778 (
            .O(N__19712),
            .I(\ALU.d_RNIRV558Z0Z_13 ));
    CascadeMux I__2777 (
            .O(N__19709),
            .I(\ALU.d_RNIRV558Z0Z_13_cascade_ ));
    InMux I__2776 (
            .O(N__19706),
            .I(N__19703));
    LocalMux I__2775 (
            .O(N__19703),
            .I(N__19700));
    Odrv4 I__2774 (
            .O(N__19700),
            .I(\ALU.madd_371 ));
    InMux I__2773 (
            .O(N__19697),
            .I(N__19691));
    InMux I__2772 (
            .O(N__19696),
            .I(N__19691));
    LocalMux I__2771 (
            .O(N__19691),
            .I(\ALU.a2_b_12 ));
    InMux I__2770 (
            .O(N__19688),
            .I(N__19685));
    LocalMux I__2769 (
            .O(N__19685),
            .I(N__19681));
    InMux I__2768 (
            .O(N__19684),
            .I(N__19678));
    Span4Mux_h I__2767 (
            .O(N__19681),
            .I(N__19672));
    LocalMux I__2766 (
            .O(N__19678),
            .I(N__19672));
    InMux I__2765 (
            .O(N__19677),
            .I(N__19669));
    Odrv4 I__2764 (
            .O(N__19672),
            .I(\ALU.madd_259 ));
    LocalMux I__2763 (
            .O(N__19669),
            .I(\ALU.madd_259 ));
    CascadeMux I__2762 (
            .O(N__19664),
            .I(\ALU.N_240_0_i_cascade_ ));
    InMux I__2761 (
            .O(N__19661),
            .I(N__19655));
    InMux I__2760 (
            .O(N__19660),
            .I(N__19655));
    LocalMux I__2759 (
            .O(N__19655),
            .I(N__19652));
    Span4Mux_h I__2758 (
            .O(N__19652),
            .I(N__19648));
    InMux I__2757 (
            .O(N__19651),
            .I(N__19645));
    Odrv4 I__2756 (
            .O(N__19648),
            .I(\ALU.N_9_0 ));
    LocalMux I__2755 (
            .O(N__19645),
            .I(\ALU.N_9_0 ));
    InMux I__2754 (
            .O(N__19640),
            .I(N__19634));
    InMux I__2753 (
            .O(N__19639),
            .I(N__19634));
    LocalMux I__2752 (
            .O(N__19634),
            .I(N__19631));
    Span4Mux_v I__2751 (
            .O(N__19631),
            .I(N__19627));
    InMux I__2750 (
            .O(N__19630),
            .I(N__19624));
    Span4Mux_h I__2749 (
            .O(N__19627),
            .I(N__19621));
    LocalMux I__2748 (
            .O(N__19624),
            .I(N__19618));
    Odrv4 I__2747 (
            .O(N__19621),
            .I(\ALU.N_10_0 ));
    Odrv4 I__2746 (
            .O(N__19618),
            .I(\ALU.N_10_0 ));
    InMux I__2745 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__2744 (
            .O(N__19610),
            .I(N__19607));
    Span4Mux_h I__2743 (
            .O(N__19607),
            .I(N__19604));
    Odrv4 I__2742 (
            .O(N__19604),
            .I(\ALU.N_253_0 ));
    InMux I__2741 (
            .O(N__19601),
            .I(N__19598));
    LocalMux I__2740 (
            .O(N__19598),
            .I(N__19595));
    Span4Mux_s2_v I__2739 (
            .O(N__19595),
            .I(N__19592));
    Odrv4 I__2738 (
            .O(N__19592),
            .I(\ALU.d_RNIUV3H4Z0Z_0 ));
    CascadeMux I__2737 (
            .O(N__19589),
            .I(N__19585));
    InMux I__2736 (
            .O(N__19588),
            .I(N__19580));
    InMux I__2735 (
            .O(N__19585),
            .I(N__19580));
    LocalMux I__2734 (
            .O(N__19580),
            .I(N__19577));
    Span4Mux_h I__2733 (
            .O(N__19577),
            .I(N__19572));
    InMux I__2732 (
            .O(N__19576),
            .I(N__19567));
    InMux I__2731 (
            .O(N__19575),
            .I(N__19567));
    Odrv4 I__2730 (
            .O(N__19572),
            .I(\ALU.N_635_0 ));
    LocalMux I__2729 (
            .O(N__19567),
            .I(\ALU.N_635_0 ));
    CascadeMux I__2728 (
            .O(N__19562),
            .I(N__19559));
    InMux I__2727 (
            .O(N__19559),
            .I(N__19550));
    InMux I__2726 (
            .O(N__19558),
            .I(N__19550));
    InMux I__2725 (
            .O(N__19557),
            .I(N__19550));
    LocalMux I__2724 (
            .O(N__19550),
            .I(N__19547));
    Span4Mux_v I__2723 (
            .O(N__19547),
            .I(N__19544));
    Span4Mux_h I__2722 (
            .O(N__19544),
            .I(N__19541));
    Span4Mux_v I__2721 (
            .O(N__19541),
            .I(N__19536));
    CascadeMux I__2720 (
            .O(N__19540),
            .I(N__19533));
    CascadeMux I__2719 (
            .O(N__19539),
            .I(N__19530));
    Sp12to4 I__2718 (
            .O(N__19536),
            .I(N__19527));
    InMux I__2717 (
            .O(N__19533),
            .I(N__19522));
    InMux I__2716 (
            .O(N__19530),
            .I(N__19522));
    Span12Mux_s3_v I__2715 (
            .O(N__19527),
            .I(N__19519));
    LocalMux I__2714 (
            .O(N__19522),
            .I(\ALU.N_724 ));
    Odrv12 I__2713 (
            .O(N__19519),
            .I(\ALU.N_724 ));
    CascadeMux I__2712 (
            .O(N__19514),
            .I(\ALU.N_220_cascade_ ));
    InMux I__2711 (
            .O(N__19511),
            .I(N__19507));
    InMux I__2710 (
            .O(N__19510),
            .I(N__19504));
    LocalMux I__2709 (
            .O(N__19507),
            .I(\ALU.N_222 ));
    LocalMux I__2708 (
            .O(N__19504),
            .I(\ALU.N_222 ));
    InMux I__2707 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__2706 (
            .O(N__19496),
            .I(N__19493));
    Span4Mux_v I__2705 (
            .O(N__19493),
            .I(N__19490));
    Odrv4 I__2704 (
            .O(N__19490),
            .I(\ALU.madd_484_4 ));
    InMux I__2703 (
            .O(N__19487),
            .I(N__19484));
    LocalMux I__2702 (
            .O(N__19484),
            .I(\ALU.N_241_0 ));
    InMux I__2701 (
            .O(N__19481),
            .I(N__19478));
    LocalMux I__2700 (
            .O(N__19478),
            .I(\ALU.lshift_3_ns_1_15 ));
    CascadeMux I__2699 (
            .O(N__19475),
            .I(N__19472));
    InMux I__2698 (
            .O(N__19472),
            .I(N__19469));
    LocalMux I__2697 (
            .O(N__19469),
            .I(\ALU.dout_3_ns_1_14 ));
    CascadeMux I__2696 (
            .O(N__19466),
            .I(\ALU.lshift_3_ns_1_14_cascade_ ));
    InMux I__2695 (
            .O(N__19463),
            .I(N__19460));
    LocalMux I__2694 (
            .O(N__19460),
            .I(\ALU.N_256 ));
    CascadeMux I__2693 (
            .O(N__19457),
            .I(\ALU.N_224_cascade_ ));
    CascadeMux I__2692 (
            .O(N__19454),
            .I(\ALU.d_RNI8DL9U1Z0Z_3_cascade_ ));
    CascadeMux I__2691 (
            .O(N__19451),
            .I(\ALU.N_221_cascade_ ));
    CascadeMux I__2690 (
            .O(N__19448),
            .I(\ALU.N_588_cascade_ ));
    InMux I__2689 (
            .O(N__19445),
            .I(N__19442));
    LocalMux I__2688 (
            .O(N__19442),
            .I(\ALU.N_575 ));
    CascadeMux I__2687 (
            .O(N__19439),
            .I(\ALU.N_575_cascade_ ));
    InMux I__2686 (
            .O(N__19436),
            .I(N__19433));
    LocalMux I__2685 (
            .O(N__19433),
            .I(\ALU.rshift_3_ns_1_8 ));
    InMux I__2684 (
            .O(N__19430),
            .I(N__19427));
    LocalMux I__2683 (
            .O(N__19427),
            .I(N__19424));
    Span4Mux_s1_v I__2682 (
            .O(N__19424),
            .I(N__19421));
    Odrv4 I__2681 (
            .O(N__19421),
            .I(\ALU.m55_bmZ0 ));
    InMux I__2680 (
            .O(N__19418),
            .I(N__19415));
    LocalMux I__2679 (
            .O(N__19415),
            .I(N__19412));
    Odrv12 I__2678 (
            .O(N__19412),
            .I(\ALU.m55_amZ0 ));
    CascadeMux I__2677 (
            .O(N__19409),
            .I(\ALU.m650_nsZ0Z_1_cascade_ ));
    InMux I__2676 (
            .O(N__19406),
            .I(N__19400));
    InMux I__2675 (
            .O(N__19405),
            .I(N__19400));
    LocalMux I__2674 (
            .O(N__19400),
            .I(\ALU.N_15_0 ));
    InMux I__2673 (
            .O(N__19397),
            .I(N__19394));
    LocalMux I__2672 (
            .O(N__19394),
            .I(N_727));
    CascadeMux I__2671 (
            .O(N__19391),
            .I(\ALU.N_577_cascade_ ));
    CascadeMux I__2670 (
            .O(N__19388),
            .I(\ALU.N_528_cascade_ ));
    InMux I__2669 (
            .O(N__19385),
            .I(N__19382));
    LocalMux I__2668 (
            .O(N__19382),
            .I(N__19379));
    Span4Mux_v I__2667 (
            .O(N__19379),
            .I(N__19375));
    InMux I__2666 (
            .O(N__19378),
            .I(N__19372));
    Odrv4 I__2665 (
            .O(N__19375),
            .I(\ALU.N_633 ));
    LocalMux I__2664 (
            .O(N__19372),
            .I(\ALU.N_633 ));
    InMux I__2663 (
            .O(N__19367),
            .I(N__19364));
    LocalMux I__2662 (
            .O(N__19364),
            .I(N__19361));
    Span4Mux_h I__2661 (
            .O(N__19361),
            .I(N__19358));
    Odrv4 I__2660 (
            .O(N__19358),
            .I(\ALU.madd_144 ));
    InMux I__2659 (
            .O(N__19355),
            .I(N__19352));
    LocalMux I__2658 (
            .O(N__19352),
            .I(N__19349));
    Span4Mux_s3_h I__2657 (
            .O(N__19349),
            .I(N__19345));
    InMux I__2656 (
            .O(N__19348),
            .I(N__19342));
    Odrv4 I__2655 (
            .O(N__19345),
            .I(\ALU.madd_113 ));
    LocalMux I__2654 (
            .O(N__19342),
            .I(\ALU.madd_113 ));
    CascadeMux I__2653 (
            .O(N__19337),
            .I(\ALU.madd_154_cascade_ ));
    InMux I__2652 (
            .O(N__19334),
            .I(N__19330));
    InMux I__2651 (
            .O(N__19333),
            .I(N__19327));
    LocalMux I__2650 (
            .O(N__19330),
            .I(N__19322));
    LocalMux I__2649 (
            .O(N__19327),
            .I(N__19322));
    Span4Mux_h I__2648 (
            .O(N__19322),
            .I(N__19319));
    Span4Mux_v I__2647 (
            .O(N__19319),
            .I(N__19316));
    Odrv4 I__2646 (
            .O(N__19316),
            .I(\ALU.madd_99 ));
    InMux I__2645 (
            .O(N__19313),
            .I(N__19310));
    LocalMux I__2644 (
            .O(N__19310),
            .I(\ALU.madd_73 ));
    InMux I__2643 (
            .O(N__19307),
            .I(N__19303));
    InMux I__2642 (
            .O(N__19306),
            .I(N__19300));
    LocalMux I__2641 (
            .O(N__19303),
            .I(\ALU.madd_109 ));
    LocalMux I__2640 (
            .O(N__19300),
            .I(\ALU.madd_109 ));
    InMux I__2639 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__2638 (
            .O(N__19292),
            .I(N__19289));
    Span4Mux_v I__2637 (
            .O(N__19289),
            .I(N__19285));
    InMux I__2636 (
            .O(N__19288),
            .I(N__19282));
    Odrv4 I__2635 (
            .O(N__19285),
            .I(\ALU.madd_154 ));
    LocalMux I__2634 (
            .O(N__19282),
            .I(\ALU.madd_154 ));
    InMux I__2633 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__2632 (
            .O(N__19274),
            .I(N__19271));
    Span4Mux_v I__2631 (
            .O(N__19271),
            .I(N__19266));
    InMux I__2630 (
            .O(N__19270),
            .I(N__19261));
    InMux I__2629 (
            .O(N__19269),
            .I(N__19261));
    Odrv4 I__2628 (
            .O(N__19266),
            .I(\ALU.madd_118 ));
    LocalMux I__2627 (
            .O(N__19261),
            .I(\ALU.madd_118 ));
    CascadeMux I__2626 (
            .O(N__19256),
            .I(N__19253));
    InMux I__2625 (
            .O(N__19253),
            .I(N__19250));
    LocalMux I__2624 (
            .O(N__19250),
            .I(N__19247));
    Odrv4 I__2623 (
            .O(N__19247),
            .I(\ALU.m641_nsZ0Z_1 ));
    InMux I__2622 (
            .O(N__19244),
            .I(N__19241));
    LocalMux I__2621 (
            .O(N__19241),
            .I(N__19238));
    Span4Mux_s0_v I__2620 (
            .O(N__19238),
            .I(N__19235));
    Odrv4 I__2619 (
            .O(N__19235),
            .I(\ALU.m645_nsZ0Z_1 ));
    CascadeMux I__2618 (
            .O(N__19232),
            .I(\ALU.N_283_0_cascade_ ));
    CascadeMux I__2617 (
            .O(N__19229),
            .I(\ALU.madd_74_0_cascade_ ));
    InMux I__2616 (
            .O(N__19226),
            .I(N__19220));
    InMux I__2615 (
            .O(N__19225),
            .I(N__19220));
    LocalMux I__2614 (
            .O(N__19220),
            .I(\ALU.madd_83 ));
    CascadeMux I__2613 (
            .O(N__19217),
            .I(N__19212));
    InMux I__2612 (
            .O(N__19216),
            .I(N__19207));
    InMux I__2611 (
            .O(N__19215),
            .I(N__19207));
    InMux I__2610 (
            .O(N__19212),
            .I(N__19204));
    LocalMux I__2609 (
            .O(N__19207),
            .I(\ALU.madd_46 ));
    LocalMux I__2608 (
            .O(N__19204),
            .I(\ALU.madd_46 ));
    InMux I__2607 (
            .O(N__19199),
            .I(N__19193));
    InMux I__2606 (
            .O(N__19198),
            .I(N__19193));
    LocalMux I__2605 (
            .O(N__19193),
            .I(\ALU.madd_69 ));
    InMux I__2604 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__2603 (
            .O(N__19187),
            .I(\ALU.madd_74_0 ));
    InMux I__2602 (
            .O(N__19184),
            .I(N__19180));
    InMux I__2601 (
            .O(N__19183),
            .I(N__19177));
    LocalMux I__2600 (
            .O(N__19180),
            .I(\ALU.madd_79_0 ));
    LocalMux I__2599 (
            .O(N__19177),
            .I(\ALU.madd_79_0 ));
    InMux I__2598 (
            .O(N__19172),
            .I(N__19164));
    InMux I__2597 (
            .O(N__19171),
            .I(N__19164));
    InMux I__2596 (
            .O(N__19170),
            .I(N__19159));
    InMux I__2595 (
            .O(N__19169),
            .I(N__19159));
    LocalMux I__2594 (
            .O(N__19164),
            .I(N__19156));
    LocalMux I__2593 (
            .O(N__19159),
            .I(\ALU.madd_51 ));
    Odrv4 I__2592 (
            .O(N__19156),
            .I(\ALU.madd_51 ));
    InMux I__2591 (
            .O(N__19151),
            .I(N__19144));
    InMux I__2590 (
            .O(N__19150),
            .I(N__19144));
    InMux I__2589 (
            .O(N__19149),
            .I(N__19141));
    LocalMux I__2588 (
            .O(N__19144),
            .I(N__19136));
    LocalMux I__2587 (
            .O(N__19141),
            .I(N__19136));
    Odrv4 I__2586 (
            .O(N__19136),
            .I(\ALU.madd_58 ));
    CascadeMux I__2585 (
            .O(N__19133),
            .I(\ALU.madd_79_0_cascade_ ));
    InMux I__2584 (
            .O(N__19130),
            .I(N__19127));
    LocalMux I__2583 (
            .O(N__19127),
            .I(\ALU.madd_56 ));
    CascadeMux I__2582 (
            .O(N__19124),
            .I(\ALU.madd_88_cascade_ ));
    InMux I__2581 (
            .O(N__19121),
            .I(N__19118));
    LocalMux I__2580 (
            .O(N__19118),
            .I(\ALU.madd_114 ));
    InMux I__2579 (
            .O(N__19115),
            .I(N__19112));
    LocalMux I__2578 (
            .O(N__19112),
            .I(\ALU.madd_41 ));
    CascadeMux I__2577 (
            .O(N__19109),
            .I(\ALU.madd_73_cascade_ ));
    CascadeMux I__2576 (
            .O(N__19106),
            .I(N__19103));
    InMux I__2575 (
            .O(N__19103),
            .I(N__19099));
    InMux I__2574 (
            .O(N__19102),
            .I(N__19095));
    LocalMux I__2573 (
            .O(N__19099),
            .I(N__19092));
    InMux I__2572 (
            .O(N__19098),
            .I(N__19086));
    LocalMux I__2571 (
            .O(N__19095),
            .I(N__19082));
    Span4Mux_v I__2570 (
            .O(N__19092),
            .I(N__19077));
    InMux I__2569 (
            .O(N__19091),
            .I(N__19074));
    InMux I__2568 (
            .O(N__19090),
            .I(N__19069));
    InMux I__2567 (
            .O(N__19089),
            .I(N__19069));
    LocalMux I__2566 (
            .O(N__19086),
            .I(N__19066));
    InMux I__2565 (
            .O(N__19085),
            .I(N__19063));
    Span4Mux_v I__2564 (
            .O(N__19082),
            .I(N__19060));
    InMux I__2563 (
            .O(N__19081),
            .I(N__19055));
    InMux I__2562 (
            .O(N__19080),
            .I(N__19055));
    Odrv4 I__2561 (
            .O(N__19077),
            .I(\ALU.operand2_7 ));
    LocalMux I__2560 (
            .O(N__19074),
            .I(\ALU.operand2_7 ));
    LocalMux I__2559 (
            .O(N__19069),
            .I(\ALU.operand2_7 ));
    Odrv4 I__2558 (
            .O(N__19066),
            .I(\ALU.operand2_7 ));
    LocalMux I__2557 (
            .O(N__19063),
            .I(\ALU.operand2_7 ));
    Odrv4 I__2556 (
            .O(N__19060),
            .I(\ALU.operand2_7 ));
    LocalMux I__2555 (
            .O(N__19055),
            .I(\ALU.operand2_7 ));
    CascadeMux I__2554 (
            .O(N__19040),
            .I(N__19037));
    InMux I__2553 (
            .O(N__19037),
            .I(N__19033));
    InMux I__2552 (
            .O(N__19036),
            .I(N__19030));
    LocalMux I__2551 (
            .O(N__19033),
            .I(\ALU.a0_b_7 ));
    LocalMux I__2550 (
            .O(N__19030),
            .I(\ALU.a0_b_7 ));
    CascadeMux I__2549 (
            .O(N__19025),
            .I(\ALU.madd_12_cascade_ ));
    InMux I__2548 (
            .O(N__19022),
            .I(N__19019));
    LocalMux I__2547 (
            .O(N__19019),
            .I(\ALU.madd_34 ));
    InMux I__2546 (
            .O(N__19016),
            .I(N__19013));
    LocalMux I__2545 (
            .O(N__19013),
            .I(N__19010));
    Odrv4 I__2544 (
            .O(N__19010),
            .I(\ALU.madd_42 ));
    CascadeMux I__2543 (
            .O(N__19007),
            .I(\ALU.madd_34_cascade_ ));
    InMux I__2542 (
            .O(N__19004),
            .I(N__18997));
    InMux I__2541 (
            .O(N__19003),
            .I(N__18997));
    InMux I__2540 (
            .O(N__19002),
            .I(N__18994));
    LocalMux I__2539 (
            .O(N__18997),
            .I(\ALU.madd_37 ));
    LocalMux I__2538 (
            .O(N__18994),
            .I(\ALU.madd_37 ));
    CascadeMux I__2537 (
            .O(N__18989),
            .I(\ALU.madd_56_cascade_ ));
    InMux I__2536 (
            .O(N__18986),
            .I(N__18983));
    LocalMux I__2535 (
            .O(N__18983),
            .I(N__18980));
    Odrv4 I__2534 (
            .O(N__18980),
            .I(\ALU.madd_52_0 ));
    CascadeMux I__2533 (
            .O(N__18977),
            .I(N__18973));
    InMux I__2532 (
            .O(N__18976),
            .I(N__18965));
    InMux I__2531 (
            .O(N__18973),
            .I(N__18965));
    InMux I__2530 (
            .O(N__18972),
            .I(N__18965));
    LocalMux I__2529 (
            .O(N__18965),
            .I(N__18962));
    Span4Mux_v I__2528 (
            .O(N__18962),
            .I(N__18959));
    Odrv4 I__2527 (
            .O(N__18959),
            .I(\ALU.madd_25 ));
    CascadeMux I__2526 (
            .O(N__18956),
            .I(N__18953));
    InMux I__2525 (
            .O(N__18953),
            .I(N__18947));
    InMux I__2524 (
            .O(N__18952),
            .I(N__18947));
    LocalMux I__2523 (
            .O(N__18947),
            .I(\ALU.madd_12 ));
    CascadeMux I__2522 (
            .O(N__18944),
            .I(\ALU.un2_addsub_axb_6_cascade_ ));
    CascadeMux I__2521 (
            .O(N__18941),
            .I(N__18936));
    InMux I__2520 (
            .O(N__18940),
            .I(N__18931));
    InMux I__2519 (
            .O(N__18939),
            .I(N__18931));
    InMux I__2518 (
            .O(N__18936),
            .I(N__18928));
    LocalMux I__2517 (
            .O(N__18931),
            .I(N__18925));
    LocalMux I__2516 (
            .O(N__18928),
            .I(N__18922));
    Span4Mux_v I__2515 (
            .O(N__18925),
            .I(N__18919));
    Span4Mux_h I__2514 (
            .O(N__18922),
            .I(N__18916));
    Odrv4 I__2513 (
            .O(N__18919),
            .I(\ALU.madd_64_0 ));
    Odrv4 I__2512 (
            .O(N__18916),
            .I(\ALU.madd_64_0 ));
    CascadeMux I__2511 (
            .O(N__18911),
            .I(\ALU.a8_b_0_cascade_ ));
    CascadeMux I__2510 (
            .O(N__18908),
            .I(\ALU.madd_10_cascade_ ));
    InMux I__2509 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__2508 (
            .O(N__18902),
            .I(N__18899));
    Odrv4 I__2507 (
            .O(N__18899),
            .I(\ALU.madd_24 ));
    InMux I__2506 (
            .O(N__18896),
            .I(N__18893));
    LocalMux I__2505 (
            .O(N__18893),
            .I(N__18890));
    Span4Mux_v I__2504 (
            .O(N__18890),
            .I(N__18887));
    Odrv4 I__2503 (
            .O(N__18887),
            .I(\ALU.madd_29 ));
    CascadeMux I__2502 (
            .O(N__18884),
            .I(\ALU.madd_24_cascade_ ));
    CascadeMux I__2501 (
            .O(N__18881),
            .I(N__18878));
    InMux I__2500 (
            .O(N__18878),
            .I(N__18875));
    LocalMux I__2499 (
            .O(N__18875),
            .I(\ALU.madd_i1_mux_1 ));
    InMux I__2498 (
            .O(N__18872),
            .I(N__18869));
    LocalMux I__2497 (
            .O(N__18869),
            .I(N__18866));
    Odrv4 I__2496 (
            .O(N__18866),
            .I(\ALU.madd_i3_mux_0 ));
    InMux I__2495 (
            .O(N__18863),
            .I(N__18859));
    InMux I__2494 (
            .O(N__18862),
            .I(N__18856));
    LocalMux I__2493 (
            .O(N__18859),
            .I(N__18853));
    LocalMux I__2492 (
            .O(N__18856),
            .I(\ALU.a4_b_2 ));
    Odrv4 I__2491 (
            .O(N__18853),
            .I(\ALU.a4_b_2 ));
    CascadeMux I__2490 (
            .O(N__18848),
            .I(N__18845));
    InMux I__2489 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__2488 (
            .O(N__18842),
            .I(\ALU.a6_b_0 ));
    CascadeMux I__2487 (
            .O(N__18839),
            .I(\ALU.operand2_10_cascade_ ));
    InMux I__2486 (
            .O(N__18836),
            .I(N__18830));
    InMux I__2485 (
            .O(N__18835),
            .I(N__18830));
    LocalMux I__2484 (
            .O(N__18830),
            .I(N__18827));
    Span4Mux_s3_h I__2483 (
            .O(N__18827),
            .I(N__18824));
    Span4Mux_v I__2482 (
            .O(N__18824),
            .I(N__18821));
    Odrv4 I__2481 (
            .O(N__18821),
            .I(\ALU.a4_b_10 ));
    InMux I__2480 (
            .O(N__18818),
            .I(N__18815));
    LocalMux I__2479 (
            .O(N__18815),
            .I(\ALU.a3_b_10 ));
    CascadeMux I__2478 (
            .O(N__18812),
            .I(\ALU.a3_b_10_cascade_ ));
    InMux I__2477 (
            .O(N__18809),
            .I(N__18806));
    LocalMux I__2476 (
            .O(N__18806),
            .I(N__18802));
    InMux I__2475 (
            .O(N__18805),
            .I(N__18799));
    Odrv4 I__2474 (
            .O(N__18802),
            .I(\ALU.madd_305 ));
    LocalMux I__2473 (
            .O(N__18799),
            .I(\ALU.madd_305 ));
    CascadeMux I__2472 (
            .O(N__18794),
            .I(\ALU.madd_5_cascade_ ));
    InMux I__2471 (
            .O(N__18791),
            .I(N__18785));
    InMux I__2470 (
            .O(N__18790),
            .I(N__18785));
    LocalMux I__2469 (
            .O(N__18785),
            .I(\ALU.madd_19 ));
    InMux I__2468 (
            .O(N__18782),
            .I(N__18775));
    InMux I__2467 (
            .O(N__18781),
            .I(N__18775));
    InMux I__2466 (
            .O(N__18780),
            .I(N__18772));
    LocalMux I__2465 (
            .O(N__18775),
            .I(\ALU.madd_17 ));
    LocalMux I__2464 (
            .O(N__18772),
            .I(\ALU.madd_17 ));
    CascadeMux I__2463 (
            .O(N__18767),
            .I(\ALU.madd_19_cascade_ ));
    InMux I__2462 (
            .O(N__18764),
            .I(N__18761));
    LocalMux I__2461 (
            .O(N__18761),
            .I(\ALU.madd_47 ));
    CascadeMux I__2460 (
            .O(N__18758),
            .I(N__18755));
    InMux I__2459 (
            .O(N__18755),
            .I(N__18752));
    LocalMux I__2458 (
            .O(N__18752),
            .I(N__18749));
    Span4Mux_v I__2457 (
            .O(N__18749),
            .I(N__18746));
    Span4Mux_s1_h I__2456 (
            .O(N__18746),
            .I(N__18743));
    Odrv4 I__2455 (
            .O(N__18743),
            .I(\ALU.g0_0_a3_0 ));
    InMux I__2454 (
            .O(N__18740),
            .I(N__18735));
    InMux I__2453 (
            .O(N__18739),
            .I(N__18732));
    InMux I__2452 (
            .O(N__18738),
            .I(N__18724));
    LocalMux I__2451 (
            .O(N__18735),
            .I(N__18721));
    LocalMux I__2450 (
            .O(N__18732),
            .I(N__18718));
    InMux I__2449 (
            .O(N__18731),
            .I(N__18713));
    InMux I__2448 (
            .O(N__18730),
            .I(N__18710));
    InMux I__2447 (
            .O(N__18729),
            .I(N__18703));
    InMux I__2446 (
            .O(N__18728),
            .I(N__18703));
    InMux I__2445 (
            .O(N__18727),
            .I(N__18703));
    LocalMux I__2444 (
            .O(N__18724),
            .I(N__18698));
    Span4Mux_v I__2443 (
            .O(N__18721),
            .I(N__18698));
    Span4Mux_h I__2442 (
            .O(N__18718),
            .I(N__18695));
    InMux I__2441 (
            .O(N__18717),
            .I(N__18690));
    InMux I__2440 (
            .O(N__18716),
            .I(N__18690));
    LocalMux I__2439 (
            .O(N__18713),
            .I(N__18685));
    LocalMux I__2438 (
            .O(N__18710),
            .I(N__18685));
    LocalMux I__2437 (
            .O(N__18703),
            .I(\ALU.operand2_8 ));
    Odrv4 I__2436 (
            .O(N__18698),
            .I(\ALU.operand2_8 ));
    Odrv4 I__2435 (
            .O(N__18695),
            .I(\ALU.operand2_8 ));
    LocalMux I__2434 (
            .O(N__18690),
            .I(\ALU.operand2_8 ));
    Odrv12 I__2433 (
            .O(N__18685),
            .I(\ALU.operand2_8 ));
    CascadeMux I__2432 (
            .O(N__18674),
            .I(N__18670));
    InMux I__2431 (
            .O(N__18673),
            .I(N__18665));
    InMux I__2430 (
            .O(N__18670),
            .I(N__18662));
    CascadeMux I__2429 (
            .O(N__18669),
            .I(N__18659));
    CascadeMux I__2428 (
            .O(N__18668),
            .I(N__18656));
    LocalMux I__2427 (
            .O(N__18665),
            .I(N__18652));
    LocalMux I__2426 (
            .O(N__18662),
            .I(N__18649));
    InMux I__2425 (
            .O(N__18659),
            .I(N__18644));
    InMux I__2424 (
            .O(N__18656),
            .I(N__18641));
    InMux I__2423 (
            .O(N__18655),
            .I(N__18637));
    Span4Mux_h I__2422 (
            .O(N__18652),
            .I(N__18632));
    Span4Mux_v I__2421 (
            .O(N__18649),
            .I(N__18632));
    CascadeMux I__2420 (
            .O(N__18648),
            .I(N__18629));
    CascadeMux I__2419 (
            .O(N__18647),
            .I(N__18624));
    LocalMux I__2418 (
            .O(N__18644),
            .I(N__18619));
    LocalMux I__2417 (
            .O(N__18641),
            .I(N__18619));
    CascadeMux I__2416 (
            .O(N__18640),
            .I(N__18615));
    LocalMux I__2415 (
            .O(N__18637),
            .I(N__18609));
    Span4Mux_v I__2414 (
            .O(N__18632),
            .I(N__18609));
    InMux I__2413 (
            .O(N__18629),
            .I(N__18600));
    InMux I__2412 (
            .O(N__18628),
            .I(N__18600));
    InMux I__2411 (
            .O(N__18627),
            .I(N__18600));
    InMux I__2410 (
            .O(N__18624),
            .I(N__18600));
    Span4Mux_v I__2409 (
            .O(N__18619),
            .I(N__18597));
    InMux I__2408 (
            .O(N__18618),
            .I(N__18592));
    InMux I__2407 (
            .O(N__18615),
            .I(N__18592));
    InMux I__2406 (
            .O(N__18614),
            .I(N__18589));
    Span4Mux_v I__2405 (
            .O(N__18609),
            .I(N__18586));
    LocalMux I__2404 (
            .O(N__18600),
            .I(\ALU.N_199_0 ));
    Odrv4 I__2403 (
            .O(N__18597),
            .I(\ALU.N_199_0 ));
    LocalMux I__2402 (
            .O(N__18592),
            .I(\ALU.N_199_0 ));
    LocalMux I__2401 (
            .O(N__18589),
            .I(\ALU.N_199_0 ));
    Odrv4 I__2400 (
            .O(N__18586),
            .I(\ALU.N_199_0 ));
    InMux I__2399 (
            .O(N__18575),
            .I(N__18572));
    LocalMux I__2398 (
            .O(N__18572),
            .I(\ALU.a3_b_8 ));
    InMux I__2397 (
            .O(N__18569),
            .I(N__18566));
    LocalMux I__2396 (
            .O(N__18566),
            .I(N__18563));
    Span4Mux_v I__2395 (
            .O(N__18563),
            .I(N__18560));
    Odrv4 I__2394 (
            .O(N__18560),
            .I(\ALU.madd_275 ));
    InMux I__2393 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__2392 (
            .O(N__18554),
            .I(N__18551));
    Span4Mux_s3_h I__2391 (
            .O(N__18551),
            .I(N__18546));
    InMux I__2390 (
            .O(N__18550),
            .I(N__18541));
    InMux I__2389 (
            .O(N__18549),
            .I(N__18541));
    Span4Mux_h I__2388 (
            .O(N__18546),
            .I(N__18538));
    LocalMux I__2387 (
            .O(N__18541),
            .I(N__18535));
    Odrv4 I__2386 (
            .O(N__18538),
            .I(\ALU.madd_217 ));
    Odrv4 I__2385 (
            .O(N__18535),
            .I(\ALU.madd_217 ));
    CascadeMux I__2384 (
            .O(N__18530),
            .I(N__18527));
    InMux I__2383 (
            .O(N__18527),
            .I(N__18522));
    InMux I__2382 (
            .O(N__18526),
            .I(N__18519));
    InMux I__2381 (
            .O(N__18525),
            .I(N__18516));
    LocalMux I__2380 (
            .O(N__18522),
            .I(N__18512));
    LocalMux I__2379 (
            .O(N__18519),
            .I(N__18509));
    LocalMux I__2378 (
            .O(N__18516),
            .I(N__18506));
    CascadeMux I__2377 (
            .O(N__18515),
            .I(N__18503));
    Span4Mux_v I__2376 (
            .O(N__18512),
            .I(N__18497));
    Span4Mux_v I__2375 (
            .O(N__18509),
            .I(N__18497));
    Span4Mux_v I__2374 (
            .O(N__18506),
            .I(N__18494));
    InMux I__2373 (
            .O(N__18503),
            .I(N__18489));
    InMux I__2372 (
            .O(N__18502),
            .I(N__18489));
    Odrv4 I__2371 (
            .O(N__18497),
            .I(\ALU.madd_222 ));
    Odrv4 I__2370 (
            .O(N__18494),
            .I(\ALU.madd_222 ));
    LocalMux I__2369 (
            .O(N__18489),
            .I(\ALU.madd_222 ));
    InMux I__2368 (
            .O(N__18482),
            .I(N__18476));
    InMux I__2367 (
            .O(N__18481),
            .I(N__18476));
    LocalMux I__2366 (
            .O(N__18476),
            .I(N__18471));
    InMux I__2365 (
            .O(N__18475),
            .I(N__18466));
    InMux I__2364 (
            .O(N__18474),
            .I(N__18466));
    Span4Mux_h I__2363 (
            .O(N__18471),
            .I(N__18463));
    LocalMux I__2362 (
            .O(N__18466),
            .I(\ALU.madd_212 ));
    Odrv4 I__2361 (
            .O(N__18463),
            .I(\ALU.madd_212 ));
    InMux I__2360 (
            .O(N__18458),
            .I(N__18454));
    InMux I__2359 (
            .O(N__18457),
            .I(N__18451));
    LocalMux I__2358 (
            .O(N__18454),
            .I(N__18448));
    LocalMux I__2357 (
            .O(N__18451),
            .I(\ALU.madd_284 ));
    Odrv4 I__2356 (
            .O(N__18448),
            .I(\ALU.madd_284 ));
    CascadeMux I__2355 (
            .O(N__18443),
            .I(\ALU.madd_279_cascade_ ));
    CascadeMux I__2354 (
            .O(N__18440),
            .I(N__18437));
    InMux I__2353 (
            .O(N__18437),
            .I(N__18434));
    LocalMux I__2352 (
            .O(N__18434),
            .I(N__18431));
    Span4Mux_s3_h I__2351 (
            .O(N__18431),
            .I(N__18427));
    InMux I__2350 (
            .O(N__18430),
            .I(N__18424));
    Odrv4 I__2349 (
            .O(N__18427),
            .I(\ALU.madd_349 ));
    LocalMux I__2348 (
            .O(N__18424),
            .I(\ALU.madd_349 ));
    InMux I__2347 (
            .O(N__18419),
            .I(N__18415));
    InMux I__2346 (
            .O(N__18418),
            .I(N__18412));
    LocalMux I__2345 (
            .O(N__18415),
            .I(\ALU.d_RNIV96U8Z0Z_13 ));
    LocalMux I__2344 (
            .O(N__18412),
            .I(\ALU.d_RNIV96U8Z0Z_13 ));
    InMux I__2343 (
            .O(N__18407),
            .I(N__18404));
    LocalMux I__2342 (
            .O(N__18404),
            .I(N__18401));
    Span4Mux_h I__2341 (
            .O(N__18401),
            .I(N__18398));
    Span4Mux_h I__2340 (
            .O(N__18398),
            .I(N__18394));
    InMux I__2339 (
            .O(N__18397),
            .I(N__18391));
    Odrv4 I__2338 (
            .O(N__18394),
            .I(\ALU.madd_310_0 ));
    LocalMux I__2337 (
            .O(N__18391),
            .I(\ALU.madd_310_0 ));
    InMux I__2336 (
            .O(N__18386),
            .I(N__18383));
    LocalMux I__2335 (
            .O(N__18383),
            .I(\ALU.madd_330_0 ));
    CascadeMux I__2334 (
            .O(N__18380),
            .I(\ALU.c_RNIF549Z0Z_10_cascade_ ));
    InMux I__2333 (
            .O(N__18377),
            .I(N__18374));
    LocalMux I__2332 (
            .O(N__18374),
            .I(\ALU.a_RNIBLBOZ0Z_10 ));
    CascadeMux I__2331 (
            .O(N__18371),
            .I(\ALU.operand2_7_ns_1_10_cascade_ ));
    CascadeMux I__2330 (
            .O(N__18368),
            .I(\ALU.un9_addsub_axb_12_cascade_ ));
    CascadeMux I__2329 (
            .O(N__18365),
            .I(\ALU.d_RNIV96U8Z0Z_13_cascade_ ));
    InMux I__2328 (
            .O(N__18362),
            .I(N__18359));
    LocalMux I__2327 (
            .O(N__18359),
            .I(N__18355));
    InMux I__2326 (
            .O(N__18358),
            .I(N__18352));
    Odrv4 I__2325 (
            .O(N__18355),
            .I(\ALU.madd_314 ));
    LocalMux I__2324 (
            .O(N__18352),
            .I(\ALU.madd_314 ));
    CascadeMux I__2323 (
            .O(N__18347),
            .I(\ALU.madd_310_0_cascade_ ));
    InMux I__2322 (
            .O(N__18344),
            .I(N__18338));
    InMux I__2321 (
            .O(N__18343),
            .I(N__18338));
    LocalMux I__2320 (
            .O(N__18338),
            .I(\ALU.madd_334 ));
    InMux I__2319 (
            .O(N__18335),
            .I(N__18332));
    LocalMux I__2318 (
            .O(N__18332),
            .I(\ALU.a1_b_12 ));
    CascadeMux I__2317 (
            .O(N__18329),
            .I(\ALU.a2_b_9_cascade_ ));
    InMux I__2316 (
            .O(N__18326),
            .I(N__18323));
    LocalMux I__2315 (
            .O(N__18323),
            .I(\ALU.a9_b_4 ));
    CascadeMux I__2314 (
            .O(N__18320),
            .I(\ALU.a10_b_3_cascade_ ));
    InMux I__2313 (
            .O(N__18317),
            .I(N__18311));
    InMux I__2312 (
            .O(N__18316),
            .I(N__18311));
    LocalMux I__2311 (
            .O(N__18311),
            .I(\ALU.madd_319 ));
    InMux I__2310 (
            .O(N__18308),
            .I(N__18305));
    LocalMux I__2309 (
            .O(N__18305),
            .I(N__18302));
    Odrv4 I__2308 (
            .O(N__18302),
            .I(\ALU.madd_366 ));
    InMux I__2307 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__2306 (
            .O(N__18296),
            .I(\ALU.madd_484_11 ));
    InMux I__2305 (
            .O(N__18293),
            .I(N__18290));
    LocalMux I__2304 (
            .O(N__18290),
            .I(N__18287));
    Odrv4 I__2303 (
            .O(N__18287),
            .I(\ALU.madd_376 ));
    CascadeMux I__2302 (
            .O(N__18284),
            .I(\ALU.madd_484_17_cascade_ ));
    InMux I__2301 (
            .O(N__18281),
            .I(N__18278));
    LocalMux I__2300 (
            .O(N__18278),
            .I(\ALU.madd_484_15 ));
    InMux I__2299 (
            .O(N__18275),
            .I(N__18272));
    LocalMux I__2298 (
            .O(N__18272),
            .I(\ALU.madd_484_20 ));
    CascadeMux I__2297 (
            .O(N__18269),
            .I(N__18266));
    InMux I__2296 (
            .O(N__18266),
            .I(N__18262));
    InMux I__2295 (
            .O(N__18265),
            .I(N__18259));
    LocalMux I__2294 (
            .O(N__18262),
            .I(N__18256));
    LocalMux I__2293 (
            .O(N__18259),
            .I(N__18253));
    Span4Mux_h I__2292 (
            .O(N__18256),
            .I(N__18250));
    Odrv4 I__2291 (
            .O(N__18253),
            .I(\ALU.madd_309 ));
    Odrv4 I__2290 (
            .O(N__18250),
            .I(\ALU.madd_309 ));
    InMux I__2289 (
            .O(N__18245),
            .I(N__18242));
    LocalMux I__2288 (
            .O(N__18242),
            .I(N__18238));
    InMux I__2287 (
            .O(N__18241),
            .I(N__18235));
    Span4Mux_v I__2286 (
            .O(N__18238),
            .I(N__18232));
    LocalMux I__2285 (
            .O(N__18235),
            .I(N__18229));
    Span4Mux_s3_h I__2284 (
            .O(N__18232),
            .I(N__18226));
    Odrv12 I__2283 (
            .O(N__18229),
            .I(\ALU.madd_362 ));
    Odrv4 I__2282 (
            .O(N__18226),
            .I(\ALU.madd_362 ));
    InMux I__2281 (
            .O(N__18221),
            .I(N__18218));
    LocalMux I__2280 (
            .O(N__18218),
            .I(\ALU.madd_391 ));
    InMux I__2279 (
            .O(N__18215),
            .I(N__18212));
    LocalMux I__2278 (
            .O(N__18212),
            .I(N__18209));
    Span4Mux_h I__2277 (
            .O(N__18209),
            .I(N__18206));
    Odrv4 I__2276 (
            .O(N__18206),
            .I(\ALU.a5_b_9 ));
    InMux I__2275 (
            .O(N__18203),
            .I(N__18200));
    LocalMux I__2274 (
            .O(N__18200),
            .I(N__18197));
    Span4Mux_h I__2273 (
            .O(N__18197),
            .I(N__18193));
    InMux I__2272 (
            .O(N__18196),
            .I(N__18190));
    Odrv4 I__2271 (
            .O(N__18193),
            .I(\ALU.a6_b_8 ));
    LocalMux I__2270 (
            .O(N__18190),
            .I(\ALU.a6_b_8 ));
    CascadeMux I__2269 (
            .O(N__18185),
            .I(\ALU.a7_b_7_cascade_ ));
    InMux I__2268 (
            .O(N__18182),
            .I(N__18179));
    LocalMux I__2267 (
            .O(N__18179),
            .I(\ALU.madd_381 ));
    InMux I__2266 (
            .O(N__18176),
            .I(N__18173));
    LocalMux I__2265 (
            .O(N__18173),
            .I(\ALU.madd_484_16 ));
    CascadeMux I__2264 (
            .O(N__18170),
            .I(\ALU.dout_6_ns_1_12_cascade_ ));
    InMux I__2263 (
            .O(N__18167),
            .I(N__18164));
    LocalMux I__2262 (
            .O(N__18164),
            .I(\ALU.N_711 ));
    CascadeMux I__2261 (
            .O(N__18161),
            .I(\ALU.N_759_cascade_ ));
    CascadeMux I__2260 (
            .O(N__18158),
            .I(\ALU.aluOut_12_cascade_ ));
    CascadeMux I__2259 (
            .O(N__18155),
            .I(N__18152));
    InMux I__2258 (
            .O(N__18152),
            .I(N__18146));
    InMux I__2257 (
            .O(N__18151),
            .I(N__18146));
    LocalMux I__2256 (
            .O(N__18146),
            .I(\ALU.a12_b_2 ));
    InMux I__2255 (
            .O(N__18143),
            .I(N__18127));
    InMux I__2254 (
            .O(N__18142),
            .I(N__18127));
    InMux I__2253 (
            .O(N__18141),
            .I(N__18127));
    InMux I__2252 (
            .O(N__18140),
            .I(N__18127));
    InMux I__2251 (
            .O(N__18139),
            .I(N__18127));
    InMux I__2250 (
            .O(N__18138),
            .I(N__18124));
    LocalMux I__2249 (
            .O(N__18127),
            .I(N__18117));
    LocalMux I__2248 (
            .O(N__18124),
            .I(N__18114));
    InMux I__2247 (
            .O(N__18123),
            .I(N__18105));
    InMux I__2246 (
            .O(N__18122),
            .I(N__18105));
    InMux I__2245 (
            .O(N__18121),
            .I(N__18105));
    InMux I__2244 (
            .O(N__18120),
            .I(N__18105));
    Span4Mux_h I__2243 (
            .O(N__18117),
            .I(N__18101));
    Span4Mux_v I__2242 (
            .O(N__18114),
            .I(N__18098));
    LocalMux I__2241 (
            .O(N__18105),
            .I(N__18095));
    InMux I__2240 (
            .O(N__18104),
            .I(N__18092));
    Span4Mux_v I__2239 (
            .O(N__18101),
            .I(N__18087));
    Sp12to4 I__2238 (
            .O(N__18098),
            .I(N__18084));
    Span12Mux_h I__2237 (
            .O(N__18095),
            .I(N__18079));
    LocalMux I__2236 (
            .O(N__18092),
            .I(N__18079));
    InMux I__2235 (
            .O(N__18091),
            .I(N__18074));
    InMux I__2234 (
            .O(N__18090),
            .I(N__18074));
    Odrv4 I__2233 (
            .O(N__18087),
            .I(\ALU.N_90_0 ));
    Odrv12 I__2232 (
            .O(N__18084),
            .I(\ALU.N_90_0 ));
    Odrv12 I__2231 (
            .O(N__18079),
            .I(\ALU.N_90_0 ));
    LocalMux I__2230 (
            .O(N__18074),
            .I(\ALU.N_90_0 ));
    InMux I__2229 (
            .O(N__18065),
            .I(N__18062));
    LocalMux I__2228 (
            .O(N__18062),
            .I(N__18058));
    InMux I__2227 (
            .O(N__18061),
            .I(N__18055));
    Span4Mux_h I__2226 (
            .O(N__18058),
            .I(N__18049));
    LocalMux I__2225 (
            .O(N__18055),
            .I(N__18046));
    InMux I__2224 (
            .O(N__18054),
            .I(N__18039));
    InMux I__2223 (
            .O(N__18053),
            .I(N__18039));
    InMux I__2222 (
            .O(N__18052),
            .I(N__18039));
    Span4Mux_v I__2221 (
            .O(N__18049),
            .I(N__18034));
    Span4Mux_h I__2220 (
            .O(N__18046),
            .I(N__18034));
    LocalMux I__2219 (
            .O(N__18039),
            .I(ctrlOut_3));
    Odrv4 I__2218 (
            .O(N__18034),
            .I(ctrlOut_3));
    CascadeMux I__2217 (
            .O(N__18029),
            .I(\ALU.N_235_0_cascade_ ));
    CascadeMux I__2216 (
            .O(N__18026),
            .I(\ALU.a12_b_3_cascade_ ));
    CascadeMux I__2215 (
            .O(N__18023),
            .I(N__18019));
    InMux I__2214 (
            .O(N__18022),
            .I(N__18014));
    InMux I__2213 (
            .O(N__18019),
            .I(N__18014));
    LocalMux I__2212 (
            .O(N__18014),
            .I(ctrlOut_4));
    CascadeMux I__2211 (
            .O(N__18011),
            .I(\ALU.a_15_m2_ns_1Z0Z_14_cascade_ ));
    CascadeMux I__2210 (
            .O(N__18008),
            .I(\ALU.lshift_15_ns_1_14_cascade_ ));
    CascadeMux I__2209 (
            .O(N__18005),
            .I(\ALU.lshift_14_cascade_ ));
    InMux I__2208 (
            .O(N__18002),
            .I(N__17999));
    LocalMux I__2207 (
            .O(N__17999),
            .I(\ALU.a_15_m2_14 ));
    CascadeMux I__2206 (
            .O(N__17996),
            .I(\ALU.a_15_m4_14_cascade_ ));
    InMux I__2205 (
            .O(N__17993),
            .I(N__17990));
    LocalMux I__2204 (
            .O(N__17990),
            .I(N__17987));
    Odrv4 I__2203 (
            .O(N__17987),
            .I(\ALU.a_15_m3_14 ));
    CascadeMux I__2202 (
            .O(N__17984),
            .I(\ALU.dout_3_ns_1_12_cascade_ ));
    CascadeMux I__2201 (
            .O(N__17981),
            .I(\ALU.rshift_3_ns_1_6_cascade_ ));
    CascadeMux I__2200 (
            .O(N__17978),
            .I(\ALU.N_474_cascade_ ));
    InMux I__2199 (
            .O(N__17975),
            .I(N__17972));
    LocalMux I__2198 (
            .O(N__17972),
            .I(\ALU.rshift_15_ns_1_6 ));
    CascadeMux I__2197 (
            .O(N__17969),
            .I(\ALU.rshift_6_cascade_ ));
    InMux I__2196 (
            .O(N__17966),
            .I(N__17963));
    LocalMux I__2195 (
            .O(N__17963),
            .I(N__17960));
    Odrv4 I__2194 (
            .O(N__17960),
            .I(\ALU.N_291_0 ));
    CascadeMux I__2193 (
            .O(N__17957),
            .I(\ALU.dout_6_ns_1_14_cascade_ ));
    CascadeMux I__2192 (
            .O(N__17954),
            .I(\ALU.aluOut_15_cascade_ ));
    InMux I__2191 (
            .O(N__17951),
            .I(N__17948));
    LocalMux I__2190 (
            .O(N__17948),
            .I(\ALU.N_761 ));
    InMux I__2189 (
            .O(N__17945),
            .I(N__17942));
    LocalMux I__2188 (
            .O(N__17942),
            .I(\ALU.N_713 ));
    InMux I__2187 (
            .O(N__17939),
            .I(N__17930));
    InMux I__2186 (
            .O(N__17938),
            .I(N__17930));
    InMux I__2185 (
            .O(N__17937),
            .I(N__17930));
    LocalMux I__2184 (
            .O(N__17930),
            .I(\ALU.a_cnv_0Z0Z_0 ));
    CascadeMux I__2183 (
            .O(N__17927),
            .I(N__17918));
    InMux I__2182 (
            .O(N__17926),
            .I(N__17914));
    InMux I__2181 (
            .O(N__17925),
            .I(N__17911));
    InMux I__2180 (
            .O(N__17924),
            .I(N__17908));
    InMux I__2179 (
            .O(N__17923),
            .I(N__17897));
    InMux I__2178 (
            .O(N__17922),
            .I(N__17897));
    InMux I__2177 (
            .O(N__17921),
            .I(N__17897));
    InMux I__2176 (
            .O(N__17918),
            .I(N__17897));
    InMux I__2175 (
            .O(N__17917),
            .I(N__17897));
    LocalMux I__2174 (
            .O(N__17914),
            .I(aluResults_1));
    LocalMux I__2173 (
            .O(N__17911),
            .I(aluResults_1));
    LocalMux I__2172 (
            .O(N__17908),
            .I(aluResults_1));
    LocalMux I__2171 (
            .O(N__17897),
            .I(aluResults_1));
    CascadeMux I__2170 (
            .O(N__17888),
            .I(N__17885));
    InMux I__2169 (
            .O(N__17885),
            .I(N__17879));
    CascadeMux I__2168 (
            .O(N__17884),
            .I(N__17876));
    CascadeMux I__2167 (
            .O(N__17883),
            .I(N__17873));
    InMux I__2166 (
            .O(N__17882),
            .I(N__17870));
    LocalMux I__2165 (
            .O(N__17879),
            .I(N__17867));
    InMux I__2164 (
            .O(N__17876),
            .I(N__17862));
    InMux I__2163 (
            .O(N__17873),
            .I(N__17862));
    LocalMux I__2162 (
            .O(N__17870),
            .I(\ALU.b_cnv_0Z0Z_0 ));
    Odrv4 I__2161 (
            .O(N__17867),
            .I(\ALU.b_cnv_0Z0Z_0 ));
    LocalMux I__2160 (
            .O(N__17862),
            .I(\ALU.b_cnv_0Z0Z_0 ));
    CascadeMux I__2159 (
            .O(N__17855),
            .I(N__17849));
    CascadeMux I__2158 (
            .O(N__17854),
            .I(N__17844));
    CascadeMux I__2157 (
            .O(N__17853),
            .I(N__17841));
    InMux I__2156 (
            .O(N__17852),
            .I(N__17836));
    InMux I__2155 (
            .O(N__17849),
            .I(N__17823));
    InMux I__2154 (
            .O(N__17848),
            .I(N__17823));
    InMux I__2153 (
            .O(N__17847),
            .I(N__17823));
    InMux I__2152 (
            .O(N__17844),
            .I(N__17823));
    InMux I__2151 (
            .O(N__17841),
            .I(N__17823));
    InMux I__2150 (
            .O(N__17840),
            .I(N__17823));
    InMux I__2149 (
            .O(N__17839),
            .I(N__17820));
    LocalMux I__2148 (
            .O(N__17836),
            .I(aluResults_2));
    LocalMux I__2147 (
            .O(N__17823),
            .I(aluResults_2));
    LocalMux I__2146 (
            .O(N__17820),
            .I(aluResults_2));
    InMux I__2145 (
            .O(N__17813),
            .I(N__17808));
    InMux I__2144 (
            .O(N__17812),
            .I(N__17803));
    InMux I__2143 (
            .O(N__17811),
            .I(N__17803));
    LocalMux I__2142 (
            .O(N__17808),
            .I(N__17799));
    LocalMux I__2141 (
            .O(N__17803),
            .I(N__17796));
    InMux I__2140 (
            .O(N__17802),
            .I(N__17793));
    Odrv4 I__2139 (
            .O(N__17799),
            .I(\ALU.N_169_0 ));
    Odrv4 I__2138 (
            .O(N__17796),
            .I(\ALU.N_169_0 ));
    LocalMux I__2137 (
            .O(N__17793),
            .I(\ALU.N_169_0 ));
    CascadeMux I__2136 (
            .O(N__17786),
            .I(\ALU.c_RNIEP354Z0Z_14_cascade_ ));
    InMux I__2135 (
            .O(N__17783),
            .I(N__17780));
    LocalMux I__2134 (
            .O(N__17780),
            .I(\ALU.c_RNIJENJ8_0Z0Z_15 ));
    CascadeMux I__2133 (
            .O(N__17777),
            .I(testClock_0_cascade_));
    CascadeMux I__2132 (
            .O(N__17774),
            .I(\ALU.a_cnv_0Z0Z_0_cascade_ ));
    InMux I__2131 (
            .O(N__17771),
            .I(N__17768));
    LocalMux I__2130 (
            .O(N__17768),
            .I(\ALU.N_53_0 ));
    InMux I__2129 (
            .O(N__17765),
            .I(N__17759));
    InMux I__2128 (
            .O(N__17764),
            .I(N__17759));
    LocalMux I__2127 (
            .O(N__17759),
            .I(N__17756));
    Odrv4 I__2126 (
            .O(N__17756),
            .I(aluResults_0));
    InMux I__2125 (
            .O(N__17753),
            .I(N__17750));
    LocalMux I__2124 (
            .O(N__17750),
            .I(testClock_0));
    InMux I__2123 (
            .O(N__17747),
            .I(N__17740));
    InMux I__2122 (
            .O(N__17746),
            .I(N__17731));
    InMux I__2121 (
            .O(N__17745),
            .I(N__17731));
    InMux I__2120 (
            .O(N__17744),
            .I(N__17731));
    InMux I__2119 (
            .O(N__17743),
            .I(N__17731));
    LocalMux I__2118 (
            .O(N__17740),
            .I(testClockZ0));
    LocalMux I__2117 (
            .O(N__17731),
            .I(testClockZ0));
    CascadeMux I__2116 (
            .O(N__17726),
            .I(\ALU.madd_41_cascade_ ));
    CascadeMux I__2115 (
            .O(N__17723),
            .I(\ALU.madd_46_cascade_ ));
    CascadeMux I__2114 (
            .O(N__17720),
            .I(\ALU.madd_39_cascade_ ));
    InMux I__2113 (
            .O(N__17717),
            .I(N__17711));
    InMux I__2112 (
            .O(N__17716),
            .I(N__17711));
    LocalMux I__2111 (
            .O(N__17711),
            .I(N__17708));
    Odrv4 I__2110 (
            .O(N__17708),
            .I(\ALU.a6_b_3 ));
    CascadeMux I__2109 (
            .O(N__17705),
            .I(\ALU.madd_78_0_tz_cascade_ ));
    InMux I__2108 (
            .O(N__17702),
            .I(N__17699));
    LocalMux I__2107 (
            .O(N__17699),
            .I(\ALU.madd_78_0 ));
    InMux I__2106 (
            .O(N__17696),
            .I(N__17693));
    LocalMux I__2105 (
            .O(N__17693),
            .I(\ALU.madd_39 ));
    CascadeMux I__2104 (
            .O(N__17690),
            .I(\ALU.madd_78_0_cascade_ ));
    CascadeMux I__2103 (
            .O(N__17687),
            .I(\ALU.madd_114_cascade_ ));
    CascadeMux I__2102 (
            .O(N__17684),
            .I(\ALU.g1_2_cascade_ ));
    InMux I__2101 (
            .O(N__17681),
            .I(N__17678));
    LocalMux I__2100 (
            .O(N__17678),
            .I(\ALU.a4_b_0_7 ));
    InMux I__2099 (
            .O(N__17675),
            .I(N__17672));
    LocalMux I__2098 (
            .O(N__17672),
            .I(N__17669));
    Odrv4 I__2097 (
            .O(N__17669),
            .I(\ALU.g2_0_0_0 ));
    CascadeMux I__2096 (
            .O(N__17666),
            .I(\ALU.un2_addsub_axb_5_cascade_ ));
    InMux I__2095 (
            .O(N__17663),
            .I(N__17660));
    LocalMux I__2094 (
            .O(N__17660),
            .I(N__17657));
    Span4Mux_v I__2093 (
            .O(N__17657),
            .I(N__17654));
    Odrv4 I__2092 (
            .O(N__17654),
            .I(\ALU.a6_b_0_7 ));
    CascadeMux I__2091 (
            .O(N__17651),
            .I(\ALU.a6_b_0_cascade_ ));
    InMux I__2090 (
            .O(N__17648),
            .I(N__17642));
    InMux I__2089 (
            .O(N__17647),
            .I(N__17642));
    LocalMux I__2088 (
            .O(N__17642),
            .I(\ALU.madd_275_0 ));
    CascadeMux I__2087 (
            .O(N__17639),
            .I(\ALU.madd_42_cascade_ ));
    InMux I__2086 (
            .O(N__17636),
            .I(N__17633));
    LocalMux I__2085 (
            .O(N__17633),
            .I(\ALU.madd_42_0 ));
    CascadeMux I__2084 (
            .O(N__17630),
            .I(\ALU.e_RNIM09HZ0Z_7_cascade_ ));
    CascadeMux I__2083 (
            .O(N__17627),
            .I(\ALU.operand2_7_ns_1_7_cascade_ ));
    InMux I__2082 (
            .O(N__17624),
            .I(N__17621));
    LocalMux I__2081 (
            .O(N__17621),
            .I(N__17618));
    Span4Mux_v I__2080 (
            .O(N__17618),
            .I(N__17615));
    Odrv4 I__2079 (
            .O(N__17615),
            .I(\ALU.a2_b_6 ));
    InMux I__2078 (
            .O(N__17612),
            .I(N__17609));
    LocalMux I__2077 (
            .O(N__17609),
            .I(N__17606));
    Span4Mux_v I__2076 (
            .O(N__17606),
            .I(N__17603));
    Odrv4 I__2075 (
            .O(N__17603),
            .I(\ALU.a0_b_8 ));
    CascadeMux I__2074 (
            .O(N__17600),
            .I(\ALU.a2_b_6_cascade_ ));
    CascadeMux I__2073 (
            .O(N__17597),
            .I(\ALU.a5_b_6_cascade_ ));
    CascadeMux I__2072 (
            .O(N__17594),
            .I(\ALU.operand2_5_cascade_ ));
    InMux I__2071 (
            .O(N__17591),
            .I(N__17585));
    InMux I__2070 (
            .O(N__17590),
            .I(N__17585));
    LocalMux I__2069 (
            .O(N__17585),
            .I(N__17582));
    Span4Mux_v I__2068 (
            .O(N__17582),
            .I(N__17579));
    Odrv4 I__2067 (
            .O(N__17579),
            .I(\ALU.madd_176_0 ));
    InMux I__2066 (
            .O(N__17576),
            .I(N__17570));
    InMux I__2065 (
            .O(N__17575),
            .I(N__17570));
    LocalMux I__2064 (
            .O(N__17570),
            .I(N__17567));
    Span4Mux_v I__2063 (
            .O(N__17567),
            .I(N__17563));
    InMux I__2062 (
            .O(N__17566),
            .I(N__17560));
    Odrv4 I__2061 (
            .O(N__17563),
            .I(\ALU.madd_218_0 ));
    LocalMux I__2060 (
            .O(N__17560),
            .I(\ALU.madd_218_0 ));
    InMux I__2059 (
            .O(N__17555),
            .I(N__17551));
    InMux I__2058 (
            .O(N__17554),
            .I(N__17548));
    LocalMux I__2057 (
            .O(N__17551),
            .I(\ALU.a7_b_4 ));
    LocalMux I__2056 (
            .O(N__17548),
            .I(\ALU.a7_b_4 ));
    InMux I__2055 (
            .O(N__17543),
            .I(N__17540));
    LocalMux I__2054 (
            .O(N__17540),
            .I(N__17537));
    Span4Mux_s1_h I__2053 (
            .O(N__17537),
            .I(N__17534));
    Span4Mux_v I__2052 (
            .O(N__17534),
            .I(N__17529));
    InMux I__2051 (
            .O(N__17533),
            .I(N__17526));
    InMux I__2050 (
            .O(N__17532),
            .I(N__17523));
    Odrv4 I__2049 (
            .O(N__17529),
            .I(\ALU.a6_b_5 ));
    LocalMux I__2048 (
            .O(N__17526),
            .I(\ALU.a6_b_5 ));
    LocalMux I__2047 (
            .O(N__17523),
            .I(\ALU.a6_b_5 ));
    InMux I__2046 (
            .O(N__17516),
            .I(N__17513));
    LocalMux I__2045 (
            .O(N__17513),
            .I(N__17510));
    Span4Mux_s2_h I__2044 (
            .O(N__17510),
            .I(N__17506));
    CascadeMux I__2043 (
            .O(N__17509),
            .I(N__17503));
    Span4Mux_h I__2042 (
            .O(N__17506),
            .I(N__17500));
    InMux I__2041 (
            .O(N__17503),
            .I(N__17497));
    Odrv4 I__2040 (
            .O(N__17500),
            .I(\ALU.a5_b_6 ));
    LocalMux I__2039 (
            .O(N__17497),
            .I(\ALU.a5_b_6 ));
    CascadeMux I__2038 (
            .O(N__17492),
            .I(N__17487));
    InMux I__2037 (
            .O(N__17491),
            .I(N__17484));
    InMux I__2036 (
            .O(N__17490),
            .I(N__17481));
    InMux I__2035 (
            .O(N__17487),
            .I(N__17478));
    LocalMux I__2034 (
            .O(N__17484),
            .I(N__17475));
    LocalMux I__2033 (
            .O(N__17481),
            .I(N__17472));
    LocalMux I__2032 (
            .O(N__17478),
            .I(N__17469));
    Span12Mux_s2_h I__2031 (
            .O(N__17475),
            .I(N__17466));
    Span4Mux_v I__2030 (
            .O(N__17472),
            .I(N__17461));
    Span4Mux_s2_h I__2029 (
            .O(N__17469),
            .I(N__17461));
    Odrv12 I__2028 (
            .O(N__17466),
            .I(\ALU.madd_320 ));
    Odrv4 I__2027 (
            .O(N__17461),
            .I(\ALU.madd_320 ));
    InMux I__2026 (
            .O(N__17456),
            .I(N__17451));
    InMux I__2025 (
            .O(N__17455),
            .I(N__17448));
    InMux I__2024 (
            .O(N__17454),
            .I(N__17445));
    LocalMux I__2023 (
            .O(N__17451),
            .I(\ALU.madd_325_0 ));
    LocalMux I__2022 (
            .O(N__17448),
            .I(\ALU.madd_325_0 ));
    LocalMux I__2021 (
            .O(N__17445),
            .I(\ALU.madd_325_0 ));
    CascadeMux I__2020 (
            .O(N__17438),
            .I(\ALU.madd_274_cascade_ ));
    InMux I__2019 (
            .O(N__17435),
            .I(N__17432));
    LocalMux I__2018 (
            .O(N__17432),
            .I(N__17428));
    InMux I__2017 (
            .O(N__17431),
            .I(N__17425));
    Span4Mux_v I__2016 (
            .O(N__17428),
            .I(N__17422));
    LocalMux I__2015 (
            .O(N__17425),
            .I(N__17419));
    Odrv4 I__2014 (
            .O(N__17422),
            .I(\ALU.madd_254 ));
    Odrv4 I__2013 (
            .O(N__17419),
            .I(\ALU.madd_254 ));
    InMux I__2012 (
            .O(N__17414),
            .I(N__17411));
    LocalMux I__2011 (
            .O(N__17411),
            .I(N__17408));
    Span4Mux_s2_h I__2010 (
            .O(N__17408),
            .I(N__17404));
    InMux I__2009 (
            .O(N__17407),
            .I(N__17401));
    Odrv4 I__2008 (
            .O(N__17404),
            .I(\ALU.madd_344 ));
    LocalMux I__2007 (
            .O(N__17401),
            .I(\ALU.madd_344 ));
    CascadeMux I__2006 (
            .O(N__17396),
            .I(\ALU.madd_29_cascade_ ));
    CascadeMux I__2005 (
            .O(N__17393),
            .I(\ALU.madd_47_cascade_ ));
    InMux I__2004 (
            .O(N__17390),
            .I(N__17387));
    LocalMux I__2003 (
            .O(N__17387),
            .I(N__17384));
    Odrv4 I__2002 (
            .O(N__17384),
            .I(\ALU.madd_265_0 ));
    CascadeMux I__2001 (
            .O(N__17381),
            .I(N__17377));
    InMux I__2000 (
            .O(N__17380),
            .I(N__17374));
    InMux I__1999 (
            .O(N__17377),
            .I(N__17371));
    LocalMux I__1998 (
            .O(N__17374),
            .I(N__17368));
    LocalMux I__1997 (
            .O(N__17371),
            .I(N__17365));
    Span12Mux_h I__1996 (
            .O(N__17368),
            .I(N__17362));
    Span4Mux_v I__1995 (
            .O(N__17365),
            .I(N__17359));
    Odrv12 I__1994 (
            .O(N__17362),
            .I(\ALU.madd_260 ));
    Odrv4 I__1993 (
            .O(N__17359),
            .I(\ALU.madd_260 ));
    InMux I__1992 (
            .O(N__17354),
            .I(N__17348));
    InMux I__1991 (
            .O(N__17353),
            .I(N__17348));
    LocalMux I__1990 (
            .O(N__17348),
            .I(\ALU.madd_329 ));
    InMux I__1989 (
            .O(N__17345),
            .I(N__17339));
    InMux I__1988 (
            .O(N__17344),
            .I(N__17339));
    LocalMux I__1987 (
            .O(N__17339),
            .I(\ALU.madd_407 ));
    InMux I__1986 (
            .O(N__17336),
            .I(N__17333));
    LocalMux I__1985 (
            .O(N__17333),
            .I(\ALU.madd_412 ));
    InMux I__1984 (
            .O(N__17330),
            .I(N__17327));
    LocalMux I__1983 (
            .O(N__17327),
            .I(\ALU.madd_i3_mux_1 ));
    InMux I__1982 (
            .O(N__17324),
            .I(N__17321));
    LocalMux I__1981 (
            .O(N__17321),
            .I(\ALU.madd_330 ));
    CascadeMux I__1980 (
            .O(N__17318),
            .I(N__17315));
    InMux I__1979 (
            .O(N__17315),
            .I(N__17312));
    LocalMux I__1978 (
            .O(N__17312),
            .I(N__17309));
    Span4Mux_v I__1977 (
            .O(N__17309),
            .I(N__17306));
    Span4Mux_s0_h I__1976 (
            .O(N__17306),
            .I(N__17303));
    Odrv4 I__1975 (
            .O(N__17303),
            .I(\ALU.madd_141_1 ));
    CascadeMux I__1974 (
            .O(N__17300),
            .I(N__17296));
    InMux I__1973 (
            .O(N__17299),
            .I(N__17291));
    InMux I__1972 (
            .O(N__17296),
            .I(N__17284));
    InMux I__1971 (
            .O(N__17295),
            .I(N__17284));
    InMux I__1970 (
            .O(N__17294),
            .I(N__17284));
    LocalMux I__1969 (
            .O(N__17291),
            .I(\ALU.madd_270_0 ));
    LocalMux I__1968 (
            .O(N__17284),
            .I(\ALU.madd_270_0 ));
    InMux I__1967 (
            .O(N__17279),
            .I(N__17276));
    LocalMux I__1966 (
            .O(N__17276),
            .I(\ALU.madd_250_0 ));
    CascadeMux I__1965 (
            .O(N__17273),
            .I(\ALU.madd_250_0_cascade_ ));
    CascadeMux I__1964 (
            .O(N__17270),
            .I(N__17267));
    InMux I__1963 (
            .O(N__17267),
            .I(N__17264));
    LocalMux I__1962 (
            .O(N__17264),
            .I(N__17261));
    Span4Mux_v I__1961 (
            .O(N__17261),
            .I(N__17258));
    Span4Mux_s0_h I__1960 (
            .O(N__17258),
            .I(N__17255));
    Odrv4 I__1959 (
            .O(N__17255),
            .I(\ALU.madd_250 ));
    CascadeMux I__1958 (
            .O(N__17252),
            .I(N__17247));
    InMux I__1957 (
            .O(N__17251),
            .I(N__17244));
    InMux I__1956 (
            .O(N__17250),
            .I(N__17239));
    InMux I__1955 (
            .O(N__17247),
            .I(N__17239));
    LocalMux I__1954 (
            .O(N__17244),
            .I(N__17236));
    LocalMux I__1953 (
            .O(N__17239),
            .I(N__17233));
    Odrv4 I__1952 (
            .O(N__17236),
            .I(\ALU.a3_b_9 ));
    Odrv4 I__1951 (
            .O(N__17233),
            .I(\ALU.a3_b_9 ));
    CascadeMux I__1950 (
            .O(N__17228),
            .I(\ALU.madd_250_cascade_ ));
    InMux I__1949 (
            .O(N__17225),
            .I(N__17221));
    InMux I__1948 (
            .O(N__17224),
            .I(N__17218));
    LocalMux I__1947 (
            .O(N__17221),
            .I(N__17215));
    LocalMux I__1946 (
            .O(N__17218),
            .I(N__17208));
    Span4Mux_s2_h I__1945 (
            .O(N__17215),
            .I(N__17205));
    InMux I__1944 (
            .O(N__17214),
            .I(N__17198));
    InMux I__1943 (
            .O(N__17213),
            .I(N__17198));
    InMux I__1942 (
            .O(N__17212),
            .I(N__17198));
    InMux I__1941 (
            .O(N__17211),
            .I(N__17195));
    Odrv4 I__1940 (
            .O(N__17208),
            .I(\ALU.madd_207 ));
    Odrv4 I__1939 (
            .O(N__17205),
            .I(\ALU.madd_207 ));
    LocalMux I__1938 (
            .O(N__17198),
            .I(\ALU.madd_207 ));
    LocalMux I__1937 (
            .O(N__17195),
            .I(\ALU.madd_207 ));
    InMux I__1936 (
            .O(N__17186),
            .I(N__17180));
    InMux I__1935 (
            .O(N__17185),
            .I(N__17180));
    LocalMux I__1934 (
            .O(N__17180),
            .I(\ALU.madd_274 ));
    InMux I__1933 (
            .O(N__17177),
            .I(N__17174));
    LocalMux I__1932 (
            .O(N__17174),
            .I(\ALU.madd_372_0 ));
    InMux I__1931 (
            .O(N__17171),
            .I(N__17165));
    InMux I__1930 (
            .O(N__17170),
            .I(N__17165));
    LocalMux I__1929 (
            .O(N__17165),
            .I(\ALU.madd_382 ));
    CascadeMux I__1928 (
            .O(N__17162),
            .I(\ALU.madd_377_cascade_ ));
    InMux I__1927 (
            .O(N__17159),
            .I(N__17156));
    LocalMux I__1926 (
            .O(N__17156),
            .I(N__17152));
    InMux I__1925 (
            .O(N__17155),
            .I(N__17149));
    Odrv4 I__1924 (
            .O(N__17152),
            .I(\ALU.a13_b_1 ));
    LocalMux I__1923 (
            .O(N__17149),
            .I(\ALU.a13_b_1 ));
    InMux I__1922 (
            .O(N__17144),
            .I(N__17141));
    LocalMux I__1921 (
            .O(N__17141),
            .I(\ALU.madd_397 ));
    InMux I__1920 (
            .O(N__17138),
            .I(N__17132));
    InMux I__1919 (
            .O(N__17137),
            .I(N__17132));
    LocalMux I__1918 (
            .O(N__17132),
            .I(\ALU.madd_392 ));
    CascadeMux I__1917 (
            .O(N__17129),
            .I(\ALU.madd_397_cascade_ ));
    InMux I__1916 (
            .O(N__17126),
            .I(N__17120));
    InMux I__1915 (
            .O(N__17125),
            .I(N__17120));
    LocalMux I__1914 (
            .O(N__17120),
            .I(N__17117));
    Odrv4 I__1913 (
            .O(N__17117),
            .I(\ALU.madd_339 ));
    InMux I__1912 (
            .O(N__17114),
            .I(N__17111));
    LocalMux I__1911 (
            .O(N__17111),
            .I(\ALU.madd_406 ));
    CascadeMux I__1910 (
            .O(N__17108),
            .I(\ALU.a5_b_8_cascade_ ));
    InMux I__1909 (
            .O(N__17105),
            .I(N__17102));
    LocalMux I__1908 (
            .O(N__17102),
            .I(\ALU.madd_387 ));
    InMux I__1907 (
            .O(N__17099),
            .I(N__17093));
    InMux I__1906 (
            .O(N__17098),
            .I(N__17093));
    LocalMux I__1905 (
            .O(N__17093),
            .I(\ALU.madd_329_0 ));
    CascadeMux I__1904 (
            .O(N__17090),
            .I(\ALU.madd_387_cascade_ ));
    InMux I__1903 (
            .O(N__17087),
            .I(N__17084));
    LocalMux I__1902 (
            .O(N__17084),
            .I(\ALU.madd_402 ));
    CascadeMux I__1901 (
            .O(N__17081),
            .I(\ALU.madd_402_cascade_ ));
    InMux I__1900 (
            .O(N__17078),
            .I(N__17075));
    LocalMux I__1899 (
            .O(N__17075),
            .I(\ALU.madd_354 ));
    CascadeMux I__1898 (
            .O(N__17072),
            .I(\ALU.madd_412_cascade_ ));
    CascadeMux I__1897 (
            .O(N__17069),
            .I(\ALU.madd_324_0_cascade_ ));
    InMux I__1896 (
            .O(N__17066),
            .I(N__17063));
    LocalMux I__1895 (
            .O(N__17063),
            .I(N__17060));
    Odrv4 I__1894 (
            .O(N__17060),
            .I(\ALU.madd_372 ));
    InMux I__1893 (
            .O(N__17057),
            .I(N__17054));
    LocalMux I__1892 (
            .O(N__17054),
            .I(\ALU.madd_396 ));
    InMux I__1891 (
            .O(N__17051),
            .I(N__17048));
    LocalMux I__1890 (
            .O(N__17048),
            .I(\ALU.madd_484_21 ));
    CascadeMux I__1889 (
            .O(N__17045),
            .I(\ALU.madd_411_cascade_ ));
    InMux I__1888 (
            .O(N__17042),
            .I(N__17039));
    LocalMux I__1887 (
            .O(N__17039),
            .I(\ALU.madd_484_24 ));
    CascadeMux I__1886 (
            .O(N__17036),
            .I(N__17032));
    InMux I__1885 (
            .O(N__17035),
            .I(N__17027));
    InMux I__1884 (
            .O(N__17032),
            .I(N__17027));
    LocalMux I__1883 (
            .O(N__17027),
            .I(\ALU.a8_b_6 ));
    InMux I__1882 (
            .O(N__17024),
            .I(N__17018));
    InMux I__1881 (
            .O(N__17023),
            .I(N__17018));
    LocalMux I__1880 (
            .O(N__17018),
            .I(\ALU.a9_b_5 ));
    CascadeMux I__1879 (
            .O(N__17015),
            .I(N__17012));
    InMux I__1878 (
            .O(N__17012),
            .I(N__17009));
    LocalMux I__1877 (
            .O(N__17009),
            .I(\ALU.madd_377 ));
    InMux I__1876 (
            .O(N__17006),
            .I(N__17003));
    LocalMux I__1875 (
            .O(N__17003),
            .I(\ALU.a11_b_3 ));
    CascadeMux I__1874 (
            .O(N__17000),
            .I(\ALU.a11_b_3_cascade_ ));
    CascadeMux I__1873 (
            .O(N__16997),
            .I(N__16993));
    InMux I__1872 (
            .O(N__16996),
            .I(N__16988));
    InMux I__1871 (
            .O(N__16993),
            .I(N__16988));
    LocalMux I__1870 (
            .O(N__16988),
            .I(ctrlOut_14));
    InMux I__1869 (
            .O(N__16985),
            .I(N__16982));
    LocalMux I__1868 (
            .O(N__16982),
            .I(N__16977));
    InMux I__1867 (
            .O(N__16981),
            .I(N__16972));
    InMux I__1866 (
            .O(N__16980),
            .I(N__16972));
    Span4Mux_v I__1865 (
            .O(N__16977),
            .I(N__16967));
    LocalMux I__1864 (
            .O(N__16972),
            .I(N__16967));
    Span4Mux_h I__1863 (
            .O(N__16967),
            .I(N__16963));
    InMux I__1862 (
            .O(N__16966),
            .I(N__16960));
    Span4Mux_s0_h I__1861 (
            .O(N__16963),
            .I(N__16957));
    LocalMux I__1860 (
            .O(N__16960),
            .I(RXbuffer_6));
    Odrv4 I__1859 (
            .O(N__16957),
            .I(RXbuffer_6));
    InMux I__1858 (
            .O(N__16952),
            .I(N__16949));
    LocalMux I__1857 (
            .O(N__16949),
            .I(N__16945));
    CascadeMux I__1856 (
            .O(N__16948),
            .I(N__16942));
    Span4Mux_s2_v I__1855 (
            .O(N__16945),
            .I(N__16939));
    InMux I__1854 (
            .O(N__16942),
            .I(N__16936));
    Odrv4 I__1853 (
            .O(N__16939),
            .I(testWordZ0Z_14));
    LocalMux I__1852 (
            .O(N__16936),
            .I(testWordZ0Z_14));
    CascadeMux I__1851 (
            .O(N__16931),
            .I(\ALU.a7_b_6_cascade_ ));
    InMux I__1850 (
            .O(N__16928),
            .I(N__16922));
    InMux I__1849 (
            .O(N__16927),
            .I(N__16922));
    LocalMux I__1848 (
            .O(N__16922),
            .I(\ALU.a6_b_7 ));
    CascadeMux I__1847 (
            .O(N__16919),
            .I(N__16916));
    InMux I__1846 (
            .O(N__16916),
            .I(N__16913));
    LocalMux I__1845 (
            .O(N__16913),
            .I(\ALU.a7_b_6 ));
    InMux I__1844 (
            .O(N__16910),
            .I(N__16907));
    LocalMux I__1843 (
            .O(N__16907),
            .I(\ALU.madd_324_0 ));
    CascadeMux I__1842 (
            .O(N__16904),
            .I(\ALU.a13_b_1_cascade_ ));
    InMux I__1841 (
            .O(N__16901),
            .I(N__16898));
    LocalMux I__1840 (
            .O(N__16898),
            .I(\ALU.un2_addsub_axb_14 ));
    CascadeMux I__1839 (
            .O(N__16895),
            .I(\ALU.un2_addsub_axb_9_cascade_ ));
    CascadeMux I__1838 (
            .O(N__16892),
            .I(N_662_0_cascade_));
    InMux I__1837 (
            .O(N__16889),
            .I(N__16886));
    LocalMux I__1836 (
            .O(N__16886),
            .I(N_665_0));
    CascadeMux I__1835 (
            .O(N__16883),
            .I(N_301_0_cascade_));
    CascadeMux I__1834 (
            .O(N__16880),
            .I(N_668_0_cascade_));
    InMux I__1833 (
            .O(N__16877),
            .I(N__16874));
    LocalMux I__1832 (
            .O(N__16874),
            .I(\ALU.m300_nsZ0Z_1 ));
    InMux I__1831 (
            .O(N__16871),
            .I(N__16868));
    LocalMux I__1830 (
            .O(N__16868),
            .I(N__16865));
    Span4Mux_v I__1829 (
            .O(N__16865),
            .I(N__16860));
    InMux I__1828 (
            .O(N__16864),
            .I(N__16855));
    InMux I__1827 (
            .O(N__16863),
            .I(N__16855));
    Odrv4 I__1826 (
            .O(N__16860),
            .I(N_662_0));
    LocalMux I__1825 (
            .O(N__16855),
            .I(N_662_0));
    CascadeMux I__1824 (
            .O(N__16850),
            .I(N_670_0_cascade_));
    CEMux I__1823 (
            .O(N__16847),
            .I(N__16844));
    LocalMux I__1822 (
            .O(N__16844),
            .I(N__16840));
    CEMux I__1821 (
            .O(N__16843),
            .I(N__16837));
    Span4Mux_s2_v I__1820 (
            .O(N__16840),
            .I(N__16834));
    LocalMux I__1819 (
            .O(N__16837),
            .I(N__16831));
    Sp12to4 I__1818 (
            .O(N__16834),
            .I(N__16828));
    Span4Mux_h I__1817 (
            .O(N__16831),
            .I(N__16825));
    Odrv12 I__1816 (
            .O(N__16828),
            .I(\CONTROL.results_cnvZ0Z_0 ));
    Odrv4 I__1815 (
            .O(N__16825),
            .I(\CONTROL.results_cnvZ0Z_0 ));
    CascadeMux I__1814 (
            .O(N__16820),
            .I(N_51_0_cascade_));
    InMux I__1813 (
            .O(N__16817),
            .I(N__16814));
    LocalMux I__1812 (
            .O(N__16814),
            .I(N__16811));
    IoSpan4Mux I__1811 (
            .O(N__16811),
            .I(N__16807));
    InMux I__1810 (
            .O(N__16810),
            .I(N__16804));
    IoSpan4Mux I__1809 (
            .O(N__16807),
            .I(N__16799));
    LocalMux I__1808 (
            .O(N__16804),
            .I(N__16799));
    Odrv4 I__1807 (
            .O(N__16799),
            .I(testWordZ0Z_15));
    InMux I__1806 (
            .O(N__16796),
            .I(N__16793));
    LocalMux I__1805 (
            .O(N__16793),
            .I(N__16789));
    InMux I__1804 (
            .O(N__16792),
            .I(N__16786));
    Odrv4 I__1803 (
            .O(N__16789),
            .I(\ALU.madd_129 ));
    LocalMux I__1802 (
            .O(N__16786),
            .I(\ALU.madd_129 ));
    InMux I__1801 (
            .O(N__16781),
            .I(N__16778));
    LocalMux I__1800 (
            .O(N__16778),
            .I(\ALU.a5_b_4 ));
    CascadeMux I__1799 (
            .O(N__16775),
            .I(\ALU.a5_b_4_cascade_ ));
    CascadeMux I__1798 (
            .O(N__16772),
            .I(\ALU.madd_133_cascade_ ));
    InMux I__1797 (
            .O(N__16769),
            .I(N__16763));
    InMux I__1796 (
            .O(N__16768),
            .I(N__16763));
    LocalMux I__1795 (
            .O(N__16763),
            .I(N__16760));
    Span4Mux_v I__1794 (
            .O(N__16760),
            .I(N__16756));
    InMux I__1793 (
            .O(N__16759),
            .I(N__16753));
    Span4Mux_v I__1792 (
            .O(N__16756),
            .I(N__16750));
    LocalMux I__1791 (
            .O(N__16753),
            .I(N__16747));
    Odrv4 I__1790 (
            .O(N__16750),
            .I(\ALU.madd_237_0_tz_0 ));
    Odrv4 I__1789 (
            .O(N__16747),
            .I(\ALU.madd_237_0_tz_0 ));
    InMux I__1788 (
            .O(N__16742),
            .I(N__16736));
    InMux I__1787 (
            .O(N__16741),
            .I(N__16736));
    LocalMux I__1786 (
            .O(N__16736),
            .I(\ALU.madd_133 ));
    InMux I__1785 (
            .O(N__16733),
            .I(N__16729));
    CascadeMux I__1784 (
            .O(N__16732),
            .I(N__16726));
    LocalMux I__1783 (
            .O(N__16729),
            .I(N__16722));
    InMux I__1782 (
            .O(N__16726),
            .I(N__16717));
    InMux I__1781 (
            .O(N__16725),
            .I(N__16717));
    Sp12to4 I__1780 (
            .O(N__16722),
            .I(N__16712));
    LocalMux I__1779 (
            .O(N__16717),
            .I(N__16712));
    Span12Mux_v I__1778 (
            .O(N__16712),
            .I(N__16709));
    Odrv12 I__1777 (
            .O(N__16709),
            .I(\ALU.madd_138 ));
    CascadeMux I__1776 (
            .O(N__16706),
            .I(\ALU.madd_128_0_0_0_cascade_ ));
    InMux I__1775 (
            .O(N__16703),
            .I(N__16694));
    InMux I__1774 (
            .O(N__16702),
            .I(N__16694));
    InMux I__1773 (
            .O(N__16701),
            .I(N__16694));
    LocalMux I__1772 (
            .O(N__16694),
            .I(\ALU.madd_70 ));
    CascadeMux I__1771 (
            .O(N__16691),
            .I(\ALU.madd_237_0_tz_0_1_cascade_ ));
    InMux I__1770 (
            .O(N__16688),
            .I(N__16682));
    InMux I__1769 (
            .O(N__16687),
            .I(N__16679));
    InMux I__1768 (
            .O(N__16686),
            .I(N__16674));
    InMux I__1767 (
            .O(N__16685),
            .I(N__16674));
    LocalMux I__1766 (
            .O(N__16682),
            .I(N__16669));
    LocalMux I__1765 (
            .O(N__16679),
            .I(N__16669));
    LocalMux I__1764 (
            .O(N__16674),
            .I(N__16666));
    Span12Mux_v I__1763 (
            .O(N__16669),
            .I(N__16663));
    Odrv4 I__1762 (
            .O(N__16666),
            .I(\ALU.g0_0_0 ));
    Odrv12 I__1761 (
            .O(N__16663),
            .I(\ALU.g0_0_0 ));
    InMux I__1760 (
            .O(N__16658),
            .I(N__16655));
    LocalMux I__1759 (
            .O(N__16655),
            .I(N__16652));
    Sp12to4 I__1758 (
            .O(N__16652),
            .I(N__16649));
    Odrv12 I__1757 (
            .O(N__16649),
            .I(\ALU.N_1537_0_0_1 ));
    CascadeMux I__1756 (
            .O(N__16646),
            .I(\ALU.i6_mux_cascade_ ));
    CascadeMux I__1755 (
            .O(N__16643),
            .I(\ALU.un2_addsub_axb_7_cascade_ ));
    CascadeMux I__1754 (
            .O(N__16640),
            .I(\ALU.a0_b_8_cascade_ ));
    InMux I__1753 (
            .O(N__16637),
            .I(N__16633));
    InMux I__1752 (
            .O(N__16636),
            .I(N__16630));
    LocalMux I__1751 (
            .O(N__16633),
            .I(\ALU.madd_103 ));
    LocalMux I__1750 (
            .O(N__16630),
            .I(\ALU.madd_103 ));
    InMux I__1749 (
            .O(N__16625),
            .I(N__16622));
    LocalMux I__1748 (
            .O(N__16622),
            .I(\ALU.madd_124 ));
    InMux I__1747 (
            .O(N__16619),
            .I(N__16610));
    InMux I__1746 (
            .O(N__16618),
            .I(N__16610));
    InMux I__1745 (
            .O(N__16617),
            .I(N__16610));
    LocalMux I__1744 (
            .O(N__16610),
            .I(\ALU.madd_148 ));
    CascadeMux I__1743 (
            .O(N__16607),
            .I(\ALU.madd_148_cascade_ ));
    InMux I__1742 (
            .O(N__16604),
            .I(N__16598));
    InMux I__1741 (
            .O(N__16603),
            .I(N__16598));
    LocalMux I__1740 (
            .O(N__16598),
            .I(\ALU.madd_247_0_tz_0 ));
    CascadeMux I__1739 (
            .O(N__16595),
            .I(N__16592));
    InMux I__1738 (
            .O(N__16592),
            .I(N__16587));
    InMux I__1737 (
            .O(N__16591),
            .I(N__16584));
    InMux I__1736 (
            .O(N__16590),
            .I(N__16581));
    LocalMux I__1735 (
            .O(N__16587),
            .I(\ALU.madd_143 ));
    LocalMux I__1734 (
            .O(N__16584),
            .I(\ALU.madd_143 ));
    LocalMux I__1733 (
            .O(N__16581),
            .I(\ALU.madd_143 ));
    InMux I__1732 (
            .O(N__16574),
            .I(N__16567));
    InMux I__1731 (
            .O(N__16573),
            .I(N__16567));
    InMux I__1730 (
            .O(N__16572),
            .I(N__16564));
    LocalMux I__1729 (
            .O(N__16567),
            .I(\ALU.madd_181 ));
    LocalMux I__1728 (
            .O(N__16564),
            .I(\ALU.madd_181 ));
    CascadeMux I__1727 (
            .O(N__16559),
            .I(\ALU.madd_280_cascade_ ));
    InMux I__1726 (
            .O(N__16556),
            .I(N__16550));
    InMux I__1725 (
            .O(N__16555),
            .I(N__16550));
    LocalMux I__1724 (
            .O(N__16550),
            .I(N__16547));
    Odrv4 I__1723 (
            .O(N__16547),
            .I(\ALU.madd_285 ));
    InMux I__1722 (
            .O(N__16544),
            .I(N__16541));
    LocalMux I__1721 (
            .O(N__16541),
            .I(\ALU.madd_326 ));
    CascadeMux I__1720 (
            .O(N__16538),
            .I(N__16534));
    CascadeMux I__1719 (
            .O(N__16537),
            .I(N__16531));
    InMux I__1718 (
            .O(N__16534),
            .I(N__16526));
    InMux I__1717 (
            .O(N__16531),
            .I(N__16526));
    LocalMux I__1716 (
            .O(N__16526),
            .I(N__16523));
    Span4Mux_v I__1715 (
            .O(N__16523),
            .I(N__16520));
    Odrv4 I__1714 (
            .O(N__16520),
            .I(\ALU.a4_b_7 ));
    CascadeMux I__1713 (
            .O(N__16517),
            .I(\ALU.a4_b_7_cascade_ ));
    CascadeMux I__1712 (
            .O(N__16514),
            .I(\ALU.madd_233_cascade_ ));
    InMux I__1711 (
            .O(N__16511),
            .I(N__16507));
    InMux I__1710 (
            .O(N__16510),
            .I(N__16504));
    LocalMux I__1709 (
            .O(N__16507),
            .I(N__16499));
    LocalMux I__1708 (
            .O(N__16504),
            .I(N__16499));
    Odrv12 I__1707 (
            .O(N__16499),
            .I(\ALU.madd_237 ));
    InMux I__1706 (
            .O(N__16496),
            .I(N__16492));
    InMux I__1705 (
            .O(N__16495),
            .I(N__16489));
    LocalMux I__1704 (
            .O(N__16492),
            .I(\ALU.madd_242 ));
    LocalMux I__1703 (
            .O(N__16489),
            .I(\ALU.madd_242 ));
    CascadeMux I__1702 (
            .O(N__16484),
            .I(\ALU.madd_247_cascade_ ));
    InMux I__1701 (
            .O(N__16481),
            .I(N__16478));
    LocalMux I__1700 (
            .O(N__16478),
            .I(\ALU.madd_295_0 ));
    CascadeMux I__1699 (
            .O(N__16475),
            .I(N__16472));
    InMux I__1698 (
            .O(N__16472),
            .I(N__16469));
    LocalMux I__1697 (
            .O(N__16469),
            .I(\ALU.madd_N_10 ));
    InMux I__1696 (
            .O(N__16466),
            .I(N__16463));
    LocalMux I__1695 (
            .O(N__16463),
            .I(\ALU.madd_247 ));
    CascadeMux I__1694 (
            .O(N__16460),
            .I(\ALU.madd_N_10_cascade_ ));
    InMux I__1693 (
            .O(N__16457),
            .I(N__16454));
    LocalMux I__1692 (
            .O(N__16454),
            .I(\ALU.madd_N_5_0 ));
    InMux I__1691 (
            .O(N__16451),
            .I(N__16444));
    InMux I__1690 (
            .O(N__16450),
            .I(N__16444));
    CascadeMux I__1689 (
            .O(N__16449),
            .I(N__16441));
    LocalMux I__1688 (
            .O(N__16444),
            .I(N__16438));
    InMux I__1687 (
            .O(N__16441),
            .I(N__16435));
    Odrv4 I__1686 (
            .O(N__16438),
            .I(\ALU.madd_190 ));
    LocalMux I__1685 (
            .O(N__16435),
            .I(\ALU.madd_190 ));
    CascadeMux I__1684 (
            .O(N__16430),
            .I(N__16427));
    InMux I__1683 (
            .O(N__16427),
            .I(N__16421));
    InMux I__1682 (
            .O(N__16426),
            .I(N__16421));
    LocalMux I__1681 (
            .O(N__16421),
            .I(N__16418));
    Odrv4 I__1680 (
            .O(N__16418),
            .I(\ALU.madd_238_0 ));
    InMux I__1679 (
            .O(N__16415),
            .I(N__16412));
    LocalMux I__1678 (
            .O(N__16412),
            .I(\ALU.madd_233 ));
    InMux I__1677 (
            .O(N__16409),
            .I(N__16404));
    InMux I__1676 (
            .O(N__16408),
            .I(N__16399));
    InMux I__1675 (
            .O(N__16407),
            .I(N__16399));
    LocalMux I__1674 (
            .O(N__16404),
            .I(\ALU.madd_327 ));
    LocalMux I__1673 (
            .O(N__16399),
            .I(\ALU.madd_327 ));
    InMux I__1672 (
            .O(N__16394),
            .I(N__16388));
    InMux I__1671 (
            .O(N__16393),
            .I(N__16388));
    LocalMux I__1670 (
            .O(N__16388),
            .I(\ALU.madd_208 ));
    CascadeMux I__1669 (
            .O(N__16385),
            .I(\ALU.N_225_0_cascade_ ));
    CascadeMux I__1668 (
            .O(N__16382),
            .I(\ALU.madd_290_0_cascade_ ));
    CascadeMux I__1667 (
            .O(N__16379),
            .I(\ALU.madd_299_cascade_ ));
    InMux I__1666 (
            .O(N__16376),
            .I(N__16373));
    LocalMux I__1665 (
            .O(N__16373),
            .I(N__16370));
    Span4Mux_h I__1664 (
            .O(N__16370),
            .I(N__16365));
    InMux I__1663 (
            .O(N__16369),
            .I(N__16360));
    InMux I__1662 (
            .O(N__16368),
            .I(N__16360));
    Span4Mux_v I__1661 (
            .O(N__16365),
            .I(N__16357));
    LocalMux I__1660 (
            .O(N__16360),
            .I(N__16354));
    Odrv4 I__1659 (
            .O(N__16357),
            .I(\ALU.g0_11 ));
    Odrv4 I__1658 (
            .O(N__16354),
            .I(\ALU.g0_11 ));
    InMux I__1657 (
            .O(N__16349),
            .I(N__16346));
    LocalMux I__1656 (
            .O(N__16346),
            .I(N__16342));
    InMux I__1655 (
            .O(N__16345),
            .I(N__16339));
    Odrv12 I__1654 (
            .O(N__16342),
            .I(\ALU.madd_299 ));
    LocalMux I__1653 (
            .O(N__16339),
            .I(\ALU.madd_299 ));
    InMux I__1652 (
            .O(N__16334),
            .I(N__16331));
    LocalMux I__1651 (
            .O(N__16331),
            .I(N__16328));
    Odrv4 I__1650 (
            .O(N__16328),
            .I(\ALU.madd_223_0 ));
    InMux I__1649 (
            .O(N__16325),
            .I(N__16321));
    InMux I__1648 (
            .O(N__16324),
            .I(N__16318));
    LocalMux I__1647 (
            .O(N__16321),
            .I(\ALU.madd_228 ));
    LocalMux I__1646 (
            .O(N__16318),
            .I(\ALU.madd_228 ));
    InMux I__1645 (
            .O(N__16313),
            .I(N__16309));
    CascadeMux I__1644 (
            .O(N__16312),
            .I(N__16304));
    LocalMux I__1643 (
            .O(N__16309),
            .I(N__16301));
    InMux I__1642 (
            .O(N__16308),
            .I(N__16296));
    InMux I__1641 (
            .O(N__16307),
            .I(N__16296));
    InMux I__1640 (
            .O(N__16304),
            .I(N__16293));
    Odrv4 I__1639 (
            .O(N__16301),
            .I(\ALU.madd_170 ));
    LocalMux I__1638 (
            .O(N__16296),
            .I(\ALU.madd_170 ));
    LocalMux I__1637 (
            .O(N__16293),
            .I(\ALU.madd_170 ));
    CascadeMux I__1636 (
            .O(N__16286),
            .I(\ALU.madd_265_0_cascade_ ));
    InMux I__1635 (
            .O(N__16283),
            .I(N__16280));
    LocalMux I__1634 (
            .O(N__16280),
            .I(N__16275));
    InMux I__1633 (
            .O(N__16279),
            .I(N__16272));
    InMux I__1632 (
            .O(N__16278),
            .I(N__16269));
    Odrv12 I__1631 (
            .O(N__16275),
            .I(\ALU.madd_280 ));
    LocalMux I__1630 (
            .O(N__16272),
            .I(\ALU.madd_280 ));
    LocalMux I__1629 (
            .O(N__16269),
            .I(\ALU.madd_280 ));
    CascadeMux I__1628 (
            .O(N__16262),
            .I(\ALU.madd_223_0_cascade_ ));
    InMux I__1627 (
            .O(N__16259),
            .I(N__16256));
    LocalMux I__1626 (
            .O(N__16256),
            .I(\ALU.N_1533_0 ));
    InMux I__1625 (
            .O(N__16253),
            .I(N__16250));
    LocalMux I__1624 (
            .O(N__16250),
            .I(N__16247));
    Span4Mux_s2_h I__1623 (
            .O(N__16247),
            .I(N__16244));
    Odrv4 I__1622 (
            .O(N__16244),
            .I(\ALU.N_1559_0 ));
    InMux I__1621 (
            .O(N__16241),
            .I(N__16235));
    InMux I__1620 (
            .O(N__16240),
            .I(N__16235));
    LocalMux I__1619 (
            .O(N__16235),
            .I(\ALU.madd_165_0_tz ));
    InMux I__1618 (
            .O(N__16232),
            .I(N__16228));
    InMux I__1617 (
            .O(N__16231),
            .I(N__16225));
    LocalMux I__1616 (
            .O(N__16228),
            .I(\ALU.madd_165_0 ));
    LocalMux I__1615 (
            .O(N__16225),
            .I(\ALU.madd_165_0 ));
    CascadeMux I__1614 (
            .O(N__16220),
            .I(N__16217));
    InMux I__1613 (
            .O(N__16217),
            .I(N__16214));
    LocalMux I__1612 (
            .O(N__16214),
            .I(\ALU.a5_b_5 ));
    CascadeMux I__1611 (
            .O(N__16211),
            .I(\ALU.a5_b_5_cascade_ ));
    InMux I__1610 (
            .O(N__16208),
            .I(N__16204));
    InMux I__1609 (
            .O(N__16207),
            .I(N__16201));
    LocalMux I__1608 (
            .O(N__16204),
            .I(N__16196));
    LocalMux I__1607 (
            .O(N__16201),
            .I(N__16196));
    Odrv4 I__1606 (
            .O(N__16196),
            .I(\ALU.a4_b_6 ));
    CascadeMux I__1605 (
            .O(N__16193),
            .I(\ALU.madd_175_cascade_ ));
    CascadeMux I__1604 (
            .O(N__16190),
            .I(N__16186));
    CascadeMux I__1603 (
            .O(N__16189),
            .I(N__16182));
    InMux I__1602 (
            .O(N__16186),
            .I(N__16178));
    InMux I__1601 (
            .O(N__16185),
            .I(N__16171));
    InMux I__1600 (
            .O(N__16182),
            .I(N__16171));
    InMux I__1599 (
            .O(N__16181),
            .I(N__16171));
    LocalMux I__1598 (
            .O(N__16178),
            .I(N__16166));
    LocalMux I__1597 (
            .O(N__16171),
            .I(N__16166));
    Odrv4 I__1596 (
            .O(N__16166),
            .I(\ALU.madd_232 ));
    InMux I__1595 (
            .O(N__16163),
            .I(N__16160));
    LocalMux I__1594 (
            .O(N__16160),
            .I(\ALU.madd_175 ));
    InMux I__1593 (
            .O(N__16157),
            .I(N__16151));
    InMux I__1592 (
            .O(N__16156),
            .I(N__16151));
    LocalMux I__1591 (
            .O(N__16151),
            .I(\ALU.madd_213_0 ));
    CascadeMux I__1590 (
            .O(N__16148),
            .I(\ALU.a7_b_4_cascade_ ));
    InMux I__1589 (
            .O(N__16145),
            .I(N__16142));
    LocalMux I__1588 (
            .O(N__16142),
            .I(\ALU.madd_i1_mux_2 ));
    InMux I__1587 (
            .O(N__16139),
            .I(N__16135));
    CascadeMux I__1586 (
            .O(N__16138),
            .I(N__16132));
    LocalMux I__1585 (
            .O(N__16135),
            .I(N__16129));
    InMux I__1584 (
            .O(N__16132),
            .I(N__16126));
    Odrv4 I__1583 (
            .O(N__16129),
            .I(\ALU.madd_289 ));
    LocalMux I__1582 (
            .O(N__16126),
            .I(\ALU.madd_289 ));
    InMux I__1581 (
            .O(N__16121),
            .I(N__16115));
    InMux I__1580 (
            .O(N__16120),
            .I(N__16115));
    LocalMux I__1579 (
            .O(N__16115),
            .I(\ALU.madd_227 ));
    CascadeMux I__1578 (
            .O(N__16112),
            .I(\ALU.madd_227_cascade_ ));
    CascadeMux I__1577 (
            .O(N__16109),
            .I(\ALU.madd_165_0_0_cascade_ ));
    CascadeMux I__1576 (
            .O(N__16106),
            .I(\ALU.madd_170_0_tz_cascade_ ));
    InMux I__1575 (
            .O(N__16103),
            .I(N__16098));
    InMux I__1574 (
            .O(N__16102),
            .I(N__16093));
    InMux I__1573 (
            .O(N__16101),
            .I(N__16093));
    LocalMux I__1572 (
            .O(N__16098),
            .I(N__16090));
    LocalMux I__1571 (
            .O(N__16093),
            .I(\ALU.madd_90 ));
    Odrv4 I__1570 (
            .O(N__16090),
            .I(\ALU.madd_90 ));
    InMux I__1569 (
            .O(N__16085),
            .I(N__16082));
    LocalMux I__1568 (
            .O(N__16082),
            .I(\ALU.madd_340_0 ));
    CascadeMux I__1567 (
            .O(N__16079),
            .I(\ALU.g0_1_cascade_ ));
    InMux I__1566 (
            .O(N__16076),
            .I(N__16073));
    LocalMux I__1565 (
            .O(N__16073),
            .I(\ALU.g2 ));
    InMux I__1564 (
            .O(N__16070),
            .I(N__16067));
    LocalMux I__1563 (
            .O(N__16067),
            .I(\ALU.N_1545_1 ));
    CascadeMux I__1562 (
            .O(N__16064),
            .I(\ALU.g0_3_cascade_ ));
    InMux I__1561 (
            .O(N__16061),
            .I(N__16058));
    LocalMux I__1560 (
            .O(N__16058),
            .I(\ALU.madd_350_0 ));
    CascadeMux I__1559 (
            .O(N__16055),
            .I(\ALU.madd_350_0_cascade_ ));
    InMux I__1558 (
            .O(N__16052),
            .I(N__16044));
    InMux I__1557 (
            .O(N__16051),
            .I(N__16044));
    InMux I__1556 (
            .O(N__16050),
            .I(N__16041));
    InMux I__1555 (
            .O(N__16049),
            .I(N__16038));
    LocalMux I__1554 (
            .O(N__16044),
            .I(\ALU.madd_335 ));
    LocalMux I__1553 (
            .O(N__16041),
            .I(\ALU.madd_335 ));
    LocalMux I__1552 (
            .O(N__16038),
            .I(\ALU.madd_335 ));
    CascadeMux I__1551 (
            .O(N__16031),
            .I(\ALU.a4_b_8_cascade_ ));
    InMux I__1550 (
            .O(N__16028),
            .I(N__16022));
    InMux I__1549 (
            .O(N__16027),
            .I(N__16022));
    LocalMux I__1548 (
            .O(N__16022),
            .I(\ALU.madd_269 ));
    CascadeMux I__1547 (
            .O(N__16019),
            .I(\ALU.madd_i1_mux_cascade_ ));
    InMux I__1546 (
            .O(N__16016),
            .I(N__16013));
    LocalMux I__1545 (
            .O(N__16013),
            .I(N__16009));
    InMux I__1544 (
            .O(N__16012),
            .I(N__16006));
    Span4Mux_v I__1543 (
            .O(N__16009),
            .I(N__16003));
    LocalMux I__1542 (
            .O(N__16006),
            .I(N__16000));
    Odrv4 I__1541 (
            .O(N__16003),
            .I(\ALU.g0_14 ));
    Odrv4 I__1540 (
            .O(N__16000),
            .I(\ALU.g0_14 ));
    CascadeMux I__1539 (
            .O(N__15995),
            .I(\ALU.madd_i3_mux_cascade_ ));
    CascadeMux I__1538 (
            .O(N__15992),
            .I(\ALU.madd_331_cascade_ ));
    CascadeMux I__1537 (
            .O(N__15989),
            .I(N__15985));
    InMux I__1536 (
            .O(N__15988),
            .I(N__15980));
    InMux I__1535 (
            .O(N__15985),
            .I(N__15980));
    LocalMux I__1534 (
            .O(N__15980),
            .I(\ALU.madd_328 ));
    CascadeMux I__1533 (
            .O(N__15977),
            .I(\ALU.N_275_0_cascade_ ));
    InMux I__1532 (
            .O(N__15974),
            .I(N__15971));
    LocalMux I__1531 (
            .O(N__15971),
            .I(\ALU.g0_0_0_N_3L3 ));
    CascadeMux I__1530 (
            .O(N__15968),
            .I(\ALU.g0_0_0_N_4L5_cascade_ ));
    InMux I__1529 (
            .O(N__15965),
            .I(N__15962));
    LocalMux I__1528 (
            .O(N__15962),
            .I(\ALU.g0_0_0_N_3L3_0 ));
    CascadeMux I__1527 (
            .O(N__15959),
            .I(\ALU.a5_b_9_cascade_ ));
    CascadeMux I__1526 (
            .O(N__15956),
            .I(\ALU.operand2_8_cascade_ ));
    CascadeMux I__1525 (
            .O(N__15953),
            .I(N__15950));
    InMux I__1524 (
            .O(N__15950),
            .I(N__15947));
    LocalMux I__1523 (
            .O(N__15947),
            .I(N__15944));
    Span4Mux_v I__1522 (
            .O(N__15944),
            .I(N__15941));
    Span4Mux_v I__1521 (
            .O(N__15941),
            .I(N__15938));
    Odrv4 I__1520 (
            .O(N__15938),
            .I(\ALU.a1_b_8 ));
    CascadeMux I__1519 (
            .O(N__15935),
            .I(\ALU.a1_b_8_cascade_ ));
    CascadeMux I__1518 (
            .O(N__15932),
            .I(N_661_0_cascade_));
    CascadeMux I__1517 (
            .O(N__15929),
            .I(\ALU.un2_addsub_axb_8_cascade_ ));
    CascadeMux I__1516 (
            .O(N__15926),
            .I(N__15922));
    InMux I__1515 (
            .O(N__15925),
            .I(N__15916));
    InMux I__1514 (
            .O(N__15922),
            .I(N__15916));
    CascadeMux I__1513 (
            .O(N__15921),
            .I(N__15913));
    LocalMux I__1512 (
            .O(N__15916),
            .I(N__15910));
    InMux I__1511 (
            .O(N__15913),
            .I(N__15907));
    Odrv4 I__1510 (
            .O(N__15910),
            .I(RXbuffer_0));
    LocalMux I__1509 (
            .O(N__15907),
            .I(RXbuffer_0));
    CascadeMux I__1508 (
            .O(N__15902),
            .I(N__15898));
    CascadeMux I__1507 (
            .O(N__15901),
            .I(N__15893));
    InMux I__1506 (
            .O(N__15898),
            .I(N__15887));
    InMux I__1505 (
            .O(N__15897),
            .I(N__15887));
    InMux I__1504 (
            .O(N__15896),
            .I(N__15884));
    InMux I__1503 (
            .O(N__15893),
            .I(N__15881));
    InMux I__1502 (
            .O(N__15892),
            .I(N__15878));
    LocalMux I__1501 (
            .O(N__15887),
            .I(N__15875));
    LocalMux I__1500 (
            .O(N__15884),
            .I(N__15870));
    LocalMux I__1499 (
            .O(N__15881),
            .I(N__15870));
    LocalMux I__1498 (
            .O(N__15878),
            .I(RXbuffer_7));
    Odrv4 I__1497 (
            .O(N__15875),
            .I(RXbuffer_7));
    Odrv4 I__1496 (
            .O(N__15870),
            .I(RXbuffer_7));
    CascadeMux I__1495 (
            .O(N__15863),
            .I(N__15858));
    CascadeMux I__1494 (
            .O(N__15862),
            .I(N__15854));
    CascadeMux I__1493 (
            .O(N__15861),
            .I(N__15851));
    InMux I__1492 (
            .O(N__15858),
            .I(N__15847));
    InMux I__1491 (
            .O(N__15857),
            .I(N__15842));
    InMux I__1490 (
            .O(N__15854),
            .I(N__15842));
    InMux I__1489 (
            .O(N__15851),
            .I(N__15839));
    InMux I__1488 (
            .O(N__15850),
            .I(N__15836));
    LocalMux I__1487 (
            .O(N__15847),
            .I(N__15833));
    LocalMux I__1486 (
            .O(N__15842),
            .I(N__15830));
    LocalMux I__1485 (
            .O(N__15839),
            .I(N__15827));
    LocalMux I__1484 (
            .O(N__15836),
            .I(RXbuffer_1));
    Odrv4 I__1483 (
            .O(N__15833),
            .I(RXbuffer_1));
    Odrv4 I__1482 (
            .O(N__15830),
            .I(RXbuffer_1));
    Odrv4 I__1481 (
            .O(N__15827),
            .I(RXbuffer_1));
    CascadeMux I__1480 (
            .O(N__15818),
            .I(N__15815));
    InMux I__1479 (
            .O(N__15815),
            .I(N__15806));
    InMux I__1478 (
            .O(N__15814),
            .I(N__15806));
    InMux I__1477 (
            .O(N__15813),
            .I(N__15803));
    InMux I__1476 (
            .O(N__15812),
            .I(N__15798));
    InMux I__1475 (
            .O(N__15811),
            .I(N__15798));
    LocalMux I__1474 (
            .O(N__15806),
            .I(N__15795));
    LocalMux I__1473 (
            .O(N__15803),
            .I(N__15788));
    LocalMux I__1472 (
            .O(N__15798),
            .I(N__15788));
    Span4Mux_v I__1471 (
            .O(N__15795),
            .I(N__15788));
    Span4Mux_v I__1470 (
            .O(N__15788),
            .I(N__15785));
    Odrv4 I__1469 (
            .O(N__15785),
            .I(RXbuffer_3));
    InMux I__1468 (
            .O(N__15782),
            .I(N__15779));
    LocalMux I__1467 (
            .O(N__15779),
            .I(N__15776));
    Span4Mux_s0_v I__1466 (
            .O(N__15776),
            .I(N__15772));
    CascadeMux I__1465 (
            .O(N__15775),
            .I(N__15769));
    Span4Mux_v I__1464 (
            .O(N__15772),
            .I(N__15766));
    InMux I__1463 (
            .O(N__15769),
            .I(N__15763));
    Odrv4 I__1462 (
            .O(N__15766),
            .I(testWordZ0Z_13));
    LocalMux I__1461 (
            .O(N__15763),
            .I(testWordZ0Z_13));
    CascadeMux I__1460 (
            .O(N__15758),
            .I(\ALU.m304_nsZ0Z_1_cascade_ ));
    CascadeMux I__1459 (
            .O(N__15755),
            .I(\ALU.i73_mux_1_cascade_ ));
    InMux I__1458 (
            .O(N__15752),
            .I(N__15749));
    LocalMux I__1457 (
            .O(N__15749),
            .I(clkdivZ0Z_16));
    InMux I__1456 (
            .O(N__15746),
            .I(bfn_1_18_0_));
    InMux I__1455 (
            .O(N__15743),
            .I(N__15740));
    LocalMux I__1454 (
            .O(N__15740),
            .I(clkdivZ0Z_17));
    InMux I__1453 (
            .O(N__15737),
            .I(clkdiv_cry_16));
    InMux I__1452 (
            .O(N__15734),
            .I(N__15731));
    LocalMux I__1451 (
            .O(N__15731),
            .I(clkdivZ0Z_18));
    InMux I__1450 (
            .O(N__15728),
            .I(clkdiv_cry_17));
    InMux I__1449 (
            .O(N__15725),
            .I(N__15722));
    LocalMux I__1448 (
            .O(N__15722),
            .I(clkdivZ0Z_19));
    InMux I__1447 (
            .O(N__15719),
            .I(clkdiv_cry_18));
    InMux I__1446 (
            .O(N__15716),
            .I(N__15713));
    LocalMux I__1445 (
            .O(N__15713),
            .I(clkdivZ0Z_20));
    InMux I__1444 (
            .O(N__15710),
            .I(clkdiv_cry_19));
    InMux I__1443 (
            .O(N__15707),
            .I(N__15704));
    LocalMux I__1442 (
            .O(N__15704),
            .I(clkdivZ0Z_21));
    InMux I__1441 (
            .O(N__15701),
            .I(clkdiv_cry_20));
    InMux I__1440 (
            .O(N__15698),
            .I(N__15695));
    LocalMux I__1439 (
            .O(N__15695),
            .I(clkdivZ0Z_22));
    InMux I__1438 (
            .O(N__15692),
            .I(clkdiv_cry_21));
    InMux I__1437 (
            .O(N__15689),
            .I(clkdiv_cry_22));
    IoInMux I__1436 (
            .O(N__15686),
            .I(N__15683));
    LocalMux I__1435 (
            .O(N__15683),
            .I(N__15680));
    Span12Mux_s7_v I__1434 (
            .O(N__15680),
            .I(N__15676));
    InMux I__1433 (
            .O(N__15679),
            .I(N__15673));
    Odrv12 I__1432 (
            .O(N__15676),
            .I(GPIO3_c));
    LocalMux I__1431 (
            .O(N__15673),
            .I(GPIO3_c));
    InMux I__1430 (
            .O(N__15668),
            .I(N__15665));
    LocalMux I__1429 (
            .O(N__15665),
            .I(clkdivZ0Z_7));
    InMux I__1428 (
            .O(N__15662),
            .I(clkdiv_cry_6));
    InMux I__1427 (
            .O(N__15659),
            .I(N__15656));
    LocalMux I__1426 (
            .O(N__15656),
            .I(clkdivZ0Z_8));
    InMux I__1425 (
            .O(N__15653),
            .I(bfn_1_17_0_));
    InMux I__1424 (
            .O(N__15650),
            .I(N__15647));
    LocalMux I__1423 (
            .O(N__15647),
            .I(clkdivZ0Z_9));
    InMux I__1422 (
            .O(N__15644),
            .I(clkdiv_cry_8));
    InMux I__1421 (
            .O(N__15641),
            .I(N__15638));
    LocalMux I__1420 (
            .O(N__15638),
            .I(clkdivZ0Z_10));
    InMux I__1419 (
            .O(N__15635),
            .I(clkdiv_cry_9));
    InMux I__1418 (
            .O(N__15632),
            .I(N__15629));
    LocalMux I__1417 (
            .O(N__15629),
            .I(clkdivZ0Z_11));
    InMux I__1416 (
            .O(N__15626),
            .I(clkdiv_cry_10));
    InMux I__1415 (
            .O(N__15623),
            .I(N__15620));
    LocalMux I__1414 (
            .O(N__15620),
            .I(clkdivZ0Z_12));
    InMux I__1413 (
            .O(N__15617),
            .I(clkdiv_cry_11));
    InMux I__1412 (
            .O(N__15614),
            .I(N__15611));
    LocalMux I__1411 (
            .O(N__15611),
            .I(clkdivZ0Z_13));
    InMux I__1410 (
            .O(N__15608),
            .I(clkdiv_cry_12));
    InMux I__1409 (
            .O(N__15605),
            .I(N__15602));
    LocalMux I__1408 (
            .O(N__15602),
            .I(clkdivZ0Z_14));
    InMux I__1407 (
            .O(N__15599),
            .I(clkdiv_cry_13));
    InMux I__1406 (
            .O(N__15596),
            .I(N__15593));
    LocalMux I__1405 (
            .O(N__15593),
            .I(clkdivZ0Z_15));
    InMux I__1404 (
            .O(N__15590),
            .I(clkdiv_cry_14));
    InMux I__1403 (
            .O(N__15587),
            .I(N__15583));
    InMux I__1402 (
            .O(N__15586),
            .I(N__15580));
    LocalMux I__1401 (
            .O(N__15583),
            .I(\ALU.madd_324 ));
    LocalMux I__1400 (
            .O(N__15580),
            .I(\ALU.madd_324 ));
    CascadeMux I__1399 (
            .O(N__15575),
            .I(\ALU.madd_326_cascade_ ));
    InMux I__1398 (
            .O(N__15572),
            .I(N__15567));
    InMux I__1397 (
            .O(N__15571),
            .I(N__15562));
    InMux I__1396 (
            .O(N__15570),
            .I(N__15562));
    LocalMux I__1395 (
            .O(N__15567),
            .I(\ALU.madd_325 ));
    LocalMux I__1394 (
            .O(N__15562),
            .I(\ALU.madd_325 ));
    InMux I__1393 (
            .O(N__15557),
            .I(N__15554));
    LocalMux I__1392 (
            .O(N__15554),
            .I(clkdivZ0Z_0));
    InMux I__1391 (
            .O(N__15551),
            .I(bfn_1_16_0_));
    InMux I__1390 (
            .O(N__15548),
            .I(N__15545));
    LocalMux I__1389 (
            .O(N__15545),
            .I(clkdivZ0Z_1));
    InMux I__1388 (
            .O(N__15542),
            .I(clkdiv_cry_0));
    InMux I__1387 (
            .O(N__15539),
            .I(N__15536));
    LocalMux I__1386 (
            .O(N__15536),
            .I(clkdivZ0Z_2));
    InMux I__1385 (
            .O(N__15533),
            .I(clkdiv_cry_1));
    InMux I__1384 (
            .O(N__15530),
            .I(N__15527));
    LocalMux I__1383 (
            .O(N__15527),
            .I(clkdivZ0Z_3));
    InMux I__1382 (
            .O(N__15524),
            .I(clkdiv_cry_2));
    InMux I__1381 (
            .O(N__15521),
            .I(N__15518));
    LocalMux I__1380 (
            .O(N__15518),
            .I(clkdivZ0Z_4));
    InMux I__1379 (
            .O(N__15515),
            .I(clkdiv_cry_3));
    InMux I__1378 (
            .O(N__15512),
            .I(N__15509));
    LocalMux I__1377 (
            .O(N__15509),
            .I(clkdivZ0Z_5));
    InMux I__1376 (
            .O(N__15506),
            .I(clkdiv_cry_4));
    InMux I__1375 (
            .O(N__15503),
            .I(N__15500));
    LocalMux I__1374 (
            .O(N__15500),
            .I(clkdivZ0Z_6));
    InMux I__1373 (
            .O(N__15497),
            .I(clkdiv_cry_5));
    CascadeMux I__1372 (
            .O(N__15494),
            .I(\ALU.madd_144_cascade_ ));
    CascadeMux I__1371 (
            .O(N__15491),
            .I(\ALU.madd_324_cascade_ ));
    CascadeMux I__1370 (
            .O(N__15488),
            .I(\ALU.madd_N_9_cascade_ ));
    InMux I__1369 (
            .O(N__15485),
            .I(N__15482));
    LocalMux I__1368 (
            .O(N__15482),
            .I(\ALU.madd_191_0 ));
    CascadeMux I__1367 (
            .O(N__15479),
            .I(N__15473));
    InMux I__1366 (
            .O(N__15478),
            .I(N__15468));
    InMux I__1365 (
            .O(N__15477),
            .I(N__15468));
    InMux I__1364 (
            .O(N__15476),
            .I(N__15463));
    InMux I__1363 (
            .O(N__15473),
            .I(N__15463));
    LocalMux I__1362 (
            .O(N__15468),
            .I(N__15460));
    LocalMux I__1361 (
            .O(N__15463),
            .I(N__15455));
    Span4Mux_s1_h I__1360 (
            .O(N__15460),
            .I(N__15455));
    Odrv4 I__1359 (
            .O(N__15455),
            .I(\ALU.madd_186 ));
    CascadeMux I__1358 (
            .O(N__15452),
            .I(\ALU.madd_191_0_cascade_ ));
    CascadeMux I__1357 (
            .O(N__15449),
            .I(\ALU.a8_b_3_cascade_ ));
    InMux I__1356 (
            .O(N__15446),
            .I(N__15441));
    InMux I__1355 (
            .O(N__15445),
            .I(N__15438));
    InMux I__1354 (
            .O(N__15444),
            .I(N__15435));
    LocalMux I__1353 (
            .O(N__15441),
            .I(\ALU.a8_b_3 ));
    LocalMux I__1352 (
            .O(N__15438),
            .I(\ALU.a8_b_3 ));
    LocalMux I__1351 (
            .O(N__15435),
            .I(\ALU.a8_b_3 ));
    InMux I__1350 (
            .O(N__15428),
            .I(N__15425));
    LocalMux I__1349 (
            .O(N__15425),
            .I(N__15422));
    Odrv12 I__1348 (
            .O(N__15422),
            .I(\ALU.g0_0_2 ));
    CascadeMux I__1347 (
            .O(N__15419),
            .I(\ALU.g0_0_cascade_ ));
    InMux I__1346 (
            .O(N__15416),
            .I(N__15413));
    LocalMux I__1345 (
            .O(N__15413),
            .I(\ALU.N_1527_1_0 ));
    CascadeMux I__1344 (
            .O(N__15410),
            .I(N__15407));
    InMux I__1343 (
            .O(N__15407),
            .I(N__15404));
    LocalMux I__1342 (
            .O(N__15404),
            .I(N__15401));
    Span4Mux_v I__1341 (
            .O(N__15401),
            .I(N__15398));
    Odrv4 I__1340 (
            .O(N__15398),
            .I(\ALU.g2_0_1 ));
    InMux I__1339 (
            .O(N__15395),
            .I(N__15392));
    LocalMux I__1338 (
            .O(N__15392),
            .I(\ALU.g1 ));
    InMux I__1337 (
            .O(N__15389),
            .I(N__15386));
    LocalMux I__1336 (
            .O(N__15386),
            .I(N__15383));
    Odrv4 I__1335 (
            .O(N__15383),
            .I(\ALU.g0_1_0 ));
    CascadeMux I__1334 (
            .O(N__15380),
            .I(\ALU.madd_124_0_cascade_ ));
    CascadeMux I__1333 (
            .O(N__15377),
            .I(\ALU.madd_124_cascade_ ));
    CascadeMux I__1332 (
            .O(N__15374),
            .I(\ALU.madd_171_cascade_ ));
    CascadeMux I__1331 (
            .O(N__15371),
            .I(\ALU.madd_161_0_cascade_ ));
    InMux I__1330 (
            .O(N__15368),
            .I(N__15365));
    LocalMux I__1329 (
            .O(N__15365),
            .I(\ALU.madd_161 ));
    InMux I__1328 (
            .O(N__15362),
            .I(N__15356));
    InMux I__1327 (
            .O(N__15361),
            .I(N__15356));
    LocalMux I__1326 (
            .O(N__15356),
            .I(N__15353));
    Odrv4 I__1325 (
            .O(N__15353),
            .I(\ALU.madd_166 ));
    InMux I__1324 (
            .O(N__15350),
            .I(N__15347));
    LocalMux I__1323 (
            .O(N__15347),
            .I(\ALU.madd_171 ));
    CascadeMux I__1322 (
            .O(N__15344),
            .I(\ALU.madd_161_cascade_ ));
    CascadeMux I__1321 (
            .O(N__15341),
            .I(\ALU.N_217_0_cascade_ ));
    CascadeMux I__1320 (
            .O(N__15338),
            .I(\ALU.un9_addsub_axb_10_cascade_ ));
    CascadeMux I__1319 (
            .O(N__15335),
            .I(\ALU.a3_b_0_10_cascade_ ));
    CascadeMux I__1318 (
            .O(N__15332),
            .I(\ALU.g0_2_cascade_ ));
    InMux I__1317 (
            .O(N__15329),
            .I(N__15326));
    LocalMux I__1316 (
            .O(N__15326),
            .I(\ALU.N_1555_0 ));
    InMux I__1315 (
            .O(N__15323),
            .I(N__15320));
    LocalMux I__1314 (
            .O(N__15320),
            .I(\ALU.N_1527_0 ));
    CascadeMux I__1313 (
            .O(N__15317),
            .I(\ALU.madd_254_0_tz_cascade_ ));
    InMux I__1312 (
            .O(N__15314),
            .I(N__15311));
    LocalMux I__1311 (
            .O(N__15311),
            .I(\ALU.madd_141 ));
    CascadeMux I__1310 (
            .O(N__15308),
            .I(\ALU.madd_254_cascade_ ));
    InMux I__1309 (
            .O(N__15305),
            .I(N__15301));
    InMux I__1308 (
            .O(N__15304),
            .I(N__15298));
    LocalMux I__1307 (
            .O(N__15301),
            .I(\ALU.madd_254_0_tz ));
    LocalMux I__1306 (
            .O(N__15298),
            .I(\ALU.madd_254_0_tz ));
    CascadeMux I__1305 (
            .O(N__15293),
            .I(N__15290));
    InMux I__1304 (
            .O(N__15290),
            .I(N__15287));
    LocalMux I__1303 (
            .O(N__15287),
            .I(\ALU.m292_nsZ0Z_1 ));
    CascadeMux I__1302 (
            .O(N__15284),
            .I(\ALU.N_90_0_cascade_ ));
    CascadeMux I__1301 (
            .O(N__15281),
            .I(N__15277));
    InMux I__1300 (
            .O(N__15280),
            .I(N__15272));
    InMux I__1299 (
            .O(N__15277),
            .I(N__15272));
    LocalMux I__1298 (
            .O(N__15272),
            .I(ctrlOut_6));
    CascadeMux I__1297 (
            .O(N__15269),
            .I(\ALU.madd_315_0_cascade_ ));
    InMux I__1296 (
            .O(N__15266),
            .I(N__15263));
    LocalMux I__1295 (
            .O(N__15263),
            .I(\ALU.a12_b_1 ));
    InMux I__1294 (
            .O(N__15260),
            .I(N__15257));
    LocalMux I__1293 (
            .O(N__15257),
            .I(\ALU.madd_315_0 ));
    CascadeMux I__1292 (
            .O(N__15254),
            .I(\ALU.a12_b_1_cascade_ ));
    InMux I__1291 (
            .O(N__15251),
            .I(N__15245));
    InMux I__1290 (
            .O(N__15250),
            .I(N__15245));
    LocalMux I__1289 (
            .O(N__15245),
            .I(\ALU.madd_264 ));
    CascadeMux I__1288 (
            .O(N__15242),
            .I(\ALU.madd_141_0_cascade_ ));
    InMux I__1287 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__1286 (
            .O(N__15236),
            .I(\ALU.N_1545_0 ));
    InMux I__1285 (
            .O(N__15233),
            .I(N__15230));
    LocalMux I__1284 (
            .O(N__15230),
            .I(\ALU.madd_166_0 ));
    InMux I__1283 (
            .O(N__15227),
            .I(N__15215));
    InMux I__1282 (
            .O(N__15226),
            .I(N__15215));
    InMux I__1281 (
            .O(N__15225),
            .I(N__15215));
    InMux I__1280 (
            .O(N__15224),
            .I(N__15215));
    LocalMux I__1279 (
            .O(N__15215),
            .I(ctrlOut_5));
    CascadeMux I__1278 (
            .O(N__15212),
            .I(\ALU.N_223_0_cascade_ ));
    CascadeMux I__1277 (
            .O(N__15209),
            .I(\ALU.a9_b_3_cascade_ ));
    InMux I__1276 (
            .O(N__15206),
            .I(N__15200));
    InMux I__1275 (
            .O(N__15205),
            .I(N__15200));
    LocalMux I__1274 (
            .O(N__15200),
            .I(\ALU.a7_b_5 ));
    CascadeMux I__1273 (
            .O(N__15197),
            .I(N__15194));
    InMux I__1272 (
            .O(N__15194),
            .I(N__15191));
    LocalMux I__1271 (
            .O(N__15191),
            .I(\ALU.a9_b_3 ));
    CascadeMux I__1270 (
            .O(N__15188),
            .I(\ALU.g0_0_a3_2_0_cascade_ ));
    CascadeMux I__1269 (
            .O(N__15185),
            .I(N__15181));
    InMux I__1268 (
            .O(N__15184),
            .I(N__15176));
    InMux I__1267 (
            .O(N__15181),
            .I(N__15176));
    LocalMux I__1266 (
            .O(N__15176),
            .I(ctrlOut_8));
    CascadeMux I__1265 (
            .O(N__15173),
            .I(\ALU.m289_nsZ0Z_1_cascade_ ));
    INV \INVFTDI.TXshift_1C  (
            .O(\INVFTDI.TXshift_1C_net ),
            .I(N__47602));
    INV \INVFTDI.TXshift_0C  (
            .O(\INVFTDI.TXshift_0C_net ),
            .I(N__47607));
    INV \INVFTDI.baudAcc_1C  (
            .O(\INVFTDI.baudAcc_1C_net ),
            .I(N__47604));
    INV \INVFTDI.TXstate_0C  (
            .O(\INVFTDI.TXstate_0C_net ),
            .I(N__47601));
    INV \INVFTDI.gap_2C  (
            .O(\INVFTDI.gap_2C_net ),
            .I(N__47599));
    INV \INVFTDI.baudAcc_0C  (
            .O(\INVFTDI.baudAcc_0C_net ),
            .I(N__47603));
    INV \INVFTDI.gap_0C  (
            .O(\INVFTDI.gap_0C_net ),
            .I(N__47609));
    INV \INVFTDI.RXreadyC  (
            .O(\INVFTDI.RXreadyC_net ),
            .I(N__47617));
    INV \INVFTDI.RXbuffer_0C  (
            .O(\INVFTDI.RXbuffer_0C_net ),
            .I(N__47667));
    INV \INVFTDI.RXbuffer_3C  (
            .O(\INVFTDI.RXbuffer_3C_net ),
            .I(N__47654));
    defparam IN_MUX_bfv_13_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_2_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\ALU.madd_cry_7 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(clkdiv_cry_7),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(clkdiv_cry_15),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\ALU.un9_addsub_cry_7 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(\ALU.un2_addsub_cry_7 ),
            .carryinitout(bfn_6_10_0_));
    ICE_GB testState_RNIB7C_0_2 (
            .USERSIGNALTOGLOBALBUFFER(N__30743),
            .GLOBALBUFFEROUTPUT(testState_i_g_2));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \FTDI.RXbuffer_3_LC_1_2_4 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_3_LC_1_2_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_3_LC_1_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_3_LC_1_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32266),
            .lcout(RXbuffer_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_3C_net ),
            .ce(N__20510),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_4_LC_1_2_7 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_4_LC_1_2_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_4_LC_1_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_4_LC_1_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25538),
            .lcout(RXbuffer_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_3C_net ),
            .ce(N__20510),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_0_LC_1_4_0 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_0_LC_1_4_0 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_0_LC_1_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_0_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15850),
            .lcout(RXbuffer_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_0C_net ),
            .ce(N__20509),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_1_LC_1_4_1 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_1_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_1_LC_1_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_1_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41534),
            .lcout(RXbuffer_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_0C_net ),
            .ce(N__20509),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_2_LC_1_4_2 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_2_LC_1_4_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_2_LC_1_4_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \FTDI.RXbuffer_2_LC_1_4_2  (
            .in0(_gnd_net_),
            .in1(N__15813),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RXbuffer_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_0C_net ),
            .ce(N__20509),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_5_LC_1_4_5 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_5_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_5_LC_1_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_5_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16966),
            .lcout(RXbuffer_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_0C_net ),
            .ce(N__20509),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_6_LC_1_4_6 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_6_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_6_LC_1_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \FTDI.RXbuffer_6_LC_1_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15892),
            .lcout(RXbuffer_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_0C_net ),
            .ce(N__20509),
            .sr(_gnd_net_));
    defparam \FTDI.RXbuffer_7_LC_1_4_7 .C_ON=1'b0;
    defparam \FTDI.RXbuffer_7_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXbuffer_7_LC_1_4_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \FTDI.RXbuffer_7_LC_1_4_7  (
            .in0(N__21938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RXbuffer_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXbuffer_0C_net ),
            .ce(N__20509),
            .sr(_gnd_net_));
    defparam \ALU.f_8_LC_1_5_0 .C_ON=1'b0;
    defparam \ALU.f_8_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \ALU.f_8_LC_1_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_8_LC_1_5_0  (
            .in0(N__48261),
            .in1(N__47893),
            .in2(_gnd_net_),
            .in3(N__47808),
            .lcout(\ALU.fZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47674),
            .ce(N__36363),
            .sr(_gnd_net_));
    defparam \ALU.m198_LC_1_6_0 .C_ON=1'b0;
    defparam \ALU.m198_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.m198_LC_1_6_0 .LUT_INIT=16'b1101111110111011;
    LogicCell40 \ALU.m198_LC_1_6_0  (
            .in0(N__30200),
            .in1(N__29739),
            .in2(N__15185),
            .in3(N__25206),
            .lcout(\ALU.N_199_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_24_LC_1_6_1.C_ON=1'b0;
    defparam testWord_24_LC_1_6_1.SEQ_MODE=4'b1000;
    defparam testWord_24_LC_1_6_1.LUT_INIT=16'b1111011110000000;
    LogicCell40 testWord_24_LC_1_6_1 (
            .in0(N__41486),
            .in1(N__41201),
            .in2(N__15926),
            .in3(N__15184),
            .lcout(ctrlOut_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__41054),
            .sr(_gnd_net_));
    defparam testWord_8_LC_1_6_2.C_ON=1'b0;
    defparam testWord_8_LC_1_6_2.SEQ_MODE=4'b1000;
    defparam testWord_8_LC_1_6_2.LUT_INIT=16'b1100111011000100;
    LogicCell40 testWord_8_LC_1_6_2 (
            .in0(N__41204),
            .in1(N__26844),
            .in2(N__41508),
            .in3(N__15925),
            .lcout(testWordZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__41054),
            .sr(_gnd_net_));
    defparam testWord_25_LC_1_6_3.C_ON=1'b0;
    defparam testWord_25_LC_1_6_3.SEQ_MODE=4'b1000;
    defparam testWord_25_LC_1_6_3.LUT_INIT=16'b1111011110000000;
    LogicCell40 testWord_25_LC_1_6_3 (
            .in0(N__41487),
            .in1(N__41202),
            .in2(N__15862),
            .in3(N__19747),
            .lcout(ctrlOut_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__41054),
            .sr(_gnd_net_));
    defparam testWord_9_LC_1_6_4.C_ON=1'b0;
    defparam testWord_9_LC_1_6_4.SEQ_MODE=4'b1000;
    defparam testWord_9_LC_1_6_4.LUT_INIT=16'b1100111011000100;
    LogicCell40 testWord_9_LC_1_6_4 (
            .in0(N__41205),
            .in1(N__27155),
            .in2(N__41509),
            .in3(N__15857),
            .lcout(testWordZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__41054),
            .sr(_gnd_net_));
    defparam testWord_13_LC_1_6_5.C_ON=1'b0;
    defparam testWord_13_LC_1_6_5.SEQ_MODE=4'b1000;
    defparam testWord_13_LC_1_6_5.LUT_INIT=16'b1110001011110000;
    LogicCell40 testWord_13_LC_1_6_5 (
            .in0(N__25534),
            .in1(N__41490),
            .in2(N__15775),
            .in3(N__41199),
            .lcout(testWordZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__41054),
            .sr(_gnd_net_));
    defparam testWord_15_LC_1_6_6.C_ON=1'b0;
    defparam testWord_15_LC_1_6_6.SEQ_MODE=4'b1000;
    defparam testWord_15_LC_1_6_6.LUT_INIT=16'b1100111011000100;
    LogicCell40 testWord_15_LC_1_6_6 (
            .in0(N__41200),
            .in1(N__16810),
            .in2(N__41507),
            .in3(N__15897),
            .lcout(testWordZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__41054),
            .sr(_gnd_net_));
    defparam testWord_31_LC_1_6_7.C_ON=1'b0;
    defparam testWord_31_LC_1_6_7.SEQ_MODE=4'b1000;
    defparam testWord_31_LC_1_6_7.LUT_INIT=16'b1111011110000000;
    LogicCell40 testWord_31_LC_1_6_7 (
            .in0(N__41488),
            .in1(N__41203),
            .in2(N__15902),
            .in3(N__20940),
            .lcout(ctrlOut_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__41054),
            .sr(_gnd_net_));
    defparam testWord_21_LC_1_7_0.C_ON=1'b0;
    defparam testWord_21_LC_1_7_0.SEQ_MODE=4'b1000;
    defparam testWord_21_LC_1_7_0.LUT_INIT=16'b1110001010101010;
    LogicCell40 testWord_21_LC_1_7_0 (
            .in0(N__15227),
            .in1(N__41489),
            .in2(N__25545),
            .in3(N__18104),
            .lcout(ctrlOut_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47683),
            .ce(N__41053),
            .sr(_gnd_net_));
    defparam \ALU.m289_ns_1_LC_1_7_1 .C_ON=1'b0;
    defparam \ALU.m289_ns_1_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.m289_ns_1_LC_1_7_1 .LUT_INIT=16'b0001100000010000;
    LogicCell40 \ALU.m289_ns_1_LC_1_7_1  (
            .in0(N__30206),
            .in1(N__26568),
            .in2(N__29756),
            .in3(N__15225),
            .lcout(),
            .ltout(\ALU.m289_nsZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1K464_5_LC_1_7_2 .C_ON=1'b0;
    defparam \ALU.d_RNI1K464_5_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1K464_5_LC_1_7_2 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \ALU.d_RNI1K464_5_LC_1_7_2  (
            .in0(N__15226),
            .in1(N__29436),
            .in2(N__15173),
            .in3(N__40390),
            .lcout(\ALU.N_290_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m222_LC_1_7_3 .C_ON=1'b0;
    defparam \ALU.m222_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m222_LC_1_7_3 .LUT_INIT=16'b1110011111101111;
    LogicCell40 \ALU.m222_LC_1_7_3  (
            .in0(N__30205),
            .in1(N__25216),
            .in2(N__29755),
            .in3(N__15224),
            .lcout(\ALU.N_223_0 ),
            .ltout(\ALU.N_223_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVULB7_5_LC_1_7_4 .C_ON=1'b0;
    defparam \ALU.d_RNIVULB7_5_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVULB7_5_LC_1_7_4 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \ALU.d_RNIVULB7_5_LC_1_7_4  (
            .in0(N__24311),
            .in1(N__46942),
            .in2(N__15212),
            .in3(N__21728),
            .lcout(\ALU.a7_b_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINF4M7_3_LC_1_7_5 .C_ON=1'b0;
    defparam \ALU.d_RNINF4M7_3_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINF4M7_3_LC_1_7_5 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNINF4M7_3_LC_1_7_5  (
            .in0(N__23916),
            .in1(N__39849),
            .in2(N__24242),
            .in3(N__24044),
            .lcout(\ALU.a9_b_3 ),
            .ltout(\ALU.a9_b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_260_LC_1_7_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_260_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_260_LC_1_7_6 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \ALU.mult_madd_260_LC_1_7_6  (
            .in0(N__42687),
            .in1(N__40102),
            .in2(N__15209),
            .in3(N__15206),
            .lcout(\ALU.madd_260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_264_LC_1_7_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_264_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_264_LC_1_7_7 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_264_LC_1_7_7  (
            .in0(N__15205),
            .in1(N__40103),
            .in2(N__15197),
            .in3(N__42688),
            .lcout(\ALU.madd_264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_166_0_LC_1_8_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_166_0_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_166_0_LC_1_8_0 .LUT_INIT=16'b0011000010011010;
    LogicCell40 \ALU.mult_madd_166_0_LC_1_8_0  (
            .in0(N__46715),
            .in1(N__41737),
            .in2(N__46973),
            .in3(N__42690),
            .lcout(\ALU.madd_166_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_a3_2_0_LC_1_8_1 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_a3_2_0_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_a3_2_0_LC_1_8_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \ALU.mult_g0_0_a3_2_0_LC_1_8_1  (
            .in0(N__42692),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46956),
            .lcout(),
            .ltout(\ALU.g0_0_a3_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g2_0_0_LC_1_8_2 .C_ON=1'b0;
    defparam \ALU.mult_g2_0_0_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g2_0_0_LC_1_8_2 .LUT_INIT=16'b0101011001101010;
    LogicCell40 \ALU.mult_g2_0_0_LC_1_8_2  (
            .in0(N__18526),
            .in1(N__17516),
            .in2(N__15188),
            .in3(N__17543),
            .lcout(\ALU.g2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_2_LC_1_8_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_2_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_2_LC_1_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_0_2_LC_1_8_3  (
            .in0(N__17454),
            .in1(N__15239),
            .in2(N__17492),
            .in3(N__16049),
            .lcout(\ALU.g0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_315_0_LC_1_8_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_315_0_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_315_0_LC_1_8_4 .LUT_INIT=16'b0010001011010010;
    LogicCell40 \ALU.mult_madd_315_0_LC_1_8_4  (
            .in0(N__27598),
            .in1(N__41738),
            .in2(N__39854),
            .in3(N__42691),
            .lcout(\ALU.madd_315_0 ),
            .ltout(\ALU.madd_315_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_335_LC_1_8_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_335_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_335_LC_1_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_335_LC_1_8_5  (
            .in0(N__16027),
            .in1(N__15250),
            .in2(N__15269),
            .in3(N__15266),
            .lcout(\ALU.madd_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI8LNC7_12_LC_1_8_6 .C_ON=1'b0;
    defparam \ALU.c_RNI8LNC7_12_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI8LNC7_12_LC_1_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.c_RNI8LNC7_12_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__25355),
            .in2(_gnd_net_),
            .in3(N__37773),
            .lcout(\ALU.a12_b_1 ),
            .ltout(\ALU.a12_b_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_339_LC_1_8_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_339_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_339_LC_1_8_7 .LUT_INIT=16'b1011111000101000;
    LogicCell40 \ALU.mult_madd_339_LC_1_8_7  (
            .in0(N__16028),
            .in1(N__15260),
            .in2(N__15254),
            .in3(N__15251),
            .lcout(\ALU.madd_339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_5_LC_1_9_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_5_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_5_LC_1_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_g0_5_LC_1_9_0  (
            .in0(N__38315),
            .in1(N__25353),
            .in2(N__39608),
            .in3(N__36984),
            .lcout(),
            .ltout(\ALU.madd_141_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_4_LC_1_9_1 .C_ON=1'b0;
    defparam \ALU.mult_g0_4_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_4_LC_1_9_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_g0_4_LC_1_9_1  (
            .in0(N__37235),
            .in1(N__27600),
            .in2(N__15242),
            .in3(N__15304),
            .lcout(\ALU.N_1545_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_166_LC_1_9_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_166_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_166_LC_1_9_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ALU.mult_madd_166_LC_1_9_2  (
            .in0(N__15233),
            .in1(N__39850),
            .in2(_gnd_net_),
            .in3(N__37757),
            .lcout(\ALU.madd_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_252_LC_1_9_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_252_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_252_LC_1_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_252_LC_1_9_3  (
            .in0(N__36983),
            .in1(N__39600),
            .in2(N__25371),
            .in3(N__38311),
            .lcout(\ALU.madd_141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_254_0_tz_LC_1_9_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_254_0_tz_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_254_0_tz_LC_1_9_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ALU.mult_madd_254_0_tz_LC_1_9_4  (
            .in0(N__39601),
            .in1(N__25352),
            .in2(N__38336),
            .in3(N__36982),
            .lcout(\ALU.madd_254_0_tz ),
            .ltout(\ALU.madd_254_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_254_LC_1_9_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_254_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_254_LC_1_9_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \ALU.mult_madd_254_LC_1_9_5  (
            .in0(N__37234),
            .in1(N__27599),
            .in2(N__15317),
            .in3(N__15314),
            .lcout(\ALU.madd_254 ),
            .ltout(\ALU.madd_254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_340_0_LC_1_9_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_340_0_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_340_0_LC_1_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_340_0_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__17491),
            .in2(N__15308),
            .in3(N__17455),
            .lcout(\ALU.madd_340_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_1_LC_1_9_7 .C_ON=1'b0;
    defparam \ALU.mult_g0_1_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_1_LC_1_9_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_g0_1_LC_1_9_7  (
            .in0(N__15305),
            .in1(N__27601),
            .in2(N__17318),
            .in3(N__37236),
            .lcout(\ALU.N_1545_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFD4D4_3_LC_1_10_0 .C_ON=1'b0;
    defparam \ALU.d_RNIFD4D4_3_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFD4D4_3_LC_1_10_0 .LUT_INIT=16'b0000111101110111;
    LogicCell40 \ALU.d_RNIFD4D4_3_LC_1_10_0  (
            .in0(N__18053),
            .in1(N__29404),
            .in2(N__15293),
            .in3(N__42012),
            .lcout(\ALU.N_293_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_3_LC_1_10_1.C_ON=1'b0;
    defparam testWord_3_LC_1_10_1.SEQ_MODE=4'b1000;
    defparam testWord_3_LC_1_10_1.LUT_INIT=16'b1100110011100100;
    LogicCell40 testWord_3_LC_1_10_1 (
            .in0(N__18091),
            .in1(N__22203),
            .in2(N__15818),
            .in3(N__41506),
            .lcout(testWordZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47688),
            .ce(N__41052),
            .sr(_gnd_net_));
    defparam testWord_19_LC_1_10_2.C_ON=1'b0;
    defparam testWord_19_LC_1_10_2.SEQ_MODE=4'b1000;
    defparam testWord_19_LC_1_10_2.LUT_INIT=16'b1100101010101010;
    LogicCell40 testWord_19_LC_1_10_2 (
            .in0(N__18054),
            .in1(N__15814),
            .in2(N__41510),
            .in3(N__18090),
            .lcout(ctrlOut_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47688),
            .ce(N__41052),
            .sr(_gnd_net_));
    defparam \ALU.m292_ns_1_LC_1_10_3 .C_ON=1'b0;
    defparam \ALU.m292_ns_1_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m292_ns_1_LC_1_10_3 .LUT_INIT=16'b0100000000001010;
    LogicCell40 \ALU.m292_ns_1_LC_1_10_3  (
            .in0(N__29729),
            .in1(N__18052),
            .in2(N__26588),
            .in3(N__30195),
            .lcout(\ALU.m292_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m89_LC_1_10_4 .C_ON=1'b0;
    defparam \ALU.m89_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m89_LC_1_10_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ALU.m89_LC_1_10_4  (
            .in0(N__21902),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30323),
            .lcout(\ALU.N_90_0 ),
            .ltout(\ALU.N_90_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_22_LC_1_10_5.C_ON=1'b0;
    defparam testWord_22_LC_1_10_5.SEQ_MODE=4'b1000;
    defparam testWord_22_LC_1_10_5.LUT_INIT=16'b1011111110000000;
    LogicCell40 testWord_22_LC_1_10_5 (
            .in0(N__16985),
            .in1(N__41502),
            .in2(N__15284),
            .in3(N__15280),
            .lcout(ctrlOut_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47688),
            .ce(N__41052),
            .sr(_gnd_net_));
    defparam \ALU.m216_LC_1_10_6 .C_ON=1'b0;
    defparam \ALU.m216_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m216_LC_1_10_6 .LUT_INIT=16'b1110111001111111;
    LogicCell40 \ALU.m216_LC_1_10_6  (
            .in0(N__30194),
            .in1(N__25225),
            .in2(N__15281),
            .in3(N__29728),
            .lcout(\ALU.N_217_0 ),
            .ltout(\ALU.N_217_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIT7NA7_6_LC_1_10_7 .C_ON=1'b0;
    defparam \ALU.d_RNIT7NA7_6_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIT7NA7_6_LC_1_10_7 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \ALU.d_RNIT7NA7_6_LC_1_10_7  (
            .in0(N__29980),
            .in1(N__42958),
            .in2(N__15341),
            .in3(N__26727),
            .lcout(\ALU.a4_b_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1DA1A_10_LC_1_11_0 .C_ON=1'b0;
    defparam \ALU.d_RNI1DA1A_10_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1DA1A_10_LC_1_11_0 .LUT_INIT=16'b0001110111100010;
    LogicCell40 \ALU.d_RNI1DA1A_10_LC_1_11_0  (
            .in0(N__20023),
            .in1(N__26498),
            .in2(N__20065),
            .in3(N__27602),
            .lcout(),
            .ltout(\ALU.un9_addsub_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIV2S0F_10_LC_1_11_1 .C_ON=1'b0;
    defparam \ALU.a_RNIV2S0F_10_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIV2S0F_10_LC_1_11_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.a_RNIV2S0F_10_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15338),
            .in3(N__39571),
            .lcout(\ALU.a_RNIV2S0FZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILMFN5_10_LC_1_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNILMFN5_10_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILMFN5_10_LC_1_11_2 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \ALU.d_RNILMFN5_10_LC_1_11_2  (
            .in0(N__20024),
            .in1(_gnd_net_),
            .in2(N__20066),
            .in3(N__26497),
            .lcout(\ALU.N_192_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVRI59_10_LC_1_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIVRI59_10_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVRI59_10_LC_1_11_3 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \ALU.d_RNIVRI59_10_LC_1_11_3  (
            .in0(N__26499),
            .in1(N__41994),
            .in2(N__20108),
            .in3(N__20022),
            .lcout(),
            .ltout(\ALU.a3_b_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_15_LC_1_11_4 .C_ON=1'b0;
    defparam \ALU.mult_g0_15_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_15_LC_1_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_15_LC_1_11_4  (
            .in0(N__28274),
            .in1(N__15389),
            .in2(N__15335),
            .in3(N__18407),
            .lcout(),
            .ltout(\ALU.g0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_14_LC_1_11_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_14_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_14_LC_1_11_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_14_LC_1_11_5  (
            .in0(N__18458),
            .in1(N__15329),
            .in2(N__15332),
            .in3(N__19688),
            .lcout(\ALU.g0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_16_LC_1_11_6 .C_ON=1'b0;
    defparam \ALU.mult_g0_16_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_16_LC_1_11_6 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_g0_16_LC_1_11_6  (
            .in0(N__15323),
            .in1(_gnd_net_),
            .in2(N__18530),
            .in3(N__18557),
            .lcout(\ALU.N_1555_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_17_LC_1_12_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_17_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_17_LC_1_12_0 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_g0_17_LC_1_12_0  (
            .in0(N__39471),
            .in1(N__15445),
            .in2(N__18758),
            .in3(N__37937),
            .lcout(\ALU.N_1527_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_165_0_tz_LC_1_12_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_165_0_tz_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_165_0_tz_LC_1_12_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \ALU.mult_madd_165_0_tz_LC_1_12_1  (
            .in0(N__37934),
            .in1(N__39595),
            .in2(N__27586),
            .in3(N__38308),
            .lcout(\ALU.madd_165_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_163_LC_1_12_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_163_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_163_LC_1_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_163_LC_1_12_2  (
            .in0(N__38309),
            .in1(N__27534),
            .in2(N__39607),
            .in3(N__37935),
            .lcout(\ALU.madd_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_171_LC_1_12_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_171_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_171_LC_1_12_3 .LUT_INIT=16'b0010110111010010;
    LogicCell40 \ALU.mult_madd_171_LC_1_12_3  (
            .in0(N__41955),
            .in1(N__47089),
            .in2(N__16220),
            .in3(N__16208),
            .lcout(\ALU.madd_171 ),
            .ltout(\ALU.madd_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_190_LC_1_12_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_190_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_190_LC_1_12_4 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_madd_190_LC_1_12_4  (
            .in0(N__17590),
            .in1(N__15368),
            .in2(N__15374),
            .in3(N__15361),
            .lcout(\ALU.madd_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_161_0_LC_1_12_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_161_0_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_161_0_LC_1_12_5 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_161_0_LC_1_12_5  (
            .in0(N__37936),
            .in1(N__39599),
            .in2(N__40112),
            .in3(N__37195),
            .lcout(),
            .ltout(\ALU.madd_161_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_161_LC_1_12_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_161_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_161_LC_1_12_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ALU.mult_madd_161_LC_1_12_6  (
            .in0(N__38310),
            .in1(_gnd_net_),
            .in2(N__15371),
            .in3(N__27535),
            .lcout(\ALU.madd_161 ),
            .ltout(\ALU.madd_161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_186_LC_1_12_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_186_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_186_LC_1_12_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_186_LC_1_12_7  (
            .in0(N__15362),
            .in1(N__15350),
            .in2(N__15344),
            .in3(N__17591),
            .lcout(\ALU.madd_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_208_LC_1_13_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_208_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_208_LC_1_13_0 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \ALU.mult_madd_208_LC_1_13_0  (
            .in0(N__27595),
            .in1(N__15444),
            .in2(N__37758),
            .in3(N__21234),
            .lcout(\ALU.madd_208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIF74M7_3_LC_1_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIF74M7_3_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIF74M7_3_LC_1_13_1 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIF74M7_3_LC_1_13_1  (
            .in0(N__23944),
            .in1(N__40093),
            .in2(N__24312),
            .in3(N__24022),
            .lcout(\ALU.a8_b_3 ),
            .ltout(\ALU.a8_b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_212_LC_1_13_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_212_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_212_LC_1_13_2 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_212_LC_1_13_2  (
            .in0(N__27596),
            .in1(N__21235),
            .in2(N__15449),
            .in3(N__37731),
            .lcout(\ALU.madd_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_24_LC_1_13_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_24_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_24_LC_1_13_3 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_g0_24_LC_1_13_3  (
            .in0(N__37732),
            .in1(N__27597),
            .in2(N__21239),
            .in3(N__15446),
            .lcout(\ALU.N_1527_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_22_LC_1_13_4 .C_ON=1'b0;
    defparam \ALU.mult_g0_22_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_22_LC_1_13_4 .LUT_INIT=16'b0011011001101100;
    LogicCell40 \ALU.mult_g0_22_LC_1_13_4  (
            .in0(N__17251),
            .in1(N__15428),
            .in2(N__17270),
            .in3(N__17225),
            .lcout(),
            .ltout(\ALU.g0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_11_LC_1_13_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_11_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_11_LC_1_13_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_11_LC_1_13_5  (
            .in0(N__16253),
            .in1(N__16012),
            .in2(N__15419),
            .in3(N__15395),
            .lcout(\ALU.g0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_LC_1_13_6 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_LC_1_13_6 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \ALU.mult_g0_0_LC_1_13_6  (
            .in0(N__15416),
            .in1(N__16279),
            .in2(N__15410),
            .in3(N__16658),
            .lcout(\ALU.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_13_LC_1_14_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_13_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_13_LC_1_14_0 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_g0_13_LC_1_14_0  (
            .in0(N__39397),
            .in1(N__37199),
            .in2(N__40772),
            .in3(N__38317),
            .lcout(\ALU.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_10_ma_LC_1_14_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_10_ma_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_10_ma_LC_1_14_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_madd_cry_10_ma_LC_1_14_1  (
            .in0(N__15571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15586),
            .lcout(\ALU.madd_cry_10_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_124_0_LC_1_14_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_124_0_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_124_0_LC_1_14_2 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_124_0_LC_1_14_2  (
            .in0(N__39814),
            .in1(N__46918),
            .in2(N__37233),
            .in3(N__38316),
            .lcout(),
            .ltout(\ALU.madd_124_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_124_LC_1_14_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_124_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_124_LC_1_14_3 .LUT_INIT=16'b0111100001111000;
    LogicCell40 \ALU.mult_madd_124_LC_1_14_3  (
            .in0(N__37742),
            .in1(N__40094),
            .in2(N__15380),
            .in3(_gnd_net_),
            .lcout(\ALU.madd_124 ),
            .ltout(\ALU.madd_124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_144_LC_1_14_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_144_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_144_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_144_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__16637),
            .in2(N__15377),
            .in3(N__16796),
            .lcout(\ALU.madd_144 ),
            .ltout(\ALU.madd_144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_158_LC_1_14_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_158_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_158_LC_1_14_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_158_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__20354),
            .in2(N__15494),
            .in3(N__19355),
            .lcout(\ALU.madd_324 ),
            .ltout(\ALU.madd_324_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_9_l_ofx_LC_1_14_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_9_l_ofx_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_9_l_ofx_LC_1_14_6 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ALU.mult_madd_axb_9_l_ofx_LC_1_14_6  (
            .in0(N__19295),
            .in1(N__15570),
            .in2(N__15491),
            .in3(N__19277),
            .lcout(\ALU.madd_axb_9_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_134_LC_1_15_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_134_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_134_LC_1_15_0 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \ALU.mult_madd_134_LC_1_15_0  (
            .in0(N__23749),
            .in1(N__36994),
            .in2(N__15953),
            .in3(N__47051),
            .lcout(\ALU.madd_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_196_0_LC_1_15_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_196_0_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_196_0_LC_1_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_196_0_LC_1_15_1  (
            .in0(N__15477),
            .in1(N__16574),
            .in2(N__16595),
            .in3(N__16617),
            .lcout(),
            .ltout(\ALU.madd_N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m4_LC_1_15_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_m4_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m4_LC_1_15_2 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \ALU.mult_madd_m4_LC_1_15_2  (
            .in0(N__15476),
            .in1(N__20318),
            .in2(N__15488),
            .in3(N__16407),
            .lcout(\ALU.madd_N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_127_LC_1_15_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_127_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_127_LC_1_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_127_LC_1_15_3  (
            .in0(N__46911),
            .in1(N__37194),
            .in2(N__40120),
            .in3(N__37741),
            .lcout(\ALU.madd_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_196_LC_1_15_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_196_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_196_LC_1_15_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_196_LC_1_15_4  (
            .in0(N__16618),
            .in1(N__20524),
            .in2(N__15479),
            .in3(N__15485),
            .lcout(\ALU.madd_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_191_0_LC_1_15_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_191_0_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_191_0_LC_1_15_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.mult_madd_191_0_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__16573),
            .in2(_gnd_net_),
            .in3(N__16591),
            .lcout(\ALU.madd_191_0 ),
            .ltout(\ALU.madd_191_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_200_LC_1_15_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_200_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_200_LC_1_15_6 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \ALU.mult_madd_200_LC_1_15_6  (
            .in0(N__16619),
            .in1(N__15478),
            .in2(N__15452),
            .in3(N__20525),
            .lcout(\ALU.madd_326 ),
            .ltout(\ALU.madd_326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_10_l_ofx_LC_1_15_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_10_l_ofx_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_10_l_ofx_LC_1_15_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \ALU.mult_madd_axb_10_l_ofx_LC_1_15_7  (
            .in0(N__16408),
            .in1(N__15587),
            .in2(N__15575),
            .in3(N__15572),
            .lcout(\ALU.madd_axb_10_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_0_LC_1_16_0.C_ON=1'b1;
    defparam clkdiv_0_LC_1_16_0.SEQ_MODE=4'b1000;
    defparam clkdiv_0_LC_1_16_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_0_LC_1_16_0 (
            .in0(_gnd_net_),
            .in1(N__15557),
            .in2(_gnd_net_),
            .in3(N__15551),
            .lcout(clkdivZ0Z_0),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(clkdiv_cry_0),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_1_LC_1_16_1.C_ON=1'b1;
    defparam clkdiv_1_LC_1_16_1.SEQ_MODE=4'b1000;
    defparam clkdiv_1_LC_1_16_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_1_LC_1_16_1 (
            .in0(_gnd_net_),
            .in1(N__15548),
            .in2(_gnd_net_),
            .in3(N__15542),
            .lcout(clkdivZ0Z_1),
            .ltout(),
            .carryin(clkdiv_cry_0),
            .carryout(clkdiv_cry_1),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_2_LC_1_16_2.C_ON=1'b1;
    defparam clkdiv_2_LC_1_16_2.SEQ_MODE=4'b1000;
    defparam clkdiv_2_LC_1_16_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_2_LC_1_16_2 (
            .in0(_gnd_net_),
            .in1(N__15539),
            .in2(_gnd_net_),
            .in3(N__15533),
            .lcout(clkdivZ0Z_2),
            .ltout(),
            .carryin(clkdiv_cry_1),
            .carryout(clkdiv_cry_2),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_3_LC_1_16_3.C_ON=1'b1;
    defparam clkdiv_3_LC_1_16_3.SEQ_MODE=4'b1000;
    defparam clkdiv_3_LC_1_16_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_3_LC_1_16_3 (
            .in0(_gnd_net_),
            .in1(N__15530),
            .in2(_gnd_net_),
            .in3(N__15524),
            .lcout(clkdivZ0Z_3),
            .ltout(),
            .carryin(clkdiv_cry_2),
            .carryout(clkdiv_cry_3),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_4_LC_1_16_4.C_ON=1'b1;
    defparam clkdiv_4_LC_1_16_4.SEQ_MODE=4'b1000;
    defparam clkdiv_4_LC_1_16_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_4_LC_1_16_4 (
            .in0(_gnd_net_),
            .in1(N__15521),
            .in2(_gnd_net_),
            .in3(N__15515),
            .lcout(clkdivZ0Z_4),
            .ltout(),
            .carryin(clkdiv_cry_3),
            .carryout(clkdiv_cry_4),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_5_LC_1_16_5.C_ON=1'b1;
    defparam clkdiv_5_LC_1_16_5.SEQ_MODE=4'b1000;
    defparam clkdiv_5_LC_1_16_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_5_LC_1_16_5 (
            .in0(_gnd_net_),
            .in1(N__15512),
            .in2(_gnd_net_),
            .in3(N__15506),
            .lcout(clkdivZ0Z_5),
            .ltout(),
            .carryin(clkdiv_cry_4),
            .carryout(clkdiv_cry_5),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_6_LC_1_16_6.C_ON=1'b1;
    defparam clkdiv_6_LC_1_16_6.SEQ_MODE=4'b1000;
    defparam clkdiv_6_LC_1_16_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_6_LC_1_16_6 (
            .in0(_gnd_net_),
            .in1(N__15503),
            .in2(_gnd_net_),
            .in3(N__15497),
            .lcout(clkdivZ0Z_6),
            .ltout(),
            .carryin(clkdiv_cry_5),
            .carryout(clkdiv_cry_6),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_7_LC_1_16_7.C_ON=1'b1;
    defparam clkdiv_7_LC_1_16_7.SEQ_MODE=4'b1000;
    defparam clkdiv_7_LC_1_16_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_7_LC_1_16_7 (
            .in0(_gnd_net_),
            .in1(N__15668),
            .in2(_gnd_net_),
            .in3(N__15662),
            .lcout(clkdivZ0Z_7),
            .ltout(),
            .carryin(clkdiv_cry_6),
            .carryout(clkdiv_cry_7),
            .clk(N__47691),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_8_LC_1_17_0.C_ON=1'b1;
    defparam clkdiv_8_LC_1_17_0.SEQ_MODE=4'b1000;
    defparam clkdiv_8_LC_1_17_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_8_LC_1_17_0 (
            .in0(_gnd_net_),
            .in1(N__15659),
            .in2(_gnd_net_),
            .in3(N__15653),
            .lcout(clkdivZ0Z_8),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(clkdiv_cry_8),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_9_LC_1_17_1.C_ON=1'b1;
    defparam clkdiv_9_LC_1_17_1.SEQ_MODE=4'b1000;
    defparam clkdiv_9_LC_1_17_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_9_LC_1_17_1 (
            .in0(_gnd_net_),
            .in1(N__15650),
            .in2(_gnd_net_),
            .in3(N__15644),
            .lcout(clkdivZ0Z_9),
            .ltout(),
            .carryin(clkdiv_cry_8),
            .carryout(clkdiv_cry_9),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_10_LC_1_17_2.C_ON=1'b1;
    defparam clkdiv_10_LC_1_17_2.SEQ_MODE=4'b1000;
    defparam clkdiv_10_LC_1_17_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_10_LC_1_17_2 (
            .in0(_gnd_net_),
            .in1(N__15641),
            .in2(_gnd_net_),
            .in3(N__15635),
            .lcout(clkdivZ0Z_10),
            .ltout(),
            .carryin(clkdiv_cry_9),
            .carryout(clkdiv_cry_10),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_11_LC_1_17_3.C_ON=1'b1;
    defparam clkdiv_11_LC_1_17_3.SEQ_MODE=4'b1000;
    defparam clkdiv_11_LC_1_17_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_11_LC_1_17_3 (
            .in0(_gnd_net_),
            .in1(N__15632),
            .in2(_gnd_net_),
            .in3(N__15626),
            .lcout(clkdivZ0Z_11),
            .ltout(),
            .carryin(clkdiv_cry_10),
            .carryout(clkdiv_cry_11),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_12_LC_1_17_4.C_ON=1'b1;
    defparam clkdiv_12_LC_1_17_4.SEQ_MODE=4'b1000;
    defparam clkdiv_12_LC_1_17_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_12_LC_1_17_4 (
            .in0(_gnd_net_),
            .in1(N__15623),
            .in2(_gnd_net_),
            .in3(N__15617),
            .lcout(clkdivZ0Z_12),
            .ltout(),
            .carryin(clkdiv_cry_11),
            .carryout(clkdiv_cry_12),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_13_LC_1_17_5.C_ON=1'b1;
    defparam clkdiv_13_LC_1_17_5.SEQ_MODE=4'b1000;
    defparam clkdiv_13_LC_1_17_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_13_LC_1_17_5 (
            .in0(_gnd_net_),
            .in1(N__15614),
            .in2(_gnd_net_),
            .in3(N__15608),
            .lcout(clkdivZ0Z_13),
            .ltout(),
            .carryin(clkdiv_cry_12),
            .carryout(clkdiv_cry_13),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_14_LC_1_17_6.C_ON=1'b1;
    defparam clkdiv_14_LC_1_17_6.SEQ_MODE=4'b1000;
    defparam clkdiv_14_LC_1_17_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_14_LC_1_17_6 (
            .in0(_gnd_net_),
            .in1(N__15605),
            .in2(_gnd_net_),
            .in3(N__15599),
            .lcout(clkdivZ0Z_14),
            .ltout(),
            .carryin(clkdiv_cry_13),
            .carryout(clkdiv_cry_14),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_15_LC_1_17_7.C_ON=1'b1;
    defparam clkdiv_15_LC_1_17_7.SEQ_MODE=4'b1000;
    defparam clkdiv_15_LC_1_17_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_15_LC_1_17_7 (
            .in0(_gnd_net_),
            .in1(N__15596),
            .in2(_gnd_net_),
            .in3(N__15590),
            .lcout(clkdivZ0Z_15),
            .ltout(),
            .carryin(clkdiv_cry_14),
            .carryout(clkdiv_cry_15),
            .clk(N__47692),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_16_LC_1_18_0.C_ON=1'b1;
    defparam clkdiv_16_LC_1_18_0.SEQ_MODE=4'b1000;
    defparam clkdiv_16_LC_1_18_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_16_LC_1_18_0 (
            .in0(_gnd_net_),
            .in1(N__15752),
            .in2(_gnd_net_),
            .in3(N__15746),
            .lcout(clkdivZ0Z_16),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(clkdiv_cry_16),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_17_LC_1_18_1.C_ON=1'b1;
    defparam clkdiv_17_LC_1_18_1.SEQ_MODE=4'b1000;
    defparam clkdiv_17_LC_1_18_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_17_LC_1_18_1 (
            .in0(_gnd_net_),
            .in1(N__15743),
            .in2(_gnd_net_),
            .in3(N__15737),
            .lcout(clkdivZ0Z_17),
            .ltout(),
            .carryin(clkdiv_cry_16),
            .carryout(clkdiv_cry_17),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_18_LC_1_18_2.C_ON=1'b1;
    defparam clkdiv_18_LC_1_18_2.SEQ_MODE=4'b1000;
    defparam clkdiv_18_LC_1_18_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_18_LC_1_18_2 (
            .in0(_gnd_net_),
            .in1(N__15734),
            .in2(_gnd_net_),
            .in3(N__15728),
            .lcout(clkdivZ0Z_18),
            .ltout(),
            .carryin(clkdiv_cry_17),
            .carryout(clkdiv_cry_18),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_19_LC_1_18_3.C_ON=1'b1;
    defparam clkdiv_19_LC_1_18_3.SEQ_MODE=4'b1000;
    defparam clkdiv_19_LC_1_18_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_19_LC_1_18_3 (
            .in0(_gnd_net_),
            .in1(N__15725),
            .in2(_gnd_net_),
            .in3(N__15719),
            .lcout(clkdivZ0Z_19),
            .ltout(),
            .carryin(clkdiv_cry_18),
            .carryout(clkdiv_cry_19),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_20_LC_1_18_4.C_ON=1'b1;
    defparam clkdiv_20_LC_1_18_4.SEQ_MODE=4'b1000;
    defparam clkdiv_20_LC_1_18_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_20_LC_1_18_4 (
            .in0(_gnd_net_),
            .in1(N__15716),
            .in2(_gnd_net_),
            .in3(N__15710),
            .lcout(clkdivZ0Z_20),
            .ltout(),
            .carryin(clkdiv_cry_19),
            .carryout(clkdiv_cry_20),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_21_LC_1_18_5.C_ON=1'b1;
    defparam clkdiv_21_LC_1_18_5.SEQ_MODE=4'b1000;
    defparam clkdiv_21_LC_1_18_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_21_LC_1_18_5 (
            .in0(_gnd_net_),
            .in1(N__15707),
            .in2(_gnd_net_),
            .in3(N__15701),
            .lcout(clkdivZ0Z_21),
            .ltout(),
            .carryin(clkdiv_cry_20),
            .carryout(clkdiv_cry_21),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_22_LC_1_18_6.C_ON=1'b1;
    defparam clkdiv_22_LC_1_18_6.SEQ_MODE=4'b1000;
    defparam clkdiv_22_LC_1_18_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clkdiv_22_LC_1_18_6 (
            .in0(_gnd_net_),
            .in1(N__15698),
            .in2(_gnd_net_),
            .in3(N__15692),
            .lcout(clkdivZ0Z_22),
            .ltout(),
            .carryin(clkdiv_cry_21),
            .carryout(clkdiv_cry_22),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam clkdiv_23_LC_1_18_7.C_ON=1'b0;
    defparam clkdiv_23_LC_1_18_7.SEQ_MODE=4'b1000;
    defparam clkdiv_23_LC_1_18_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 clkdiv_23_LC_1_18_7 (
            .in0(_gnd_net_),
            .in1(N__15679),
            .in2(_gnd_net_),
            .in3(N__15689),
            .lcout(GPIO3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47693),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.results_e_0_0_LC_2_1_0 .C_ON=1'b0;
    defparam \CONTROL.results_e_0_0_LC_2_1_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.results_e_0_0_LC_2_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.results_e_0_0_LC_2_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15782),
            .lcout(aluResults_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47642),
            .ce(N__16847),
            .sr(_gnd_net_));
    defparam testWord_18_LC_2_2_0.C_ON=1'b0;
    defparam testWord_18_LC_2_2_0.SEQ_MODE=4'b1000;
    defparam testWord_18_LC_2_2_0.LUT_INIT=16'b1110001010101010;
    LogicCell40 testWord_18_LC_2_2_0 (
            .in0(N__20277),
            .in1(N__41431),
            .in2(N__41544),
            .in3(N__18120),
            .lcout(ctrlOut_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47648),
            .ce(N__41059),
            .sr(_gnd_net_));
    defparam \ALU.m304_ns_1_LC_2_2_1 .C_ON=1'b0;
    defparam \ALU.m304_ns_1_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.m304_ns_1_LC_2_2_1 .LUT_INIT=16'b0001010111110101;
    LogicCell40 \ALU.m304_ns_1_LC_2_2_1  (
            .in0(N__22402),
            .in1(N__22687),
            .in2(N__33300),
            .in3(N__20276),
            .lcout(),
            .ltout(\ALU.m304_nsZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m304_ns_LC_2_2_2 .C_ON=1'b0;
    defparam \ALU.m304_ns_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.m304_ns_LC_2_2_2 .LUT_INIT=16'b1010011011110111;
    LogicCell40 \ALU.m304_ns_LC_2_2_2  (
            .in0(N__33261),
            .in1(N__22280),
            .in2(N__15758),
            .in3(N__38733),
            .lcout(N_305_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_2_LC_2_2_3.C_ON=1'b0;
    defparam testWord_2_LC_2_2_3.SEQ_MODE=4'b1000;
    defparam testWord_2_LC_2_2_3.LUT_INIT=16'b1111110100001000;
    LogicCell40 testWord_2_LC_2_2_3 (
            .in0(N__18122),
            .in1(N__41538),
            .in2(N__41475),
            .in3(N__22409),
            .lcout(testWordZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47648),
            .ce(N__41059),
            .sr(_gnd_net_));
    defparam testWord_1_LC_2_2_4.C_ON=1'b0;
    defparam testWord_1_LC_2_2_4.SEQ_MODE=4'b1000;
    defparam testWord_1_LC_2_2_4.LUT_INIT=16'b1011100010101010;
    LogicCell40 testWord_1_LC_2_2_4 (
            .in0(N__22692),
            .in1(N__41430),
            .in2(N__15863),
            .in3(N__18121),
            .lcout(testWordZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47648),
            .ce(N__41059),
            .sr(_gnd_net_));
    defparam testWord_5_LC_2_2_5.C_ON=1'b0;
    defparam testWord_5_LC_2_2_5.SEQ_MODE=4'b1000;
    defparam testWord_5_LC_2_2_5.LUT_INIT=16'b1111110100001000;
    LogicCell40 testWord_5_LC_2_2_5 (
            .in0(N__18123),
            .in1(N__25546),
            .in2(N__41476),
            .in3(N__33263),
            .lcout(testWordZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47648),
            .ce(N__41059),
            .sr(_gnd_net_));
    defparam \ALU.m656_LC_2_2_6 .C_ON=1'b0;
    defparam \ALU.m656_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m656_LC_2_2_6 .LUT_INIT=16'b0100011101111100;
    LogicCell40 \ALU.m656_LC_2_2_6  (
            .in0(N__21568),
            .in1(N__33259),
            .in2(N__22719),
            .in3(N__22403),
            .lcout(),
            .ltout(\ALU.i73_mux_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m657_LC_2_2_7 .C_ON=1'b0;
    defparam \ALU.m657_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m657_LC_2_2_7 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \ALU.m657_LC_2_2_7  (
            .in0(N__22281),
            .in1(N__33262),
            .in2(N__15755),
            .in3(N__22691),
            .lcout(i53_mux_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_8_LC_2_3_0 .C_ON=1'b0;
    defparam \ALU.g_8_LC_2_3_0 .SEQ_MODE=4'b1000;
    defparam \ALU.g_8_LC_2_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_8_LC_2_3_0  (
            .in0(N__48109),
            .in1(N__47894),
            .in2(_gnd_net_),
            .in3(N__47809),
            .lcout(\ALU.gZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47655),
            .ce(N__36069),
            .sr(_gnd_net_));
    defparam testWord_16_LC_2_4_0.C_ON=1'b0;
    defparam testWord_16_LC_2_4_0.SEQ_MODE=4'b1000;
    defparam testWord_16_LC_2_4_0.LUT_INIT=16'b1111011110000000;
    LogicCell40 testWord_16_LC_2_4_0 (
            .in0(N__41423),
            .in1(N__18139),
            .in2(N__15921),
            .in3(N__21564),
            .lcout(ctrlOut_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(N__41058),
            .sr(_gnd_net_));
    defparam testWord_23_LC_2_4_1.C_ON=1'b0;
    defparam testWord_23_LC_2_4_1.SEQ_MODE=4'b1000;
    defparam testWord_23_LC_2_4_1.LUT_INIT=16'b1111011110000000;
    LogicCell40 testWord_23_LC_2_4_1 (
            .in0(N__18141),
            .in1(N__41425),
            .in2(N__15901),
            .in3(N__19867),
            .lcout(ctrlOut_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(N__41058),
            .sr(_gnd_net_));
    defparam testWord_7_LC_2_4_2.C_ON=1'b0;
    defparam testWord_7_LC_2_4_2.SEQ_MODE=4'b1000;
    defparam testWord_7_LC_2_4_2.LUT_INIT=16'b1110001011110000;
    LogicCell40 testWord_7_LC_2_4_2 (
            .in0(N__15896),
            .in1(N__41429),
            .in2(N__27745),
            .in3(N__18143),
            .lcout(testWordZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(N__41058),
            .sr(_gnd_net_));
    defparam testWord_17_LC_2_4_3.C_ON=1'b0;
    defparam testWord_17_LC_2_4_3.SEQ_MODE=4'b1000;
    defparam testWord_17_LC_2_4_3.LUT_INIT=16'b1111011110000000;
    LogicCell40 testWord_17_LC_2_4_3 (
            .in0(N__18140),
            .in1(N__41424),
            .in2(N__15861),
            .in3(N__21846),
            .lcout(ctrlOut_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(N__41058),
            .sr(_gnd_net_));
    defparam testWord_4_LC_2_4_4.C_ON=1'b0;
    defparam testWord_4_LC_2_4_4.SEQ_MODE=4'b1000;
    defparam testWord_4_LC_2_4_4.LUT_INIT=16'b1011100010101010;
    LogicCell40 testWord_4_LC_2_4_4 (
            .in0(N__22504),
            .in1(N__41428),
            .in2(N__32291),
            .in3(N__18142),
            .lcout(testWordZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(N__41058),
            .sr(_gnd_net_));
    defparam testWord_11_LC_2_4_6.C_ON=1'b0;
    defparam testWord_11_LC_2_4_6.SEQ_MODE=4'b1000;
    defparam testWord_11_LC_2_4_6.LUT_INIT=16'b1110001011110000;
    LogicCell40 testWord_11_LC_2_4_6 (
            .in0(N__15811),
            .in1(N__41427),
            .in2(N__34545),
            .in3(N__41206),
            .lcout(testWordZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(N__41058),
            .sr(_gnd_net_));
    defparam testWord_27_LC_2_4_7.C_ON=1'b0;
    defparam testWord_27_LC_2_4_7.SEQ_MODE=4'b1000;
    defparam testWord_27_LC_2_4_7.LUT_INIT=16'b1111100001110000;
    LogicCell40 testWord_27_LC_2_4_7 (
            .in0(N__41207),
            .in1(N__41426),
            .in2(N__24892),
            .in3(N__15812),
            .lcout(ctrlOut_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(N__41058),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_rep2_e_LC_2_5_0 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_rep2_e_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluReadBus_rep2_e_LC_2_5_0 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \CONTROL.aluReadBus_rep2_e_LC_2_5_0  (
            .in0(N__33296),
            .in1(N__19576),
            .in2(N__19540),
            .in3(N__22257),
            .lcout(aluReadBus_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47668),
            .ce(N__34710),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_N_3L3_LC_2_5_1 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_N_3L3_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_N_3L3_LC_2_5_1 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.mult_g0_0_0_N_3L3_LC_2_5_1  (
            .in0(N__21097),
            .in1(N__32738),
            .in2(N__29898),
            .in3(N__37484),
            .lcout(\ALU.g0_0_0_N_3L3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_e_0_LC_2_5_2 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_e_0_LC_2_5_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluReadBus_e_0_LC_2_5_2 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \CONTROL.aluReadBus_e_0_LC_2_5_2  (
            .in0(N__33295),
            .in1(N__19575),
            .in2(N__19539),
            .in3(N__22256),
            .lcout(aluReadBus),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47668),
            .ce(N__34710),
            .sr(_gnd_net_));
    defparam \ALU.m8_LC_2_5_3 .C_ON=1'b0;
    defparam \ALU.m8_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m8_LC_2_5_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \ALU.m8_LC_2_5_3  (
            .in0(N__29837),
            .in1(_gnd_net_),
            .in2(N__30217),
            .in3(N__29746),
            .lcout(\ALU.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m660_LC_2_5_4 .C_ON=1'b0;
    defparam \ALU.m660_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m660_LC_2_5_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \ALU.m660_LC_2_5_4  (
            .in0(N__22492),
            .in1(N__22430),
            .in2(_gnd_net_),
            .in3(N__22255),
            .lcout(),
            .ltout(N_661_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_cnv_0_LC_2_5_5 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_cnv_0_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_cnv_0_LC_2_5_5 .LUT_INIT=16'b1000101100000000;
    LogicCell40 \CONTROL.aluOperation_cnv_0_LC_2_5_5  (
            .in0(N__16871),
            .in1(N__33294),
            .in2(N__15932),
            .in3(N__34668),
            .lcout(\CONTROL.aluOperation_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m9_LC_2_5_6 .C_ON=1'b0;
    defparam \ALU.m9_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m9_LC_2_5_6 .LUT_INIT=16'b1011101111011101;
    LogicCell40 \ALU.m9_LC_2_5_6  (
            .in0(N__29745),
            .in1(N__30207),
            .in2(_gnd_net_),
            .in3(N__29836),
            .lcout(\ALU.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m634_LC_2_5_7 .C_ON=1'b0;
    defparam \ALU.m634_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m634_LC_2_5_7 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \ALU.m634_LC_2_5_7  (
            .in0(N__22431),
            .in1(N__22493),
            .in2(_gnd_net_),
            .in3(N__22720),
            .lcout(\ALU.N_635_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIR21R7_8_LC_2_6_0 .C_ON=1'b0;
    defparam \ALU.d_RNIR21R7_8_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIR21R7_8_LC_2_6_0 .LUT_INIT=16'b0011101011000101;
    LogicCell40 \ALU.d_RNIR21R7_8_LC_2_6_0  (
            .in0(N__18728),
            .in1(N__18627),
            .in2(N__26535),
            .in3(N__40079),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQ74VB_8_LC_2_6_1 .C_ON=1'b0;
    defparam \ALU.d_RNIQ74VB_8_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQ74VB_8_LC_2_6_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNIQ74VB_8_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15929),
            .in3(N__21484),
            .lcout(\ALU.d_RNIQ74VBZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN2L24_8_LC_2_6_2 .C_ON=1'b0;
    defparam \ALU.d_RNIN2L24_8_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN2L24_8_LC_2_6_2 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \ALU.d_RNIN2L24_8_LC_2_6_2  (
            .in0(N__18729),
            .in1(_gnd_net_),
            .in2(N__26536),
            .in3(N__18628),
            .lcout(\ALU.N_201_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI60794_8_LC_2_6_3 .C_ON=1'b0;
    defparam \ALU.d_RNI60794_8_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI60794_8_LC_2_6_3 .LUT_INIT=16'b1111000011110101;
    LogicCell40 \ALU.d_RNI60794_8_LC_2_6_3  (
            .in0(N__40080),
            .in1(_gnd_net_),
            .in2(N__18648),
            .in3(N__29435),
            .lcout(),
            .ltout(\ALU.N_275_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIUSVB61_8_LC_2_6_4 .C_ON=1'b0;
    defparam \ALU.d_RNIUSVB61_8_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIUSVB61_8_LC_2_6_4 .LUT_INIT=16'b0100011100000011;
    LogicCell40 \ALU.d_RNIUSVB61_8_LC_2_6_4  (
            .in0(N__44448),
            .in1(N__43165),
            .in2(N__15977),
            .in3(N__19385),
            .lcout(\ALU.a_15_m3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_N_4L5_LC_2_6_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_N_4L5_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_N_4L5_LC_2_6_5 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_g0_0_0_N_4L5_LC_2_6_5  (
            .in0(N__27593),
            .in1(N__37244),
            .in2(N__40107),
            .in3(N__38332),
            .lcout(),
            .ltout(\ALU.g0_0_0_N_4L5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_LC_2_6_6 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_LC_2_6_6 .LUT_INIT=16'b1110100010001110;
    LogicCell40 \ALU.mult_g0_0_0_LC_2_6_6  (
            .in0(N__15974),
            .in1(N__15965),
            .in2(N__15968),
            .in3(N__21617),
            .lcout(\ALU.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_N_3L3_0_LC_2_6_7 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_N_3L3_0_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_N_3L3_0_LC_2_6_7 .LUT_INIT=16'b0100111000000000;
    LogicCell40 \ALU.mult_g0_0_0_N_3L3_0_LC_2_6_7  (
            .in0(N__24325),
            .in1(N__18727),
            .in2(N__18647),
            .in3(N__36995),
            .lcout(\ALU.g0_0_0_N_3L3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRAM58_9_LC_2_7_0 .C_ON=1'b0;
    defparam \ALU.d_RNIRAM58_9_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRAM58_9_LC_2_7_0 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNIRAM58_9_LC_2_7_0  (
            .in0(N__21089),
            .in1(N__20868),
            .in2(N__30023),
            .in3(N__40388),
            .lcout(\ALU.a5_b_9 ),
            .ltout(\ALU.a5_b_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_382_LC_2_7_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_382_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_382_LC_2_7_1 .LUT_INIT=16'b0110100100111100;
    LogicCell40 \ALU.mult_madd_382_LC_2_7_1  (
            .in0(N__47099),
            .in1(N__18196),
            .in2(N__15959),
            .in3(N__46944),
            .lcout(\ALU.madd_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVPQD3_8_LC_2_7_2 .C_ON=1'b0;
    defparam \ALU.d_RNIVPQD3_8_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVPQD3_8_LC_2_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIVPQD3_8_LC_2_7_2  (
            .in0(N__32996),
            .in1(N__25604),
            .in2(_gnd_net_),
            .in3(N__30875),
            .lcout(\ALU.operand2_8 ),
            .ltout(\ALU.operand2_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC54P6_8_LC_2_7_3 .C_ON=1'b0;
    defparam \ALU.d_RNIC54P6_8_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC54P6_8_LC_2_7_3 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \ALU.d_RNIC54P6_8_LC_2_7_3  (
            .in0(N__24232),
            .in1(N__18614),
            .in2(N__15956),
            .in3(N__37447),
            .lcout(\ALU.a1_b_8 ),
            .ltout(\ALU.a1_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_138_LC_2_7_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_138_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_138_LC_2_7_4 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_138_LC_2_7_4  (
            .in0(N__23750),
            .in1(N__36996),
            .in2(N__15935),
            .in3(N__47097),
            .lcout(\ALU.madd_138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGG5I7_8_LC_2_7_5 .C_ON=1'b0;
    defparam \ALU.d_RNIGG5I7_8_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGG5I7_8_LC_2_7_5 .LUT_INIT=16'b0100111000000000;
    LogicCell40 \ALU.d_RNIGG5I7_8_LC_2_7_5  (
            .in0(N__24233),
            .in1(N__18716),
            .in2(N__18640),
            .in3(N__42959),
            .lcout(),
            .ltout(\ALU.a4_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_269_LC_2_7_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_269_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_269_LC_2_7_6 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_269_LC_2_7_6  (
            .in0(N__23783),
            .in1(N__40389),
            .in2(N__16031),
            .in3(N__47098),
            .lcout(\ALU.madd_269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2AVH7_8_LC_2_7_7 .C_ON=1'b0;
    defparam \ALU.d_RNI2AVH7_8_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2AVH7_8_LC_2_7_7 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNI2AVH7_8_LC_2_7_7  (
            .in0(N__18618),
            .in1(N__18717),
            .in2(N__30024),
            .in3(N__46736),
            .lcout(\ALU.a6_b_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m3_1_LC_2_8_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_m3_1_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m3_1_LC_2_8_0 .LUT_INIT=16'b0010000110110111;
    LogicCell40 \ALU.mult_madd_m3_1_LC_2_8_0  (
            .in0(N__17575),
            .in1(N__16686),
            .in2(N__16537),
            .in3(N__16768),
            .lcout(),
            .ltout(\ALU.madd_i1_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m6_0_LC_2_8_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_m6_0_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m6_0_LC_2_8_1 .LUT_INIT=16'b0011000011110011;
    LogicCell40 \ALU.mult_madd_m6_0_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__18569),
            .in2(N__16019),
            .in3(N__16283),
            .lcout(),
            .ltout(\ALU.madd_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_LC_2_8_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_LC_2_8_2 .LUT_INIT=16'b0100110110001110;
    LogicCell40 \ALU.mult_madd_LC_2_8_2  (
            .in0(N__16061),
            .in1(N__16016),
            .in2(N__15995),
            .in3(N__16139),
            .lcout(\ALU.madd_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_LC_2_8_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_LC_2_8_3 .LUT_INIT=16'b0101011001101010;
    LogicCell40 \ALU.mult_madd_484_LC_2_8_3  (
            .in0(N__17042),
            .in1(N__17414),
            .in2(N__18440),
            .in3(N__17087),
            .lcout(),
            .ltout(\ALU.madd_331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_14_LC_2_8_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_14_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_14_LC_2_8_4 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ALU.mult_madd_axb_14_LC_2_8_4  (
            .in0(N__17354),
            .in1(N__15988),
            .in2(N__15992),
            .in3(N__17324),
            .lcout(\ALU.madd_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_13_l_ofx_LC_2_8_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_13_l_ofx_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_13_l_ofx_LC_2_8_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_axb_13_l_ofx_LC_2_8_5  (
            .in0(N__16349),
            .in1(N__16376),
            .in2(N__15989),
            .in3(N__17353),
            .lcout(\ALU.madd_axb_13_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_237_LC_2_8_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_237_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_237_LC_2_8_6 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \ALU.mult_madd_237_LC_2_8_6  (
            .in0(N__17576),
            .in1(N__16685),
            .in2(N__16538),
            .in3(N__16769),
            .lcout(\ALU.madd_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_325_0_LC_2_9_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_325_0_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_325_0_LC_2_9_0 .LUT_INIT=16'b0110001101010000;
    LogicCell40 \ALU.mult_madd_325_0_LC_2_9_0  (
            .in0(N__22048),
            .in1(N__21444),
            .in2(N__42990),
            .in3(N__40432),
            .lcout(\ALU.madd_325_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_354_LC_2_9_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_354_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_354_LC_2_9_1 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \ALU.mult_madd_354_LC_2_9_1  (
            .in0(N__16051),
            .in1(N__17186),
            .in2(N__16138),
            .in3(N__16085),
            .lcout(\ALU.madd_354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g2_LC_2_9_2 .C_ON=1'b0;
    defparam \ALU.mult_g2_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g2_LC_2_9_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ALU.mult_g2_LC_2_9_2  (
            .in0(N__40084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28084),
            .lcout(\ALU.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_10_LC_2_9_3 .C_ON=1'b0;
    defparam \ALU.mult_g0_10_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_10_LC_2_9_3 .LUT_INIT=16'b0000101011000110;
    LogicCell40 \ALU.mult_g0_10_LC_2_9_3  (
            .in0(N__40431),
            .in1(N__42957),
            .in2(N__21469),
            .in3(N__22047),
            .lcout(),
            .ltout(\ALU.g0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_3_2_LC_2_9_4 .C_ON=1'b0;
    defparam \ALU.mult_g0_3_2_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_3_2_LC_2_9_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_3_2_LC_2_9_4  (
            .in0(N__20201),
            .in1(N__17663),
            .in2(N__16079),
            .in3(N__16076),
            .lcout(),
            .ltout(\ALU.g0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_LC_2_9_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_LC_2_9_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_g0_LC_2_9_5  (
            .in0(N__16070),
            .in1(N__16050),
            .in2(N__16064),
            .in3(N__17185),
            .lcout(\ALU.madd_350_0 ),
            .ltout(\ALU.madd_350_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m6_2_LC_2_9_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_m6_2_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m6_2_LC_2_9_6 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \ALU.mult_madd_m6_2_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__16145),
            .in2(N__16055),
            .in3(N__16052),
            .lcout(\ALU.madd_i3_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICJE9B_8_LC_2_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNICJE9B_8_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICJE9B_8_LC_2_9_7 .LUT_INIT=16'b1001010100101011;
    LogicCell40 \ALU.d_RNICJE9B_8_LC_2_9_7  (
            .in0(N__40043),
            .in1(N__20642),
            .in2(N__21470),
            .in3(N__47308),
            .lcout(\ALU.d_RNICJE9BZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIV4344_8_LC_2_10_0 .C_ON=1'b0;
    defparam \ALU.d_RNIV4344_8_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIV4344_8_LC_2_10_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \ALU.d_RNIV4344_8_LC_2_10_0  (
            .in0(N__24318),
            .in1(N__18655),
            .in2(_gnd_net_),
            .in3(N__18731),
            .lcout(\ALU.N_201_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m3_3_LC_2_10_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_m3_3_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m3_3_LC_2_10_1 .LUT_INIT=16'b0100000111010111;
    LogicCell40 \ALU.mult_madd_m3_3_LC_2_10_1  (
            .in0(N__16121),
            .in1(N__17214),
            .in2(N__17300),
            .in3(N__16185),
            .lcout(\ALU.madd_i1_mux_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_289_LC_2_10_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_289_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_289_LC_2_10_2 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_madd_289_LC_2_10_2  (
            .in0(N__17213),
            .in1(N__17295),
            .in2(N__16189),
            .in3(N__16120),
            .lcout(\ALU.madd_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIJ8B8_9_LC_2_10_3 .C_ON=1'b0;
    defparam \ALU.d_RNIIJ8B8_9_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIJ8B8_9_LC_2_10_3 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \ALU.d_RNIIJ8B8_9_LC_2_10_3  (
            .in0(N__20867),
            .in1(N__21096),
            .in2(N__26494),
            .in3(N__42011),
            .lcout(\ALU.a3_b_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_227_LC_2_10_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_227_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_227_LC_2_10_4 .LUT_INIT=16'b1111101011101000;
    LogicCell40 \ALU.mult_madd_227_LC_2_10_4  (
            .in0(N__19980),
            .in1(N__16103),
            .in2(N__16312),
            .in3(N__16231),
            .lcout(\ALU.madd_227 ),
            .ltout(\ALU.madd_227_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_285_LC_2_10_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_285_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_285_LC_2_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_285_LC_2_10_5  (
            .in0(N__17294),
            .in1(N__17212),
            .in2(N__16112),
            .in3(N__16181),
            .lcout(\ALU.madd_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_21_LC_2_11_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_21_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_21_LC_2_11_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \ALU.mult_g0_21_LC_2_11_0  (
            .in0(N__16241),
            .in1(_gnd_net_),
            .in2(N__37237),
            .in3(N__40086),
            .lcout(),
            .ltout(\ALU.madd_165_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_18_LC_2_11_1 .C_ON=1'b0;
    defparam \ALU.mult_g0_18_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_18_LC_2_11_1 .LUT_INIT=16'b1111111011001000;
    LogicCell40 \ALU.mult_g0_18_LC_2_11_1  (
            .in0(N__16102),
            .in1(N__19982),
            .in2(N__16109),
            .in3(N__16307),
            .lcout(\ALU.N_1533_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_170_0_tz_LC_2_11_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_170_0_tz_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_170_0_tz_LC_2_11_2 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \ALU.mult_madd_170_0_tz_LC_2_11_2  (
            .in0(N__39807),
            .in1(N__46686),
            .in2(N__37767),
            .in3(N__42662),
            .lcout(),
            .ltout(\ALU.madd_170_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_170_LC_2_11_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_170_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_170_LC_2_11_3 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \ALU.mult_madd_170_LC_2_11_3  (
            .in0(N__46963),
            .in1(N__41726),
            .in2(N__16106),
            .in3(N__23390),
            .lcout(\ALU.madd_170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_223_0_LC_2_11_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_223_0_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_223_0_LC_2_11_4 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \ALU.mult_madd_223_0_LC_2_11_4  (
            .in0(N__19981),
            .in1(N__16101),
            .in2(_gnd_net_),
            .in3(N__16232),
            .lcout(\ALU.madd_223_0 ),
            .ltout(\ALU.madd_223_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_238_0_LC_2_11_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_238_0_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_238_0_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_238_0_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__16324),
            .in2(N__16262),
            .in3(N__16308),
            .lcout(\ALU.madd_238_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_12_LC_2_11_6 .C_ON=1'b0;
    defparam \ALU.mult_g0_12_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_12_LC_2_11_6 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_g0_12_LC_2_11_6  (
            .in0(N__17299),
            .in1(N__17224),
            .in2(N__16190),
            .in3(N__16259),
            .lcout(\ALU.N_1559_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_165_0_LC_2_11_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_165_0_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_165_0_LC_2_11_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ALU.mult_madd_165_0_LC_2_11_7  (
            .in0(N__40085),
            .in1(N__37214),
            .in2(_gnd_net_),
            .in3(N__16240),
            .lcout(\ALU.madd_165_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_213_0_LC_2_12_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_213_0_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_213_0_LC_2_12_0 .LUT_INIT=16'b0101000010011100;
    LogicCell40 \ALU.mult_madd_213_0_LC_2_12_0  (
            .in0(N__46463),
            .in1(N__46693),
            .in2(N__40409),
            .in3(N__28027),
            .lcout(\ALU.madd_213_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIU9R47_5_LC_2_12_1 .C_ON=1'b0;
    defparam \ALU.d_RNIU9R47_5_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIU9R47_5_LC_2_12_1 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIU9R47_5_LC_2_12_1  (
            .in0(N__21766),
            .in1(N__40362),
            .in2(N__29967),
            .in3(N__21700),
            .lcout(\ALU.a5_b_5 ),
            .ltout(\ALU.a5_b_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_175_LC_2_12_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_175_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_175_LC_2_12_2 .LUT_INIT=16'b1111001000100000;
    LogicCell40 \ALU.mult_madd_175_LC_2_12_2  (
            .in0(N__41943),
            .in1(N__47088),
            .in2(N__16211),
            .in3(N__16207),
            .lcout(\ALU.madd_175 ),
            .ltout(\ALU.madd_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_232_LC_2_12_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_232_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_232_LC_2_12_3 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_madd_232_LC_2_12_3  (
            .in0(N__17554),
            .in1(N__16156),
            .in2(N__16193),
            .in3(N__16393),
            .lcout(\ALU.madd_232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI07LK7_4_LC_2_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNI07LK7_4_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI07LK7_4_LC_2_12_4 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNI07LK7_4_LC_2_12_4  (
            .in0(N__23486),
            .in1(N__46962),
            .in2(N__26576),
            .in3(N__23569),
            .lcout(\ALU.a7_b_4 ),
            .ltout(\ALU.a7_b_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_228_LC_2_12_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_228_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_228_LC_2_12_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_228_LC_2_12_5  (
            .in0(N__16163),
            .in1(N__16157),
            .in2(N__16148),
            .in3(N__16394),
            .lcout(\ALU.madd_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAMNM3_5_LC_2_12_6 .C_ON=1'b0;
    defparam \ALU.d_RNIAMNM3_5_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAMNM3_5_LC_2_12_6 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \ALU.d_RNIAMNM3_5_LC_2_12_6  (
            .in0(N__21699),
            .in1(N__21765),
            .in2(_gnd_net_),
            .in3(N__25229),
            .lcout(\ALU.N_225_0 ),
            .ltout(\ALU.N_225_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_64_0_LC_2_12_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_64_0_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_64_0_LC_2_12_7 .LUT_INIT=16'b0000101011000110;
    LogicCell40 \ALU.mult_madd_64_0_LC_2_12_7  (
            .in0(N__36962),
            .in1(N__41942),
            .in2(N__16385),
            .in3(N__42689),
            .lcout(\ALU.madd_64_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_290_0_LC_2_13_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_290_0_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_290_0_LC_2_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_290_0_LC_2_13_0  (
            .in0(N__18475),
            .in1(N__17648),
            .in2(_gnd_net_),
            .in3(N__16278),
            .lcout(),
            .ltout(\ALU.madd_290_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_299_LC_2_13_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_299_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_299_LC_2_13_1 .LUT_INIT=16'b1011111000101000;
    LogicCell40 \ALU.mult_madd_299_LC_2_13_1  (
            .in0(N__16496),
            .in1(N__16511),
            .in2(N__16382),
            .in3(N__16556),
            .lcout(\ALU.madd_299 ),
            .ltout(\ALU.madd_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_360_LC_2_13_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_360_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_360_LC_2_13_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_360_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16379),
            .in3(N__16368),
            .lcout(\ALU.madd_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_13_ma_LC_2_13_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_13_ma_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_13_ma_LC_2_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_madd_cry_13_ma_LC_2_13_3  (
            .in0(N__16369),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16345),
            .lcout(\ALU.madd_cry_13_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_242_LC_2_13_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_242_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_242_LC_2_13_4 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \ALU.mult_madd_242_LC_2_13_4  (
            .in0(N__16334),
            .in1(N__16325),
            .in2(N__16449),
            .in3(N__16313),
            .lcout(\ALU.madd_242 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_265_0_LC_2_13_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_265_0_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_265_0_LC_2_13_5 .LUT_INIT=16'b0000110010100110;
    LogicCell40 \ALU.mult_madd_265_0_LC_2_13_5  (
            .in0(N__40419),
            .in1(N__42933),
            .in2(N__21486),
            .in3(N__47087),
            .lcout(\ALU.madd_265_0 ),
            .ltout(\ALU.madd_265_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_280_LC_2_13_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_280_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_280_LC_2_13_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_280_LC_2_13_6  (
            .in0(N__17380),
            .in1(N__23775),
            .in2(N__16286),
            .in3(N__19919),
            .lcout(\ALU.madd_280 ),
            .ltout(\ALU.madd_280_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_295_0_LC_2_13_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_295_0_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_295_0_LC_2_13_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_295_0_LC_2_13_7  (
            .in0(N__17647),
            .in1(N__18474),
            .in2(N__16559),
            .in3(N__16555),
            .lcout(\ALU.madd_295_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_11_LC_2_14_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_11_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_11_LC_2_14_0 .LUT_INIT=16'b0111100001111000;
    LogicCell40 \ALU.mult_madd_axb_11_LC_2_14_0  (
            .in0(N__16544),
            .in1(N__16409),
            .in2(N__16475),
            .in3(_gnd_net_),
            .lcout(\ALU.madd_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI698B8_7_LC_2_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNI698B8_7_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI698B8_7_LC_2_14_1 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNI698B8_7_LC_2_14_1  (
            .in0(N__19849),
            .in1(N__42906),
            .in2(N__26496),
            .in3(N__19091),
            .lcout(\ALU.a4_b_7 ),
            .ltout(\ALU.a4_b_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_233_LC_2_14_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_233_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_233_LC_2_14_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_233_LC_2_14_2  (
            .in0(N__16688),
            .in1(N__17566),
            .in2(N__16517),
            .in3(N__16759),
            .lcout(\ALU.madd_233 ),
            .ltout(\ALU.madd_233_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_247_LC_2_14_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_247_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_247_LC_2_14_3 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \ALU.mult_madd_247_LC_2_14_3  (
            .in0(N__16604),
            .in1(N__16450),
            .in2(N__16514),
            .in3(N__16426),
            .lcout(\ALU.madd_247 ),
            .ltout(\ALU.madd_247_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_300_0_LC_2_14_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_300_0_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_300_0_LC_2_14_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_300_0_LC_2_14_4  (
            .in0(N__16510),
            .in1(N__16495),
            .in2(N__16484),
            .in3(N__16481),
            .lcout(\ALU.madd_N_10 ),
            .ltout(\ALU.madd_N_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_12_l_fx_LC_2_14_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_12_l_fx_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_12_l_fx_LC_2_14_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ALU.mult_madd_axb_12_l_fx_LC_2_14_5  (
            .in0(N__16466),
            .in1(N__25933),
            .in2(N__16460),
            .in3(N__16457),
            .lcout(\ALU.madd_axb_12_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_243_LC_2_14_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_243_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_243_LC_2_14_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_243_LC_2_14_6  (
            .in0(N__16451),
            .in1(N__16603),
            .in2(N__16430),
            .in3(N__16415),
            .lcout(\ALU.madd_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0B2B8_7_LC_2_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNI0B2B8_7_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0B2B8_7_LC_2_15_0 .LUT_INIT=16'b0101110010100011;
    LogicCell40 \ALU.d_RNI0B2B8_7_LC_2_15_0  (
            .in0(N__19838),
            .in1(N__19081),
            .in2(N__26495),
            .in3(N__46912),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITAM9D_7_LC_2_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNITAM9D_7_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITAM9D_7_LC_2_15_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNITAM9D_7_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16643),
            .in3(N__47049),
            .lcout(\ALU.d_RNITAM9DZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGF4I7_8_LC_2_15_2 .C_ON=1'b0;
    defparam \ALU.d_RNIGF4I7_8_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGF4I7_8_LC_2_15_2 .LUT_INIT=16'b0100111000000000;
    LogicCell40 \ALU.d_RNIGF4I7_8_LC_2_15_2  (
            .in0(N__24298),
            .in1(N__18730),
            .in2(N__18674),
            .in3(N__37985),
            .lcout(\ALU.a0_b_8 ),
            .ltout(\ALU.a0_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_103_LC_2_15_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_103_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_103_LC_2_15_3 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_103_LC_2_15_3  (
            .in0(N__17624),
            .in1(N__37503),
            .in2(N__16640),
            .in3(N__47050),
            .lcout(\ALU.madd_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITVJU4_7_LC_2_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNITVJU4_7_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITVJU4_7_LC_2_15_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \ALU.d_RNITVJU4_7_LC_2_15_4  (
            .in0(N__19837),
            .in1(N__24297),
            .in2(_gnd_net_),
            .in3(N__19080),
            .lcout(\ALU.N_213_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_148_LC_2_15_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_148_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_148_LC_2_15_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_148_LC_2_15_5  (
            .in0(N__16636),
            .in1(N__16792),
            .in2(_gnd_net_),
            .in3(N__16625),
            .lcout(\ALU.madd_148 ),
            .ltout(\ALU.madd_148_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_195_LC_2_15_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_195_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_195_LC_2_15_6 .LUT_INIT=16'b1110100011101000;
    LogicCell40 \ALU.mult_madd_195_LC_2_15_6  (
            .in0(N__16590),
            .in1(N__16572),
            .in2(N__16607),
            .in3(_gnd_net_),
            .lcout(\ALU.madd_247_0_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_143_LC_2_15_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_143_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_143_LC_2_15_7 .LUT_INIT=16'b1100111000001000;
    LogicCell40 \ALU.mult_madd_143_LC_2_15_7  (
            .in0(N__37986),
            .in1(N__22085),
            .in2(N__22073),
            .in3(N__21977),
            .lcout(\ALU.madd_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_181_LC_2_16_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_181_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_181_LC_2_16_0 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \ALU.mult_madd_181_LC_2_16_0  (
            .in0(N__16741),
            .in1(N__16702),
            .in2(N__16732),
            .in3(N__20329),
            .lcout(\ALU.madd_181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_129_LC_2_16_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_129_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_129_LC_2_16_1 .LUT_INIT=16'b0110100101100110;
    LogicCell40 \ALU.mult_madd_129_LC_2_16_1  (
            .in0(N__17717),
            .in1(N__16781),
            .in2(N__28088),
            .in3(N__42973),
            .lcout(\ALU.madd_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6I7F7_4_LC_2_16_2 .C_ON=1'b0;
    defparam \ALU.d_RNI6I7F7_4_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6I7F7_4_LC_2_16_2 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNI6I7F7_4_LC_2_16_2  (
            .in0(N__23501),
            .in1(N__40368),
            .in2(N__24283),
            .in3(N__23573),
            .lcout(\ALU.a5_b_4 ),
            .ltout(\ALU.a5_b_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_133_LC_2_16_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_133_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_133_LC_2_16_3 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_133_LC_2_16_3  (
            .in0(N__17716),
            .in1(N__42972),
            .in2(N__16775),
            .in3(N__28071),
            .lcout(\ALU.madd_133 ),
            .ltout(\ALU.madd_133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_185_LC_2_16_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_185_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_185_LC_2_16_4 .LUT_INIT=16'b1111101011101000;
    LogicCell40 \ALU.mult_madd_185_LC_2_16_4  (
            .in0(N__16725),
            .in1(N__16701),
            .in2(N__16772),
            .in3(N__20330),
            .lcout(\ALU.madd_237_0_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_23_LC_2_16_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_23_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_23_LC_2_16_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ALU.mult_g0_23_LC_2_16_5  (
            .in0(N__38318),
            .in1(N__39853),
            .in2(_gnd_net_),
            .in3(N__20375),
            .lcout(),
            .ltout(\ALU.madd_128_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_7_LC_2_16_6 .C_ON=1'b0;
    defparam \ALU.mult_g0_7_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_7_LC_2_16_6 .LUT_INIT=16'b1110111011101000;
    LogicCell40 \ALU.mult_g0_7_LC_2_16_6  (
            .in0(N__16742),
            .in1(N__16733),
            .in2(N__16706),
            .in3(N__16703),
            .lcout(),
            .ltout(\ALU.madd_237_0_tz_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_6_LC_2_16_7 .C_ON=1'b0;
    defparam \ALU.mult_g0_6_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_6_LC_2_16_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_g0_6_LC_2_16_7  (
            .in0(N__17675),
            .in1(_gnd_net_),
            .in2(N__16691),
            .in3(N__16687),
            .lcout(\ALU.N_1537_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m48_LC_3_1_0 .C_ON=1'b0;
    defparam \ALU.m48_LC_3_1_0 .SEQ_MODE=4'b0000;
    defparam \ALU.m48_LC_3_1_0 .LUT_INIT=16'b0110111101101000;
    LogicCell40 \ALU.m48_LC_3_1_0  (
            .in0(N__22698),
            .in1(N__22408),
            .in2(N__22600),
            .in3(N__48029),
            .lcout(),
            .ltout(\ALU.i6_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m50_LC_3_1_1 .C_ON=1'b0;
    defparam \ALU.m50_LC_3_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.m50_LC_3_1_1 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \ALU.m50_LC_3_1_1  (
            .in0(N__22324),
            .in1(N__22594),
            .in2(N__16646),
            .in3(N__22699),
            .lcout(),
            .ltout(N_51_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_0_LC_3_1_2 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_0_LC_3_1_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_0_LC_3_1_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CONTROL.aluOperation_0_LC_3_1_2  (
            .in0(N__33275),
            .in1(N__33434),
            .in2(N__16820),
            .in3(N__48030),
            .lcout(aluOperation_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47637),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m55_am_LC_3_1_4 .C_ON=1'b0;
    defparam \ALU.m55_am_LC_3_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m55_am_LC_3_1_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ALU.m55_am_LC_3_1_4  (
            .in0(N__22407),
            .in1(N__22322),
            .in2(N__22601),
            .in3(N__17771),
            .lcout(\ALU.m55_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m641_ns_1_LC_3_1_6 .C_ON=1'b0;
    defparam \ALU.m641_ns_1_LC_3_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m641_ns_1_LC_3_1_6 .LUT_INIT=16'b0111000001111111;
    LogicCell40 \ALU.m641_ns_1_LC_3_1_6  (
            .in0(N__22697),
            .in1(N__22323),
            .in2(N__33303),
            .in3(N__20483),
            .lcout(\ALU.m641_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m645_ns_1_LC_3_1_7 .C_ON=1'b0;
    defparam \ALU.m645_ns_1_LC_3_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m645_ns_1_LC_3_1_7 .LUT_INIT=16'b0010001000001111;
    LogicCell40 \ALU.m645_ns_1_LC_3_1_7  (
            .in0(N__22321),
            .in1(N__22696),
            .in2(N__43180),
            .in3(N__33271),
            .lcout(\ALU.m645_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_cnv_0_LC_3_2_0 .C_ON=1'b0;
    defparam \ALU.h_cnv_0_LC_3_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.h_cnv_0_LC_3_2_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.h_cnv_0_LC_3_2_0  (
            .in0(N__17924),
            .in1(N__20459),
            .in2(N__17888),
            .in3(N__17839),
            .lcout(\ALU.h_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.results_e_0_1_LC_3_2_1 .C_ON=1'b0;
    defparam \CONTROL.results_e_0_1_LC_3_2_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.results_e_0_1_LC_3_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.results_e_0_1_LC_3_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16952),
            .lcout(aluResults_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47643),
            .ce(N__16843),
            .sr(_gnd_net_));
    defparam \CONTROL.results_e_0_2_LC_3_2_2 .C_ON=1'b0;
    defparam \CONTROL.results_e_0_2_LC_3_2_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.results_e_0_2_LC_3_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.results_e_0_2_LC_3_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16817),
            .lcout(aluResults_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47643),
            .ce(N__16843),
            .sr(_gnd_net_));
    defparam \ALU.m16_LC_3_2_3 .C_ON=1'b0;
    defparam \ALU.m16_LC_3_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m16_LC_3_2_3 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \ALU.m16_LC_3_2_3  (
            .in0(N__22387),
            .in1(N__22276),
            .in2(N__22584),
            .in3(N__22676),
            .lcout(N_723),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m55_bm_LC_3_2_4 .C_ON=1'b0;
    defparam \ALU.m55_bm_LC_3_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m55_bm_LC_3_2_4 .LUT_INIT=16'b0000000000011111;
    LogicCell40 \ALU.m55_bm_LC_3_2_4  (
            .in0(N__22677),
            .in1(N__22388),
            .in2(N__22298),
            .in3(N__22555),
            .lcout(\ALU.m55_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m661_LC_3_2_5 .C_ON=1'b0;
    defparam \ALU.m661_LC_3_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.m661_LC_3_2_5 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \ALU.m661_LC_3_2_5  (
            .in0(N__22386),
            .in1(N__22275),
            .in2(N__22582),
            .in3(N__22675),
            .lcout(N_662_0),
            .ltout(N_662_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_cnv_0_LC_3_2_6 .C_ON=1'b0;
    defparam \CONTROL.operand1_cnv_0_LC_3_2_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.operand1_cnv_0_LC_3_2_6 .LUT_INIT=16'b1101000100000000;
    LogicCell40 \CONTROL.operand1_cnv_0_LC_3_2_6  (
            .in0(N__16889),
            .in1(N__33245),
            .in2(N__16892),
            .in3(N__34604),
            .lcout(\CONTROL.operand1_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m664_LC_3_2_7 .C_ON=1'b0;
    defparam \ALU.m664_LC_3_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m664_LC_3_2_7 .LUT_INIT=16'b0100100101011001;
    LogicCell40 \ALU.m664_LC_3_2_7  (
            .in0(N__22385),
            .in1(N__22274),
            .in2(N__22583),
            .in3(N__22674),
            .lcout(N_665_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m300_ns_LC_3_3_0 .C_ON=1'b0;
    defparam \ALU.m300_ns_LC_3_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.m300_ns_LC_3_3_0 .LUT_INIT=16'b1011010010111111;
    LogicCell40 \ALU.m300_ns_LC_3_3_0  (
            .in0(N__16877),
            .in1(N__22320),
            .in2(N__33302),
            .in3(N__44324),
            .lcout(),
            .ltout(N_301_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_3_LC_3_3_1 .C_ON=1'b0;
    defparam \CONTROL.aluParams_3_LC_3_3_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluParams_3_LC_3_3_1 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \CONTROL.aluParams_3_LC_3_3_1  (
            .in0(N__44325),
            .in1(_gnd_net_),
            .in2(N__16883),
            .in3(N__22124),
            .lcout(aluParams_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47649),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m667_LC_3_3_2 .C_ON=1'b0;
    defparam \ALU.m667_LC_3_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.m667_LC_3_3_2 .LUT_INIT=16'b0100100101011011;
    LogicCell40 \ALU.m667_LC_3_3_2  (
            .in0(N__22405),
            .in1(N__22319),
            .in2(N__22525),
            .in3(N__22685),
            .lcout(),
            .ltout(N_668_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_cnv_0_LC_3_3_3 .C_ON=1'b0;
    defparam \CONTROL.aluParams_cnv_0_LC_3_3_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluParams_cnv_0_LC_3_3_3 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \CONTROL.aluParams_cnv_0_LC_3_3_3  (
            .in0(N__34617),
            .in1(N__33264),
            .in2(N__16880),
            .in3(N__16863),
            .lcout(\CONTROL.aluParams_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m300_ns_1_LC_3_3_4 .C_ON=1'b0;
    defparam \ALU.m300_ns_1_LC_3_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m300_ns_1_LC_3_3_4 .LUT_INIT=16'b0001010111110101;
    LogicCell40 \ALU.m300_ns_1_LC_3_3_4  (
            .in0(N__22406),
            .in1(N__22686),
            .in2(N__33301),
            .in3(N__18065),
            .lcout(\ALU.m300_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m669_LC_3_3_5 .C_ON=1'b0;
    defparam \ALU.m669_LC_3_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.m669_LC_3_3_5 .LUT_INIT=16'b0011000111000001;
    LogicCell40 \ALU.m669_LC_3_3_5  (
            .in0(N__22684),
            .in1(N__22497),
            .in2(N__22325),
            .in3(N__22404),
            .lcout(),
            .ltout(N_670_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.results_cnv_0_LC_3_3_6 .C_ON=1'b0;
    defparam \CONTROL.results_cnv_0_LC_3_3_6 .SEQ_MODE=4'b0000;
    defparam \CONTROL.results_cnv_0_LC_3_3_6 .LUT_INIT=16'b1000101100000000;
    LogicCell40 \CONTROL.results_cnv_0_LC_3_3_6  (
            .in0(N__16864),
            .in1(N__33260),
            .in2(N__16850),
            .in3(N__34616),
            .lcout(\CONTROL.results_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1M3JE_14_LC_3_3_7 .C_ON=1'b0;
    defparam \ALU.d_RNI1M3JE_14_LC_3_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1M3JE_14_LC_3_3_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.d_RNI1M3JE_14_LC_3_3_7  (
            .in0(_gnd_net_),
            .in1(N__16901),
            .in2(_gnd_net_),
            .in3(N__21312),
            .lcout(\ALU.d_RNI1M3JEZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKNU29_14_LC_3_4_0 .C_ON=1'b0;
    defparam \ALU.d_RNIKNU29_14_LC_3_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKNU29_14_LC_3_4_0 .LUT_INIT=16'b0110011011000011;
    LogicCell40 \ALU.d_RNIKNU29_14_LC_3_4_0  (
            .in0(N__17811),
            .in1(N__40615),
            .in2(N__30646),
            .in3(N__26375),
            .lcout(\ALU.un2_addsub_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m636_LC_3_4_1 .C_ON=1'b0;
    defparam \ALU.m636_LC_3_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.m636_LC_3_4_1 .LUT_INIT=16'b0000011100001100;
    LogicCell40 \ALU.m636_LC_3_4_1  (
            .in0(N__22715),
            .in1(N__22419),
            .in2(N__22526),
            .in3(N__22285),
            .lcout(\ALU.N_724 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5SME5_14_LC_3_4_2 .C_ON=1'b0;
    defparam \ALU.d_RNI5SME5_14_LC_3_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5SME5_14_LC_3_4_2 .LUT_INIT=16'b0111010001110100;
    LogicCell40 \ALU.d_RNI5SME5_14_LC_3_4_2  (
            .in0(N__17812),
            .in1(N__26380),
            .in2(N__30647),
            .in3(_gnd_net_),
            .lcout(\ALU.N_171_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9G6T4_9_LC_3_4_4 .C_ON=1'b0;
    defparam \ALU.d_RNI9G6T4_9_LC_3_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9G6T4_9_LC_3_4_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ALU.d_RNI9G6T4_9_LC_3_4_4  (
            .in0(N__20870),
            .in1(N__26379),
            .in2(_gnd_net_),
            .in3(N__21094),
            .lcout(\ALU.N_207_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILOIL8_9_LC_3_4_5 .C_ON=1'b0;
    defparam \ALU.d_RNILOIL8_9_LC_3_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILOIL8_9_LC_3_4_5 .LUT_INIT=16'b0101110010100011;
    LogicCell40 \ALU.d_RNILOIL8_9_LC_3_4_5  (
            .in0(N__21093),
            .in1(N__20869),
            .in2(N__26445),
            .in3(N__39847),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6B7KD_9_LC_3_4_6 .C_ON=1'b0;
    defparam \ALU.d_RNI6B7KD_9_LC_3_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6B7KD_9_LC_3_4_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNI6B7KD_9_LC_3_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16895),
            .in3(N__22065),
            .lcout(\ALU.d_RNI6B7KDZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIF9794_9_LC_3_4_7 .C_ON=1'b0;
    defparam \ALU.d_RNIF9794_9_LC_3_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIF9794_9_LC_3_4_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \ALU.d_RNIF9794_9_LC_3_4_7  (
            .in0(N__21095),
            .in1(N__29405),
            .in2(_gnd_net_),
            .in3(N__39848),
            .lcout(\ALU.N_274_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m252_LC_3_5_0 .C_ON=1'b0;
    defparam \ALU.m252_LC_3_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.m252_LC_3_5_0 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \ALU.m252_LC_3_5_0  (
            .in0(N__19630),
            .in1(N__19651),
            .in2(_gnd_net_),
            .in3(N__21563),
            .lcout(\ALU.N_253_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_362_LC_3_5_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_362_LC_3_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_362_LC_3_5_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \ALU.mult_madd_362_LC_3_5_1  (
            .in0(N__40599),
            .in1(N__18835),
            .in2(N__38337),
            .in3(N__18151),
            .lcout(\ALU.madd_362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_366_LC_3_5_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_366_LC_3_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_366_LC_3_5_2 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_366_LC_3_5_2  (
            .in0(N__18836),
            .in1(N__38322),
            .in2(N__18155),
            .in3(N__40600),
            .lcout(\ALU.madd_366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_0_ma_LC_3_5_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_0_ma_LC_3_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_0_ma_LC_3_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_madd_cry_0_ma_LC_3_5_3  (
            .in0(N__38323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37471),
            .lcout(\ALU.madd_cry_0_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIH1R53_1_LC_3_5_4 .C_ON=1'b0;
    defparam \ALU.d_RNIH1R53_1_LC_3_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIH1R53_1_LC_3_5_4 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \ALU.d_RNIH1R53_1_LC_3_5_4  (
            .in0(N__37472),
            .in1(_gnd_net_),
            .in2(N__29434),
            .in3(N__23342),
            .lcout(\ALU.N_292_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI21MU3_6_LC_3_5_5 .C_ON=1'b0;
    defparam \ALU.d_RNI21MU3_6_LC_3_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI21MU3_6_LC_3_5_5 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \ALU.d_RNI21MU3_6_LC_3_5_5  (
            .in0(N__26283),
            .in1(N__29413),
            .in2(_gnd_net_),
            .in3(N__46670),
            .lcout(\ALU.N_291_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICCNU3_7_LC_3_5_6 .C_ON=1'b0;
    defparam \ALU.d_RNICCNU3_7_LC_3_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICCNU3_7_LC_3_5_6 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \ALU.d_RNICCNU3_7_LC_3_5_6  (
            .in0(N__46966),
            .in1(_gnd_net_),
            .in2(N__29433),
            .in3(N__19822),
            .lcout(\ALU.N_264_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAB477_6_LC_3_5_7 .C_ON=1'b0;
    defparam \ALU.d_RNIAB477_6_LC_3_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAB477_6_LC_3_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNIAB477_6_LC_3_5_7  (
            .in0(N__43688),
            .in1(N__46965),
            .in2(_gnd_net_),
            .in3(N__46669),
            .lcout(\ALU.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIGTNC7_13_LC_3_6_0 .C_ON=1'b0;
    defparam \ALU.c_RNIGTNC7_13_LC_3_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIGTNC7_13_LC_3_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.c_RNIGTNC7_13_LC_3_6_0  (
            .in0(_gnd_net_),
            .in1(N__40763),
            .in2(_gnd_net_),
            .in3(N__37759),
            .lcout(\ALU.a13_b_1 ),
            .ltout(\ALU.a13_b_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_376_LC_3_6_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_376_LC_3_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_376_LC_3_6_1 .LUT_INIT=16'b1011001010100000;
    LogicCell40 \ALU.mult_madd_376_LC_3_6_1  (
            .in0(N__17006),
            .in1(N__21296),
            .in2(N__16904),
            .in3(N__38026),
            .lcout(\ALU.madd_376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDU4G5_14_LC_3_6_2 .C_ON=1'b0;
    defparam \ALU.d_RNIDU4G5_14_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDU4G5_14_LC_3_6_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \ALU.d_RNIDU4G5_14_LC_3_6_2  (
            .in0(N__17802),
            .in1(N__24234),
            .in2(_gnd_net_),
            .in3(N__30634),
            .lcout(\ALU.N_171_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m168_LC_3_6_3 .C_ON=1'b0;
    defparam \ALU.m168_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m168_LC_3_6_3 .LUT_INIT=16'b1110111001111111;
    LogicCell40 \ALU.m168_LC_3_6_3  (
            .in0(N__30201),
            .in1(N__25205),
            .in2(N__16997),
            .in3(N__29740),
            .lcout(\ALU.N_169_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIDMS7_3_LC_3_6_4 .C_ON=1'b0;
    defparam \ALU.d_RNIIDMS7_3_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIDMS7_3_LC_3_6_4 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIIDMS7_3_LC_3_6_4  (
            .in0(N__23920),
            .in1(N__39375),
            .in2(N__29914),
            .in3(N__24029),
            .lcout(\ALU.a11_b_3 ),
            .ltout(\ALU.a11_b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_372_LC_3_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_372_LC_3_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_372_LC_3_6_5 .LUT_INIT=16'b0110100101011010;
    LogicCell40 \ALU.mult_madd_372_LC_3_6_5  (
            .in0(N__17155),
            .in1(N__21297),
            .in2(N__17000),
            .in3(N__38027),
            .lcout(\ALU.madd_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_30_LC_3_6_6.C_ON=1'b0;
    defparam testWord_30_LC_3_6_6.SEQ_MODE=4'b1000;
    defparam testWord_30_LC_3_6_6.LUT_INIT=16'b1110110001001100;
    LogicCell40 testWord_30_LC_3_6_6 (
            .in0(N__41219),
            .in1(N__16996),
            .in2(N__41477),
            .in3(N__16981),
            .lcout(ctrlOut_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__41056),
            .sr(_gnd_net_));
    defparam testWord_14_LC_3_6_7.C_ON=1'b0;
    defparam testWord_14_LC_3_6_7.SEQ_MODE=4'b1000;
    defparam testWord_14_LC_3_6_7.LUT_INIT=16'b1110001011110000;
    LogicCell40 testWord_14_LC_3_6_7 (
            .in0(N__16980),
            .in1(N__41438),
            .in2(N__16948),
            .in3(N__41218),
            .lcout(testWordZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__41056),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI05GC8_7_LC_3_7_0 .C_ON=1'b0;
    defparam \ALU.d_RNI05GC8_7_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI05GC8_7_LC_3_7_0 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNI05GC8_7_LC_3_7_0  (
            .in0(N__19842),
            .in1(N__19102),
            .in2(N__30012),
            .in3(N__46728),
            .lcout(\ALU.a6_b_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN9HA7_6_LC_3_7_1 .C_ON=1'b0;
    defparam \ALU.d_RNIN9HA7_6_LC_3_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN9HA7_6_LC_3_7_1 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \ALU.d_RNIN9HA7_6_LC_3_7_1  (
            .in0(N__26732),
            .in1(N__26276),
            .in2(N__29956),
            .in3(N__46943),
            .lcout(\ALU.a7_b_6 ),
            .ltout(\ALU.a7_b_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_320_LC_3_7_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_320_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_320_LC_3_7_2 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \ALU.mult_madd_320_LC_3_7_2  (
            .in0(N__16928),
            .in1(N__40082),
            .in2(N__16931),
            .in3(N__28085),
            .lcout(\ALU.madd_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_392_LC_3_7_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_392_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_392_LC_3_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_392_LC_3_7_3  (
            .in0(N__16910),
            .in1(N__19733),
            .in2(_gnd_net_),
            .in3(N__18317),
            .lcout(\ALU.madd_392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_324_LC_3_7_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_324_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_324_LC_3_7_4 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_324_LC_3_7_4  (
            .in0(N__16927),
            .in1(N__40083),
            .in2(N__16919),
            .in3(N__28086),
            .lcout(\ALU.madd_324_0 ),
            .ltout(\ALU.madd_324_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_396_LC_3_7_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_396_LC_3_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_396_LC_3_7_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_396_LC_3_7_5  (
            .in0(_gnd_net_),
            .in1(N__19732),
            .in2(N__17069),
            .in3(N__18316),
            .lcout(\ALU.madd_396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGS0L7_6_LC_3_7_6 .C_ON=1'b0;
    defparam \ALU.d_RNIGS0L7_6_LC_3_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGS0L7_6_LC_3_7_6 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIGS0L7_6_LC_3_7_6  (
            .in0(N__26277),
            .in1(N__40081),
            .in2(N__30013),
            .in3(N__26731),
            .lcout(\ALU.a8_b_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_372_0_LC_3_7_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_372_0_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_372_0_LC_3_7_7 .LUT_INIT=16'b0100010010110100;
    LogicCell40 \ALU.mult_madd_372_0_LC_3_7_7  (
            .in0(N__21311),
            .in1(N__38035),
            .in2(N__39396),
            .in3(N__41736),
            .lcout(\ALU.madd_372_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_21_LC_3_8_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_21_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_21_LC_3_8_0 .LUT_INIT=16'b0001011111101000;
    LogicCell40 \ALU.mult_madd_484_21_LC_3_8_0  (
            .in0(N__17066),
            .in1(N__17171),
            .in2(N__17015),
            .in3(N__17057),
            .lcout(\ALU.madd_484_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1S6M7_5_LC_3_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNI1S6M7_5_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1S6M7_5_LC_3_8_1 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNI1S6M7_5_LC_3_8_1  (
            .in0(N__21785),
            .in1(N__39808),
            .in2(N__30022),
            .in3(N__21721),
            .lcout(\ALU.a9_b_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_411_LC_3_8_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_411_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_411_LC_3_8_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_411_LC_3_8_2  (
            .in0(N__17125),
            .in1(N__17144),
            .in2(_gnd_net_),
            .in3(N__17137),
            .lcout(),
            .ltout(\ALU.madd_411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_24_LC_3_8_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_24_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_24_LC_3_8_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_484_24_LC_3_8_3  (
            .in0(N__17051),
            .in1(N__17114),
            .in2(N__17045),
            .in3(N__18275),
            .lcout(\ALU.madd_484_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_381_LC_3_8_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_381_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_381_LC_3_8_4 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_381_LC_3_8_4  (
            .in0(N__17023),
            .in1(N__27554),
            .in2(N__17036),
            .in3(N__42675),
            .lcout(\ALU.madd_381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_377_LC_3_8_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_377_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_377_LC_3_8_5 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \ALU.mult_madd_377_LC_3_8_5  (
            .in0(N__42676),
            .in1(N__17035),
            .in2(N__27594),
            .in3(N__17024),
            .lcout(\ALU.madd_377 ),
            .ltout(\ALU.madd_377_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_397_LC_3_8_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_397_LC_3_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_397_LC_3_8_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_397_LC_3_8_6  (
            .in0(N__17177),
            .in1(N__17170),
            .in2(N__17162),
            .in3(N__17159),
            .lcout(\ALU.madd_397 ),
            .ltout(\ALU.madd_397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_407_LC_3_8_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_407_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_407_LC_3_8_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_407_LC_3_8_7  (
            .in0(N__17138),
            .in1(_gnd_net_),
            .in2(N__17129),
            .in3(N__17126),
            .lcout(\ALU.madd_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_406_LC_3_9_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_406_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_406_LC_3_9_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_406_LC_3_9_0  (
            .in0(N__17105),
            .in1(N__18344),
            .in2(_gnd_net_),
            .in3(N__17098),
            .lcout(\ALU.madd_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0PL97_8_LC_3_9_1 .C_ON=1'b0;
    defparam \ALU.d_RNI0PL97_8_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0PL97_8_LC_3_9_1 .LUT_INIT=16'b0010111000000000;
    LogicCell40 \ALU.d_RNI0PL97_8_LC_3_9_1  (
            .in0(N__18738),
            .in1(N__26514),
            .in2(N__18669),
            .in3(N__40430),
            .lcout(),
            .ltout(\ALU.a5_b_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_329_LC_3_9_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_329_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_329_LC_3_9_2 .LUT_INIT=16'b1111001000100000;
    LogicCell40 \ALU.mult_madd_329_LC_3_9_2  (
            .in0(N__42927),
            .in1(N__22064),
            .in2(N__17108),
            .in3(N__17431),
            .lcout(\ALU.madd_329_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_387_LC_3_9_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_387_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_387_LC_3_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_387_LC_3_9_3  (
            .in0(N__18358),
            .in1(N__18241),
            .in2(_gnd_net_),
            .in3(N__18265),
            .lcout(\ALU.madd_387 ),
            .ltout(\ALU.madd_387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_402_LC_3_9_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_402_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_402_LC_3_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_402_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(N__17099),
            .in2(N__17090),
            .in3(N__18343),
            .lcout(\ALU.madd_402 ),
            .ltout(\ALU.madd_402_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_412_LC_3_9_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_412_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_412_LC_3_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_412_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__18430),
            .in2(N__17081),
            .in3(N__17407),
            .lcout(\ALU.madd_412 ),
            .ltout(\ALU.madd_412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_417_LC_3_9_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_417_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_417_LC_3_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_417_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__17078),
            .in2(N__17072),
            .in3(N__17344),
            .lcout(\ALU.madd_329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_573_LC_3_9_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_573_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_573_LC_3_9_7 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \ALU.mult_madd_573_LC_3_9_7  (
            .in0(N__17345),
            .in1(N__17336),
            .in2(_gnd_net_),
            .in3(N__17330),
            .lcout(\ALU.madd_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_9_LC_3_10_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_9_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_9_LC_3_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_g0_9_LC_3_10_0  (
            .in0(N__38329),
            .in1(N__25372),
            .in2(N__37000),
            .in3(N__39594),
            .lcout(\ALU.madd_141_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_270_0_LC_3_10_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_270_0_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_270_0_LC_3_10_1 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_270_0_LC_3_10_1  (
            .in0(N__25373),
            .in1(N__17279),
            .in2(N__17252),
            .in3(N__38330),
            .lcout(\ALU.madd_270_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_0_rep1_LC_3_10_2 .C_ON=1'b0;
    defparam \CONTROL.operand2_0_rep1_LC_3_10_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_0_rep1_LC_3_10_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \CONTROL.operand2_0_rep1_LC_3_10_2  (
            .in0(N__34681),
            .in1(N__34798),
            .in2(N__31250),
            .in3(N__41112),
            .lcout(aluOperand2_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47686),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_207_LC_3_10_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_207_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_207_LC_3_10_3 .LUT_INIT=16'b1110110010000000;
    LogicCell40 \ALU.mult_madd_207_LC_3_10_3  (
            .in0(N__39394),
            .in1(N__19997),
            .in2(N__38339),
            .in3(N__19961),
            .lcout(\ALU.madd_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_250_0_LC_3_10_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_250_0_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_250_0_LC_3_10_4 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_250_0_LC_3_10_4  (
            .in0(N__27539),
            .in1(N__39593),
            .in2(N__36999),
            .in3(N__37232),
            .lcout(\ALU.madd_250_0 ),
            .ltout(\ALU.madd_250_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_250_LC_3_10_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_250_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_250_LC_3_10_5 .LUT_INIT=16'b0011110011110000;
    LogicCell40 \ALU.mult_madd_250_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(N__25354),
            .in2(N__17273),
            .in3(N__38331),
            .lcout(\ALU.madd_250 ),
            .ltout(\ALU.madd_250_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_274_LC_3_10_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_274_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_274_LC_3_10_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_274_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(N__17250),
            .in2(N__17228),
            .in3(N__17211),
            .lcout(\ALU.madd_274 ),
            .ltout(\ALU.madd_274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_344_LC_3_10_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_344_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_344_LC_3_10_7 .LUT_INIT=16'b1011001011101000;
    LogicCell40 \ALU.mult_madd_344_LC_3_10_7  (
            .in0(N__17490),
            .in1(N__17456),
            .in2(N__17438),
            .in3(N__17435),
            .lcout(\ALU.madd_344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_25_LC_3_11_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_25_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_25_LC_3_11_0 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \ALU.mult_madd_25_LC_3_11_0  (
            .in0(N__23617),
            .in1(N__38029),
            .in2(N__24065),
            .in3(N__28026),
            .lcout(\ALU.madd_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_29_LC_3_11_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_29_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_29_LC_3_11_1 .LUT_INIT=16'b1101110001000000;
    LogicCell40 \ALU.mult_madd_29_LC_3_11_1  (
            .in0(N__28025),
            .in1(N__24064),
            .in2(N__38046),
            .in3(N__23618),
            .lcout(\ALU.madd_29 ),
            .ltout(\ALU.madd_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_47_LC_3_11_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_47_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_47_LC_3_11_2 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \ALU.mult_madd_47_LC_3_11_2  (
            .in0(N__18905),
            .in1(N__38033),
            .in2(N__17396),
            .in3(N__46473),
            .lcout(\ALU.madd_47 ),
            .ltout(\ALU.madd_47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_5_l_fx_LC_3_11_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_5_l_fx_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_5_l_fx_LC_3_11_3 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ALU.mult_madd_axb_5_l_fx_LC_3_11_3  (
            .in0(N__18782),
            .in1(N__26183),
            .in2(N__17393),
            .in3(N__18791),
            .lcout(\ALU.madd_axb_5_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_4_l_fx_LC_3_11_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_4_l_fx_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_4_l_fx_LC_3_11_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.mult_madd_axb_4_l_fx_LC_3_11_4  (
            .in0(N__18790),
            .in1(N__25741),
            .in2(_gnd_net_),
            .in3(N__18781),
            .lcout(\ALU.madd_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_284_LC_3_11_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_284_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_284_LC_3_11_5 .LUT_INIT=16'b1111011001100000;
    LogicCell40 \ALU.mult_madd_284_LC_3_11_5  (
            .in0(N__17390),
            .in1(N__23779),
            .in2(N__17381),
            .in3(N__19915),
            .lcout(\ALU.madd_284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_309_LC_3_11_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_309_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_309_LC_3_11_6 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_madd_309_LC_3_11_6  (
            .in0(N__37205),
            .in1(N__39322),
            .in2(N__35069),
            .in3(N__18818),
            .lcout(\ALU.madd_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGGQ26_1_LC_3_11_7 .C_ON=1'b0;
    defparam \ALU.d_RNIGGQ26_1_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGGQ26_1_LC_3_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIGGQ26_1_LC_3_11_7  (
            .in0(N__37485),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37204),
            .lcout(\ALU.a1_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIG1A7_6_LC_3_12_0 .C_ON=1'b0;
    defparam \ALU.d_RNIIG1A7_6_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIG1A7_6_LC_3_12_0 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIIG1A7_6_LC_3_12_0  (
            .in0(N__26284),
            .in1(N__36958),
            .in2(N__30054),
            .in3(N__26729),
            .lcout(\ALU.a2_b_6 ),
            .ltout(\ALU.a2_b_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_99_LC_3_12_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_99_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_99_LC_3_12_1 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \ALU.mult_madd_99_LC_3_12_1  (
            .in0(N__37486),
            .in1(N__17612),
            .in2(N__17600),
            .in3(N__47096),
            .lcout(\ALU.madd_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILIL37_6_LC_3_12_2 .C_ON=1'b0;
    defparam \ALU.d_RNILIL37_6_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILIL37_6_LC_3_12_2 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNILIL37_6_LC_3_12_2  (
            .in0(N__26285),
            .in1(N__40410),
            .in2(N__30055),
            .in3(N__26730),
            .lcout(\ALU.a5_b_6 ),
            .ltout(\ALU.a5_b_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_217_LC_3_12_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_217_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_217_LC_3_12_3 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_217_LC_3_12_3  (
            .in0(N__17532),
            .in1(N__46961),
            .in2(N__17597),
            .in3(N__42666),
            .lcout(\ALU.madd_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_42_0_LC_3_12_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_42_0_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_42_0_LC_3_12_5 .LUT_INIT=16'b0010001011010010;
    LogicCell40 \ALU.mult_madd_42_0_LC_3_12_5  (
            .in0(N__37487),
            .in1(N__28034),
            .in2(N__36998),
            .in3(N__42667),
            .lcout(\ALU.madd_42_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN9H73_5_LC_3_12_6 .C_ON=1'b0;
    defparam \ALU.d_RNIN9H73_5_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN9H73_5_LC_3_12_6 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.d_RNIN9H73_5_LC_3_12_6  (
            .in0(N__28541),
            .in1(N__31655),
            .in2(N__33096),
            .in3(N__28883),
            .lcout(\ALU.operand2_5 ),
            .ltout(\ALU.operand2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINMLB7_5_LC_3_12_7 .C_ON=1'b0;
    defparam \ALU.d_RNINMLB7_5_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINMLB7_5_LC_3_12_7 .LUT_INIT=16'b0010000010101000;
    LogicCell40 \ALU.d_RNINMLB7_5_LC_3_12_7  (
            .in0(N__46672),
            .in1(N__30032),
            .in2(N__17594),
            .in3(N__21784),
            .lcout(\ALU.a6_b_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_176_0_LC_3_13_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_176_0_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_176_0_LC_3_13_0 .LUT_INIT=16'b0000101011000110;
    LogicCell40 \ALU.mult_madd_176_0_LC_3_13_0  (
            .in0(N__36964),
            .in1(N__37488),
            .in2(N__21485),
            .in3(N__22066),
            .lcout(\ALU.madd_176_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_218_0_LC_3_13_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_218_0_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_218_0_LC_3_13_1 .LUT_INIT=16'b0100101101000100;
    LogicCell40 \ALU.mult_madd_218_0_LC_3_13_1  (
            .in0(N__22067),
            .in1(N__36966),
            .in2(N__21487),
            .in3(N__41927),
            .lcout(\ALU.madd_218_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_275_0_LC_3_13_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_275_0_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_275_0_LC_3_13_2 .LUT_INIT=16'b0001011111101000;
    LogicCell40 \ALU.mult_madd_275_0_LC_3_13_2  (
            .in0(N__17555),
            .in1(N__17533),
            .in2(N__17509),
            .in3(N__18525),
            .lcout(\ALU.madd_275_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_42_LC_3_13_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_42_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_42_LC_3_13_3 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \ALU.mult_madd_42_LC_3_13_3  (
            .in0(N__37489),
            .in1(N__23605),
            .in2(N__24376),
            .in3(N__28035),
            .lcout(\ALU.madd_42 ),
            .ltout(\ALU.madd_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m3_2_LC_3_13_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_m3_2_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m3_2_LC_3_13_4 .LUT_INIT=16'b0000001100111111;
    LogicCell40 \ALU.mult_madd_m3_2_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(N__19003),
            .in2(N__17639),
            .in3(N__19022),
            .lcout(\ALU.madd_i1_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_52_0_LC_3_13_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_52_0_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_52_0_LC_3_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_52_0_LC_3_13_5  (
            .in0(N__19004),
            .in1(_gnd_net_),
            .in2(N__24377),
            .in3(N__17636),
            .lcout(\ALU.madd_52_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_1_ma_LC_3_13_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_1_ma_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_1_ma_LC_3_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_madd_cry_1_ma_LC_3_13_6  (
            .in0(N__37703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37490),
            .lcout(\ALU.madd_cry_1_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVQ5R6_2_LC_3_13_7 .C_ON=1'b0;
    defparam \ALU.d_RNIVQ5R6_2_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVQ5R6_2_LC_3_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIVQ5R6_2_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(N__36965),
            .in2(_gnd_net_),
            .in3(N__37702),
            .lcout(\ALU.a2_b_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFDNC8_7_LC_3_14_0 .C_ON=1'b0;
    defparam \ALU.d_RNIFDNC8_7_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFDNC8_7_LC_3_14_0 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIFDNC8_7_LC_3_14_0  (
            .in0(N__19819),
            .in1(N__42905),
            .in2(N__30056),
            .in3(N__19085),
            .lcout(\ALU.a4_b_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIM09H_7_LC_3_14_1 .C_ON=1'b0;
    defparam \ALU.e_RNIM09H_7_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIM09H_7_LC_3_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.e_RNIM09H_7_LC_3_14_1  (
            .in0(N__27875),
            .in1(N__28805),
            .in2(_gnd_net_),
            .in3(N__32079),
            .lcout(),
            .ltout(\ALU.e_RNIM09HZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIKJH32_7_LC_3_14_2 .C_ON=1'b0;
    defparam \ALU.e_RNIKJH32_7_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIKJH32_7_LC_3_14_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.e_RNIKJH32_7_LC_3_14_2  (
            .in0(N__33085),
            .in1(N__34512),
            .in2(N__17630),
            .in3(N__31670),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIULB84_7_LC_3_14_3 .C_ON=1'b0;
    defparam \ALU.d_RNIULB84_7_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIULB84_7_LC_3_14_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIULB84_7_LC_3_14_3  (
            .in0(N__32963),
            .in1(N__45203),
            .in2(N__17627),
            .in3(N__26897),
            .lcout(\ALU.operand2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g1_2_LC_3_14_4 .C_ON=1'b0;
    defparam \ALU.mult_g1_2_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g1_2_LC_3_14_4 .LUT_INIT=16'b1010001111111111;
    LogicCell40 \ALU.mult_g1_2_LC_3_14_4  (
            .in0(N__18673),
            .in1(N__18740),
            .in2(N__30057),
            .in3(N__41919),
            .lcout(),
            .ltout(\ALU.g1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_25_LC_3_14_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_25_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_25_LC_3_14_5 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \ALU.mult_g0_25_LC_3_14_5  (
            .in0(N__22072),
            .in1(N__36963),
            .in2(N__17684),
            .in3(N__17681),
            .lcout(\ALU.g2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIL5C37_5_LC_3_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNIL5C37_5_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIL5C37_5_LC_3_15_0 .LUT_INIT=16'b0101110010100011;
    LogicCell40 \ALU.d_RNIL5C37_5_LC_3_15_0  (
            .in0(N__21786),
            .in1(N__21722),
            .in2(N__26603),
            .in3(N__40367),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVR3QA_5_LC_3_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIVR3QA_5_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVR3QA_5_LC_3_15_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNIVR3QA_5_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17666),
            .in3(N__28070),
            .lcout(\ALU.d_RNIVR3QAZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICFBS3_5_LC_3_15_2 .C_ON=1'b0;
    defparam \ALU.d_RNICFBS3_5_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICFBS3_5_LC_3_15_2 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \ALU.d_RNICFBS3_5_LC_3_15_2  (
            .in0(N__21787),
            .in1(N__21723),
            .in2(_gnd_net_),
            .in3(N__26575),
            .lcout(\ALU.N_225_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILT5T4_7_LC_3_15_3 .C_ON=1'b0;
    defparam \ALU.d_RNILT5T4_7_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILT5T4_7_LC_3_15_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ALU.d_RNILT5T4_7_LC_3_15_3  (
            .in0(N__19089),
            .in1(N__26564),
            .in2(_gnd_net_),
            .in3(N__19821),
            .lcout(\ALU.N_213_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN01B8_7_LC_3_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNIN01B8_7_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN01B8_7_LC_3_15_4 .LUT_INIT=16'b0010101000100000;
    LogicCell40 \ALU.d_RNIN01B8_7_LC_3_15_4  (
            .in0(N__46616),
            .in1(N__19820),
            .in2(N__26604),
            .in3(N__19090),
            .lcout(\ALU.a6_b_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNII0KR6_6_LC_3_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNII0KR6_6_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNII0KR6_6_LC_3_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNII0KR6_6_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__46615),
            .in2(_gnd_net_),
            .in3(N__38291),
            .lcout(\ALU.a6_b_0 ),
            .ltout(\ALU.a6_b_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_41_LC_3_15_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_41_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_41_LC_3_15_6 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_41_LC_3_15_6  (
            .in0(N__18863),
            .in1(N__40366),
            .in2(N__17651),
            .in3(N__37730),
            .lcout(\ALU.madd_41 ),
            .ltout(\ALU.madd_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_69_LC_3_15_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_69_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_69_LC_3_15_7 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \ALU.mult_madd_69_LC_3_15_7  (
            .in0(N__19036),
            .in1(N__37514),
            .in2(N__17726),
            .in3(N__46448),
            .lcout(\ALU.madd_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_46_LC_3_16_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_46_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_46_LC_3_16_0 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_46_LC_3_16_0  (
            .in0(N__23606),
            .in1(N__37513),
            .in2(N__24375),
            .in3(N__28087),
            .lcout(\ALU.madd_46 ),
            .ltout(\ALU.madd_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_76_LC_3_16_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_76_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_76_LC_3_16_1 .LUT_INIT=16'b1011000001000000;
    LogicCell40 \ALU.mult_madd_76_LC_3_16_1  (
            .in0(N__41721),
            .in1(N__42995),
            .in2(N__17723),
            .in3(N__18940),
            .lcout(\ALU.madd_39 ),
            .ltout(\ALU.madd_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_118_LC_3_16_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_118_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_118_LC_3_16_2 .LUT_INIT=16'b1111111010101000;
    LogicCell40 \ALU.mult_madd_118_LC_3_16_2  (
            .in0(N__20366),
            .in1(N__17702),
            .in2(N__17720),
            .in3(N__19226),
            .lcout(\ALU.madd_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDAJB7_3_LC_3_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNIDAJB7_3_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDAJB7_3_LC_3_16_3 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNIDAJB7_3_LC_3_16_3  (
            .in0(N__23945),
            .in1(N__24030),
            .in2(N__24317),
            .in3(N__46671),
            .lcout(\ALU.a6_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_78_0_tz_LC_3_16_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_78_0_tz_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_78_0_tz_LC_3_16_4 .LUT_INIT=16'b1111101011110110;
    LogicCell40 \ALU.mult_madd_78_0_tz_LC_3_16_4  (
            .in0(N__18939),
            .in1(N__42994),
            .in2(N__19217),
            .in3(N__41720),
            .lcout(),
            .ltout(\ALU.madd_78_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_78_0_LC_3_16_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_78_0_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_78_0_LC_3_16_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.mult_madd_78_0_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17705),
            .in3(N__20414),
            .lcout(\ALU.madd_78_0 ),
            .ltout(\ALU.madd_78_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_114_LC_3_16_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_114_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_114_LC_3_16_6 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \ALU.mult_madd_114_LC_3_16_6  (
            .in0(N__20365),
            .in1(N__17696),
            .in2(N__17690),
            .in3(N__19225),
            .lcout(\ALU.madd_114 ),
            .ltout(\ALU.madd_114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_8_l_fx_LC_3_16_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_8_l_fx_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_8_l_fx_LC_3_16_7 .LUT_INIT=16'b1100000011111100;
    LogicCell40 \ALU.mult_madd_axb_8_l_fx_LC_3_16_7  (
            .in0(N__26068),
            .in1(N__19307),
            .in2(N__17687),
            .in3(N__18872),
            .lcout(\ALU.madd_axb_8_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testClock_RNIAQVB_LC_4_1_1.C_ON=1'b0;
    defparam testClock_RNIAQVB_LC_4_1_1.SEQ_MODE=4'b0000;
    defparam testClock_RNIAQVB_LC_4_1_1.LUT_INIT=16'b1110111101000000;
    LogicCell40 testClock_RNIAQVB_LC_4_1_1 (
            .in0(N__41338),
            .in1(N__30290),
            .in2(N__30780),
            .in3(N__17743),
            .lcout(testClock_0),
            .ltout(testClock_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_cnv_0_0_LC_4_1_2 .C_ON=1'b0;
    defparam \ALU.a_cnv_0_0_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.a_cnv_0_0_LC_4_1_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \ALU.a_cnv_0_0_LC_4_1_2  (
            .in0(N__17744),
            .in1(_gnd_net_),
            .in2(N__17777),
            .in3(N__17764),
            .lcout(\ALU.a_cnv_0Z0Z_0 ),
            .ltout(\ALU.a_cnv_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_cnv_0_LC_4_1_3 .C_ON=1'b0;
    defparam \ALU.a_cnv_0_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.a_cnv_0_LC_4_1_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.a_cnv_0_LC_4_1_3  (
            .in0(N__20435),
            .in1(N__17852),
            .in2(N__17774),
            .in3(N__17925),
            .lcout(\ALU.a_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m52_LC_4_1_4 .C_ON=1'b0;
    defparam \ALU.m52_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m52_LC_4_1_4 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \ALU.m52_LC_4_1_4  (
            .in0(N__22438),
            .in1(N__22729),
            .in2(N__22599),
            .in3(N__44038),
            .lcout(\ALU.N_53_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testClock_LC_4_1_5.C_ON=1'b0;
    defparam testClock_LC_4_1_5.SEQ_MODE=4'b1000;
    defparam testClock_LC_4_1_5.LUT_INIT=16'b1110111101000000;
    LogicCell40 testClock_LC_4_1_5 (
            .in0(N__41340),
            .in1(N__30291),
            .in2(N__30782),
            .in3(N__17746),
            .lcout(testClockZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47630),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_cnv_0_0_LC_4_1_6 .C_ON=1'b0;
    defparam \ALU.b_cnv_0_0_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.b_cnv_0_0_LC_4_1_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \ALU.b_cnv_0_0_LC_4_1_6  (
            .in0(N__17745),
            .in1(N__17765),
            .in2(_gnd_net_),
            .in3(N__17753),
            .lcout(\ALU.b_cnv_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_2_LC_4_1_7.C_ON=1'b0;
    defparam testState_2_LC_4_1_7.SEQ_MODE=4'b1000;
    defparam testState_2_LC_4_1_7.LUT_INIT=16'b0101100001010000;
    LogicCell40 testState_2_LC_4_1_7 (
            .in0(N__41339),
            .in1(N__21895),
            .in2(N__30781),
            .in3(N__30292),
            .lcout(testStateZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47630),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_cnv_0_LC_4_2_1 .C_ON=1'b0;
    defparam \ALU.e_cnv_0_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_cnv_0_LC_4_2_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ALU.e_cnv_0_LC_4_2_1  (
            .in0(N__17938),
            .in1(N__17847),
            .in2(N__17927),
            .in3(N__20455),
            .lcout(\ALU.e_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_cnv_0_LC_4_2_2 .C_ON=1'b0;
    defparam \ALU.c_cnv_0_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_cnv_0_LC_4_2_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ALU.c_cnv_0_LC_4_2_2  (
            .in0(N__20454),
            .in1(N__17921),
            .in2(N__17853),
            .in3(N__17937),
            .lcout(\ALU.c_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.G_566_LC_4_2_3 .C_ON=1'b0;
    defparam \ALU.G_566_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.G_566_LC_4_2_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ALU.G_566_LC_4_2_3  (
            .in0(N__41399),
            .in1(N__30314),
            .in2(N__30783),
            .in3(N__17747),
            .lcout(G_566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_cnv_0_LC_4_2_4 .C_ON=1'b0;
    defparam \ALU.g_cnv_0_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.g_cnv_0_LC_4_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.g_cnv_0_LC_4_2_4  (
            .in0(N__17926),
            .in1(N__17939),
            .in2(N__17855),
            .in3(N__20458),
            .lcout(\ALU.g_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_cnv_0_LC_4_2_5 .C_ON=1'b0;
    defparam \ALU.b_cnv_0_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.b_cnv_0_LC_4_2_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \ALU.b_cnv_0_LC_4_2_5  (
            .in0(N__17917),
            .in1(N__20453),
            .in2(N__17883),
            .in3(N__17840),
            .lcout(\ALU.b_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_cnv_0_LC_4_2_6 .C_ON=1'b0;
    defparam \ALU.d_cnv_0_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_cnv_0_LC_4_2_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ALU.d_cnv_0_LC_4_2_6  (
            .in0(N__17882),
            .in1(N__17922),
            .in2(N__17854),
            .in3(N__20457),
            .lcout(\ALU.d_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_cnv_0_LC_4_2_7 .C_ON=1'b0;
    defparam \ALU.f_cnv_0_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.f_cnv_0_LC_4_2_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ALU.f_cnv_0_LC_4_2_7  (
            .in0(N__17923),
            .in1(N__20456),
            .in2(N__17884),
            .in3(N__17848),
            .lcout(\ALU.f_cnvZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIEP354_14_LC_4_3_0 .C_ON=1'b0;
    defparam \ALU.c_RNIEP354_14_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIEP354_14_LC_4_3_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \ALU.c_RNIEP354_14_LC_4_3_0  (
            .in0(N__17813),
            .in1(N__40616),
            .in2(_gnd_net_),
            .in3(N__29377),
            .lcout(),
            .ltout(\ALU.c_RNIEP354Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI25K7D_14_LC_4_3_1 .C_ON=1'b0;
    defparam \ALU.c_RNI25K7D_14_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI25K7D_14_LC_4_3_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.c_RNI25K7D_14_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(N__43109),
            .in2(N__17786),
            .in3(N__17783),
            .lcout(\ALU.a_15_m3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJENJ8_0_15_LC_4_3_2 .C_ON=1'b0;
    defparam \ALU.c_RNIJENJ8_0_15_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJENJ8_0_15_LC_4_3_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \ALU.c_RNIJENJ8_0_15_LC_4_3_2  (
            .in0(N__38432),
            .in1(N__38647),
            .in2(N__39082),
            .in3(N__44334),
            .lcout(\ALU.c_RNIJENJ8_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJENJ8_15_LC_4_3_3 .C_ON=1'b0;
    defparam \ALU.c_RNIJENJ8_15_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJENJ8_15_LC_4_3_3 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \ALU.c_RNIJENJ8_15_LC_4_3_3  (
            .in0(N__38646),
            .in1(N__39053),
            .in2(N__44403),
            .in3(N__38431),
            .lcout(\ALU.rshift_15_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIR45G7_6_LC_4_3_4 .C_ON=1'b0;
    defparam \ALU.d_RNIR45G7_6_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIR45G7_6_LC_4_3_4 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.d_RNIR45G7_6_LC_4_3_4  (
            .in0(N__43697),
            .in1(N__46960),
            .in2(N__39081),
            .in3(N__46735),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIS6U9F_9_LC_4_3_5 .C_ON=1'b0;
    defparam \ALU.d_RNIS6U9F_9_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIS6U9F_9_LC_4_3_5 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNIS6U9F_9_LC_4_3_5  (
            .in0(N__39851),
            .in1(N__39054),
            .in2(N__17981),
            .in3(N__40071),
            .lcout(\ALU.N_474 ),
            .ltout(\ALU.N_474_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNII2IF91_9_LC_4_3_6 .C_ON=1'b0;
    defparam \ALU.d_RNII2IF91_9_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNII2IF91_9_LC_4_3_6 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \ALU.d_RNII2IF91_9_LC_4_3_6  (
            .in0(N__44323),
            .in1(N__19445),
            .in2(N__17978),
            .in3(N__17975),
            .lcout(),
            .ltout(\ALU.rshift_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIL01TD1_6_LC_4_3_7 .C_ON=1'b0;
    defparam \ALU.d_RNIL01TD1_6_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIL01TD1_6_LC_4_3_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \ALU.d_RNIL01TD1_6_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__43110),
            .in2(N__17969),
            .in3(N__17966),
            .lcout(\ALU.d_RNIL01TD1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIKJTS7_15_LC_4_4_0 .C_ON=1'b0;
    defparam \ALU.c_RNIKJTS7_15_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIKJTS7_15_LC_4_4_0 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \ALU.c_RNIKJTS7_15_LC_4_4_0  (
            .in0(N__40619),
            .in1(N__39076),
            .in2(N__32665),
            .in3(N__43667),
            .lcout(\ALU.lshift_3_ns_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3FQF1_14_LC_4_4_1 .C_ON=1'b0;
    defparam \ALU.c_RNI3FQF1_14_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3FQF1_14_LC_4_4_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNI3FQF1_14_LC_4_4_1  (
            .in0(N__35401),
            .in1(N__33692),
            .in2(N__19475),
            .in3(N__31556),
            .lcout(\ALU.N_713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNITDBD1_14_LC_4_4_2 .C_ON=1'b0;
    defparam \ALU.b_RNITDBD1_14_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNITDBD1_14_LC_4_4_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.b_RNITDBD1_14_LC_4_4_2  (
            .in0(N__28298),
            .in1(N__35761),
            .in2(N__28322),
            .in3(N__35588),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI81K02_14_LC_4_4_3 .C_ON=1'b0;
    defparam \ALU.d_RNI81K02_14_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI81K02_14_LC_4_4_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI81K02_14_LC_4_4_3  (
            .in0(N__35402),
            .in1(N__30620),
            .in2(N__17957),
            .in3(N__30596),
            .lcout(\ALU.N_761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIN38K3_15_LC_4_4_4 .C_ON=1'b0;
    defparam \ALU.c_RNIN38K3_15_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIN38K3_15_LC_4_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIN38K3_15_LC_4_4_4  (
            .in0(N__30556),
            .in1(N__30536),
            .in2(_gnd_net_),
            .in3(N__35243),
            .lcout(\ALU.aluOut_15 ),
            .ltout(\ALU.aluOut_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3QSJ7_15_LC_4_4_5 .C_ON=1'b0;
    defparam \ALU.c_RNI3QSJ7_15_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3QSJ7_15_LC_4_4_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNI3QSJ7_15_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(N__43653),
            .in2(N__17954),
            .in3(N__40618),
            .lcout(\ALU.N_590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFR7K3_14_LC_4_4_6 .C_ON=1'b0;
    defparam \ALU.c_RNIFR7K3_14_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFR7K3_14_LC_4_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIFR7K3_14_LC_4_4_6  (
            .in0(N__17951),
            .in1(N__17945),
            .in2(_gnd_net_),
            .in3(N__35242),
            .lcout(\ALU.aluOut_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_14_LC_4_5_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_14_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_14_LC_4_5_0 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.a_15_m2_ns_1_14_LC_4_5_0  (
            .in0(N__47292),
            .in1(N__44089),
            .in2(N__43919),
            .in3(N__43668),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI58CHC_14_LC_4_5_1 .C_ON=1'b0;
    defparam \ALU.c_RNI58CHC_14_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI58CHC_14_LC_4_5_1 .LUT_INIT=16'b1000011001100111;
    LogicCell40 \ALU.c_RNI58CHC_14_LC_4_5_1  (
            .in0(N__47293),
            .in1(N__40617),
            .in2(N__18011),
            .in3(N__21304),
            .lcout(\ALU.a_15_m2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIB9KD11_11_LC_4_5_2 .C_ON=1'b0;
    defparam \ALU.c_RNIB9KD11_11_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIB9KD11_11_LC_4_5_2 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.c_RNIB9KD11_11_LC_4_5_2  (
            .in0(N__38732),
            .in1(N__19463),
            .in2(N__44523),
            .in3(N__20789),
            .lcout(),
            .ltout(\ALU.lshift_15_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAD5QQ1_0_LC_4_5_3 .C_ON=1'b0;
    defparam \ALU.d_RNIAD5QQ1_0_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAD5QQ1_0_LC_4_5_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.d_RNIAD5QQ1_0_LC_4_5_3  (
            .in0(N__44491),
            .in1(N__39200),
            .in2(N__18008),
            .in3(N__39185),
            .lcout(),
            .ltout(\ALU.lshift_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIEGAQ72_14_LC_4_5_4 .C_ON=1'b0;
    defparam \ALU.c_RNIEGAQ72_14_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIEGAQ72_14_LC_4_5_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.c_RNIEGAQ72_14_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__44090),
            .in2(N__18005),
            .in3(N__18002),
            .lcout(),
            .ltout(\ALU.a_15_m4_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFCGVL2_14_LC_4_5_5 .C_ON=1'b0;
    defparam \ALU.c_RNIFCGVL2_14_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFCGVL2_14_LC_4_5_5 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \ALU.c_RNIFCGVL2_14_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__46331),
            .in2(N__17996),
            .in3(N__17993),
            .lcout(c_RNIFCGVL2_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI63LF1_12_LC_4_6_0 .C_ON=1'b0;
    defparam \ALU.a_RNI63LF1_12_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI63LF1_12_LC_4_6_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.a_RNI63LF1_12_LC_4_6_0  (
            .in0(N__35910),
            .in1(N__28565),
            .in2(N__36005),
            .in3(N__28211),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBAHQ1_12_LC_4_6_1 .C_ON=1'b0;
    defparam \ALU.c_RNIBAHQ1_12_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBAHQ1_12_LC_4_6_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNIBAHQ1_12_LC_4_6_1  (
            .in0(N__35394),
            .in1(N__33962),
            .in2(N__17984),
            .in3(N__31286),
            .lcout(\ALU.N_711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIP9BD1_12_LC_4_6_2 .C_ON=1'b0;
    defparam \ALU.b_RNIP9BD1_12_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIP9BD1_12_LC_4_6_2 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \ALU.b_RNIP9BD1_12_LC_4_6_2  (
            .in0(N__35762),
            .in1(N__28370),
            .in2(N__28349),
            .in3(N__35577),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0PJ02_12_LC_4_6_3 .C_ON=1'b0;
    defparam \ALU.d_RNI0PJ02_12_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0PJ02_12_LC_4_6_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI0PJ02_12_LC_4_6_3  (
            .in0(N__35395),
            .in1(N__25499),
            .in2(N__18170),
            .in3(N__28394),
            .lcout(),
            .ltout(\ALU.N_759_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFEUU3_12_LC_4_6_4 .C_ON=1'b0;
    defparam \ALU.c_RNIFEUU3_12_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFEUU3_12_LC_4_6_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.c_RNIFEUU3_12_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(N__18167),
            .in2(N__18161),
            .in3(N__35241),
            .lcout(\ALU.aluOut_12 ),
            .ltout(\ALU.aluOut_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIIUNC7_12_LC_4_6_5 .C_ON=1'b0;
    defparam \ALU.c_RNIIUNC7_12_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIIUNC7_12_LC_4_6_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ALU.c_RNIIUNC7_12_LC_4_6_5  (
            .in0(N__37245),
            .in1(_gnd_net_),
            .in2(N__18158),
            .in3(_gnd_net_),
            .lcout(\ALU.a12_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA6K08_4_LC_4_7_0 .C_ON=1'b0;
    defparam \ALU.d_RNIA6K08_4_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA6K08_4_LC_4_7_0 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIA6K08_4_LC_4_7_0  (
            .in0(N__23446),
            .in1(N__39821),
            .in2(N__30014),
            .in3(N__23567),
            .lcout(\ALU.a9_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_20_LC_4_7_1.C_ON=1'b0;
    defparam testWord_20_LC_4_7_1.SEQ_MODE=4'b1000;
    defparam testWord_20_LC_4_7_1.LUT_INIT=16'b1100101010101010;
    LogicCell40 testWord_20_LC_4_7_1 (
            .in0(N__18022),
            .in1(N__32292),
            .in2(N__41478),
            .in3(N__18138),
            .lcout(ctrlOut_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47670),
            .ce(N__41057),
            .sr(_gnd_net_));
    defparam \ALU.m234_LC_4_7_2 .C_ON=1'b0;
    defparam \ALU.m234_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.m234_LC_4_7_2 .LUT_INIT=16'b1011111111110101;
    LogicCell40 \ALU.m234_LC_4_7_2  (
            .in0(N__29681),
            .in1(N__18061),
            .in2(N__25164),
            .in3(N__30136),
            .lcout(\ALU.N_235_0 ),
            .ltout(\ALU.N_235_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRNNS7_3_LC_4_7_3 .C_ON=1'b0;
    defparam \ALU.d_RNIRNNS7_3_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRNNS7_3_LC_4_7_3 .LUT_INIT=16'b0100110000001000;
    LogicCell40 \ALU.d_RNIRNNS7_3_LC_4_7_3  (
            .in0(N__29955),
            .in1(N__25288),
            .in2(N__18029),
            .in3(N__24043),
            .lcout(),
            .ltout(\ALU.a12_b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_11_LC_4_7_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_11_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_11_LC_4_7_4 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_484_11_LC_4_7_4  (
            .in0(N__40626),
            .in1(N__23366),
            .in2(N__18026),
            .in3(N__37761),
            .lcout(\ALU.madd_484_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m228_LC_4_7_5 .C_ON=1'b0;
    defparam \ALU.m228_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.m228_LC_4_7_5 .LUT_INIT=16'b1110111001111111;
    LogicCell40 \ALU.m228_LC_4_7_5  (
            .in0(N__30135),
            .in1(N__25118),
            .in2(N__18023),
            .in3(N__29682),
            .lcout(\ALU.N_229_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIOVJ78_3_LC_4_7_6 .C_ON=1'b0;
    defparam \ALU.d_RNIOVJ78_3_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIOVJ78_3_LC_4_7_6 .LUT_INIT=16'b0010111000000000;
    LogicCell40 \ALU.d_RNIOVJ78_3_LC_4_7_6  (
            .in0(N__24042),
            .in1(N__29954),
            .in2(N__23921),
            .in3(N__27587),
            .lcout(),
            .ltout(\ALU.a10_b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_319_LC_4_7_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_319_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_319_LC_4_7_7 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_319_LC_4_7_7  (
            .in0(N__37760),
            .in1(N__18326),
            .in2(N__18320),
            .in3(N__25289),
            .lcout(\ALU.madd_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_15_LC_4_8_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_15_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_15_LC_4_8_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_484_15_LC_4_8_0  (
            .in0(N__18308),
            .in1(N__19499),
            .in2(N__20396),
            .in3(N__18299),
            .lcout(\ALU.madd_484_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_17_LC_4_8_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_17_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_17_LC_4_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_484_17_LC_4_8_1  (
            .in0(N__19706),
            .in1(N__18293),
            .in2(_gnd_net_),
            .in3(N__20984),
            .lcout(),
            .ltout(\ALU.madd_484_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_20_LC_4_8_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_20_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_20_LC_4_8_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_484_20_LC_4_8_2  (
            .in0(N__18176),
            .in1(N__18221),
            .in2(N__18284),
            .in3(N__18281),
            .lcout(\ALU.madd_484_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_391_LC_4_8_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_391_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_391_LC_4_8_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_391_LC_4_8_3  (
            .in0(N__18362),
            .in1(_gnd_net_),
            .in2(N__18269),
            .in3(N__18245),
            .lcout(\ALU.madd_391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0B2B8_0_7_LC_4_8_4 .C_ON=1'b0;
    defparam \ALU.d_RNI0B2B8_0_7_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0B2B8_0_7_LC_4_8_4 .LUT_INIT=16'b0010001010100000;
    LogicCell40 \ALU.d_RNI0B2B8_0_7_LC_4_8_4  (
            .in0(N__46907),
            .in1(N__19788),
            .in2(N__19106),
            .in3(N__26523),
            .lcout(),
            .ltout(\ALU.a7_b_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_16_LC_4_8_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_16_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_16_LC_4_8_5 .LUT_INIT=16'b0001011111101000;
    LogicCell40 \ALU.mult_madd_484_16_LC_4_8_5  (
            .in0(N__18215),
            .in1(N__18203),
            .in2(N__18185),
            .in3(N__18182),
            .lcout(\ALU.madd_484_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIB0KD9_12_LC_4_9_0 .C_ON=1'b0;
    defparam \ALU.d_RNIB0KD9_12_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIB0KD9_12_LC_4_9_0 .LUT_INIT=16'b0011010111001010;
    LogicCell40 \ALU.d_RNIB0KD9_12_LC_4_9_0  (
            .in0(N__25462),
            .in1(N__20917),
            .in2(N__26597),
            .in3(N__25326),
            .lcout(),
            .ltout(\ALU.un9_addsub_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFKNTE_12_LC_4_9_1 .C_ON=1'b0;
    defparam \ALU.d_RNIFKNTE_12_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFKNTE_12_LC_4_9_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNIFKNTE_12_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18368),
            .in3(N__40848),
            .lcout(\ALU.d_RNIFKNTEZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISHLE5_12_LC_4_9_2 .C_ON=1'b0;
    defparam \ALU.d_RNISHLE5_12_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISHLE5_12_LC_4_9_2 .LUT_INIT=16'b0000010111110101;
    LogicCell40 \ALU.d_RNISHLE5_12_LC_4_9_2  (
            .in0(N__25463),
            .in1(_gnd_net_),
            .in2(N__26596),
            .in3(N__20918),
            .lcout(\ALU.N_180_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIV96U8_13_LC_4_9_3 .C_ON=1'b0;
    defparam \ALU.d_RNIV96U8_13_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIV96U8_13_LC_4_9_3 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNIV96U8_13_LC_4_9_3  (
            .in0(N__25061),
            .in1(N__25008),
            .in2(N__30031),
            .in3(N__38002),
            .lcout(\ALU.d_RNIV96U8Z0Z_13 ),
            .ltout(\ALU.d_RNIV96U8Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_314_LC_4_9_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_314_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_314_LC_4_9_4 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_madd_314_LC_4_9_4  (
            .in0(N__39448),
            .in1(N__36989),
            .in2(N__18365),
            .in3(N__18335),
            .lcout(\ALU.madd_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_310_0_LC_4_9_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_310_0_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_310_0_LC_4_9_5 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_310_0_LC_4_9_5  (
            .in0(N__37418),
            .in1(N__40847),
            .in2(N__37003),
            .in3(N__39447),
            .lcout(\ALU.madd_310_0 ),
            .ltout(\ALU.madd_310_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_334_LC_4_9_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_334_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_334_LC_4_9_6 .LUT_INIT=16'b1011111000101000;
    LogicCell40 \ALU.mult_madd_334_LC_4_9_6  (
            .in0(N__18809),
            .in1(N__18419),
            .in2(N__18347),
            .in3(N__19677),
            .lcout(\ALU.madd_334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIM558_12_LC_4_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNIIM558_12_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIM558_12_LC_4_9_7 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.d_RNIIM558_12_LC_4_9_7  (
            .in0(N__20916),
            .in1(N__37417),
            .in2(N__30030),
            .in3(N__25461),
            .lcout(\ALU.a1_b_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO82C8_9_LC_4_10_0 .C_ON=1'b0;
    defparam \ALU.d_RNIO82C8_9_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO82C8_9_LC_4_10_0 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNIO82C8_9_LC_4_10_0  (
            .in0(N__21098),
            .in1(N__20866),
            .in2(N__30050),
            .in3(N__36985),
            .lcout(),
            .ltout(\ALU.a2_b_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_222_LC_4_10_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_222_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_222_LC_4_10_1 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_222_LC_4_10_1  (
            .in0(N__18575),
            .in1(N__42891),
            .in2(N__18329),
            .in3(N__47100),
            .lcout(\ALU.madd_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI885I7_8_LC_4_10_2 .C_ON=1'b0;
    defparam \ALU.d_RNI885I7_8_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI885I7_8_LC_4_10_2 .LUT_INIT=16'b0100111000000000;
    LogicCell40 \ALU.d_RNI885I7_8_LC_4_10_2  (
            .in0(N__24231),
            .in1(N__18739),
            .in2(N__18668),
            .in3(N__41941),
            .lcout(\ALU.a3_b_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_275_LC_4_10_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_275_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_275_LC_4_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_275_LC_4_10_3  (
            .in0(N__18482),
            .in1(_gnd_net_),
            .in2(N__18515),
            .in3(N__18550),
            .lcout(\ALU.madd_275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_279_LC_4_10_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_279_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_279_LC_4_10_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.mult_madd_279_LC_4_10_4  (
            .in0(N__18549),
            .in1(N__18502),
            .in2(_gnd_net_),
            .in3(N__18481),
            .lcout(),
            .ltout(\ALU.madd_279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_349_LC_4_10_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_349_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_349_LC_4_10_5 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \ALU.mult_madd_349_LC_4_10_5  (
            .in0(N__19684),
            .in1(N__18457),
            .in2(N__18443),
            .in3(N__18386),
            .lcout(\ALU.madd_349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_330_0_LC_4_10_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_330_0_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_330_0_LC_4_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_330_0_LC_4_10_6  (
            .in0(N__18418),
            .in1(N__18397),
            .in2(_gnd_net_),
            .in3(N__18805),
            .lcout(\ALU.madd_330_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIBLBO_10_LC_4_11_0 .C_ON=1'b0;
    defparam \ALU.a_RNIBLBO_10_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIBLBO_10_LC_4_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.a_RNIBLBO_10_LC_4_11_0  (
            .in0(N__28601),
            .in1(N__23708),
            .in2(_gnd_net_),
            .in3(N__45136),
            .lcout(\ALU.a_RNIBLBOZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIF549_10_LC_4_11_1 .C_ON=1'b0;
    defparam \ALU.c_RNIF549_10_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIF549_10_LC_4_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIF549_10_LC_4_11_1  (
            .in0(N__45137),
            .in1(N__34282),
            .in2(_gnd_net_),
            .in3(N__34934),
            .lcout(),
            .ltout(\ALU.c_RNIF549Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIVSRV1_10_LC_4_11_2 .C_ON=1'b0;
    defparam \ALU.c_RNIVSRV1_10_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIVSRV1_10_LC_4_11_2 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \ALU.c_RNIVSRV1_10_LC_4_11_2  (
            .in0(N__32992),
            .in1(N__34513),
            .in2(N__18380),
            .in3(N__18377),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHGJR4_10_LC_4_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIHGJR4_10_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHGJR4_10_LC_4_11_3 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNIHGJR4_10_LC_4_11_3  (
            .in0(N__24404),
            .in1(N__32993),
            .in2(N__18371),
            .in3(N__26801),
            .lcout(\ALU.operand2_10 ),
            .ltout(\ALU.operand2_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIF6179_10_LC_4_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNIF6179_10_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIF6179_10_LC_4_11_4 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \ALU.d_RNIF6179_10_LC_4_11_4  (
            .in0(N__42787),
            .in1(N__30045),
            .in2(N__18839),
            .in3(N__20040),
            .lcout(\ALU.a4_b_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7U079_10_LC_4_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNI7U079_10_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7U079_10_LC_4_11_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.d_RNI7U079_10_LC_4_11_5  (
            .in0(N__20041),
            .in1(N__41959),
            .in2(N__30058),
            .in3(N__20014),
            .lcout(\ALU.a3_b_10 ),
            .ltout(\ALU.a3_b_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_305_LC_4_11_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_305_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_305_LC_4_11_6 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ALU.mult_madd_305_LC_4_11_6  (
            .in0(N__37218),
            .in1(N__39395),
            .in2(N__18812),
            .in3(N__35065),
            .lcout(\ALU.madd_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIV0CK1_7_LC_4_12_0 .C_ON=1'b0;
    defparam \ALU.d_RNIV0CK1_7_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIV0CK1_7_LC_4_12_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.d_RNIV0CK1_7_LC_4_12_0  (
            .in0(N__45374),
            .in1(N__45356),
            .in2(N__35365),
            .in3(N__26906),
            .lcout(\ALU.N_754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_17_LC_4_12_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_17_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_17_LC_4_12_1 .LUT_INIT=16'b1110100011000000;
    LogicCell40 \ALU.mult_madd_17_LC_4_12_1  (
            .in0(N__23188),
            .in1(N__22970),
            .in2(N__23209),
            .in3(N__23165),
            .lcout(\ALU.madd_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_5_LC_4_12_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_5_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_5_LC_4_12_2 .LUT_INIT=16'b1110100010001000;
    LogicCell40 \ALU.mult_madd_5_LC_4_12_2  (
            .in0(N__24481),
            .in1(N__24460),
            .in2(N__37004),
            .in3(N__37651),
            .lcout(\ALU.madd_5 ),
            .ltout(\ALU.madd_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_19_LC_4_12_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_19_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_19_LC_4_12_3 .LUT_INIT=16'b0110000011000000;
    LogicCell40 \ALU.mult_madd_19_LC_4_12_3  (
            .in0(N__37652),
            .in1(N__20240),
            .in2(N__18794),
            .in3(N__41992),
            .lcout(\ALU.madd_19 ),
            .ltout(\ALU.madd_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_58_LC_4_12_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_58_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_58_LC_4_12_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \ALU.mult_madd_58_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__18780),
            .in2(N__18767),
            .in3(N__18764),
            .lcout(\ALU.madd_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_a3_0_1_LC_4_13_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_a3_0_1_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_a3_0_1_LC_4_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.mult_g0_0_a3_0_1_LC_4_13_0  (
            .in0(N__27566),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37659),
            .lcout(\ALU.g0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKRRR6_4_LC_4_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIKRRR6_4_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKRRR6_4_LC_4_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIKRRR6_4_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__42789),
            .in2(_gnd_net_),
            .in3(N__37115),
            .lcout(\ALU.a4_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKT467_8_LC_4_13_2 .C_ON=1'b0;
    defparam \ALU.d_RNIKT467_8_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKT467_8_LC_4_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIKT467_8_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__40056),
            .in2(_gnd_net_),
            .in3(N__38225),
            .lcout(),
            .ltout(\ALU.a8_b_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_93_LC_4_13_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_93_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_93_LC_4_13_3 .LUT_INIT=16'b1111100010000000;
    LogicCell40 \ALU.mult_madd_93_LC_4_13_3  (
            .in0(N__46681),
            .in1(N__37116),
            .in2(N__18911),
            .in3(N__20566),
            .lcout(\ALU.madd_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4KLR6_7_LC_4_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNI4KLR6_7_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4KLR6_7_LC_4_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNI4KLR6_7_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__46813),
            .in2(_gnd_net_),
            .in3(N__37658),
            .lcout(\ALU.a7_b_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_23_LC_4_13_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_23_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_23_LC_4_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_23_LC_4_13_5  (
            .in0(N__37660),
            .in1(N__42788),
            .in2(N__41975),
            .in3(N__37114),
            .lcout(),
            .ltout(\ALU.madd_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_24_LC_4_13_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_24_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_24_LC_4_13_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ALU.mult_madd_24_LC_4_13_6  (
            .in0(N__40425),
            .in1(N__20246),
            .in2(N__18908),
            .in3(N__38226),
            .lcout(\ALU.madd_24 ),
            .ltout(\ALU.madd_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_51_LC_4_13_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_51_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_51_LC_4_13_7 .LUT_INIT=16'b1010000011101000;
    LogicCell40 \ALU.mult_madd_51_LC_4_13_7  (
            .in0(N__18896),
            .in1(N__38001),
            .in2(N__18884),
            .in3(N__46462),
            .lcout(\ALU.madd_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m6_1_LC_4_14_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_m6_1_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m6_1_LC_4_14_0 .LUT_INIT=16'b1101010001110001;
    LogicCell40 \ALU.mult_madd_m6_1_LC_4_14_0  (
            .in0(N__19150),
            .in1(N__19183),
            .in2(N__18881),
            .in3(N__19169),
            .lcout(\ALU.madd_i3_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_37_LC_4_14_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_37_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_37_LC_4_14_1 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_37_LC_4_14_1  (
            .in0(N__40426),
            .in1(N__18862),
            .in2(N__18848),
            .in3(N__37653),
            .lcout(\ALU.madd_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_12_LC_4_14_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_12_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_12_LC_4_14_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \ALU.mult_madd_12_LC_4_14_2  (
            .in0(N__21635),
            .in1(N__21644),
            .in2(N__42971),
            .in3(N__38299),
            .lcout(\ALU.madd_12 ),
            .ltout(\ALU.madd_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_34_LC_4_14_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_34_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_34_LC_4_14_3 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_34_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__18972),
            .in2(N__19025),
            .in3(N__20301),
            .lcout(\ALU.madd_34 ),
            .ltout(\ALU.madd_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_56_LC_4_14_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_56_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_56_LC_4_14_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_56_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__19016),
            .in2(N__19007),
            .in3(N__19002),
            .lcout(\ALU.madd_56 ),
            .ltout(\ALU.madd_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_6_LC_4_14_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_6_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_6_LC_4_14_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_axb_6_LC_4_14_5  (
            .in0(N__19170),
            .in1(N__19151),
            .in2(N__18989),
            .in3(N__19184),
            .lcout(\ALU.madd_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_30_LC_4_14_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_30_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_30_LC_4_14_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_30_LC_4_14_6  (
            .in0(N__20302),
            .in1(_gnd_net_),
            .in2(N__18977),
            .in3(N__18952),
            .lcout(\ALU.madd_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_52_LC_4_14_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_52_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_52_LC_4_14_7 .LUT_INIT=16'b0101011001101010;
    LogicCell40 \ALU.mult_madd_52_LC_4_14_7  (
            .in0(N__18986),
            .in1(N__18976),
            .in2(N__18956),
            .in3(N__20303),
            .lcout(\ALU.madd_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5R097_6_LC_4_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNI5R097_6_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5R097_6_LC_4_15_0 .LUT_INIT=16'b0110110001100011;
    LogicCell40 \ALU.d_RNI5R097_6_LC_4_15_0  (
            .in0(N__26282),
            .in1(N__46626),
            .in2(N__26602),
            .in3(N__26716),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGLK5B_6_LC_4_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIGLK5B_6_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGLK5B_6_LC_4_15_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNIGLK5B_6_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18944),
            .in3(N__46443),
            .lcout(\ALU.d_RNIGLK5BZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_74_0_LC_4_15_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_74_0_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_74_0_LC_4_15_2 .LUT_INIT=16'b0010110111010010;
    LogicCell40 \ALU.mult_madd_74_0_LC_4_15_2  (
            .in0(N__42926),
            .in1(N__41706),
            .in2(N__18941),
            .in3(N__20407),
            .lcout(\ALU.madd_74_0 ),
            .ltout(\ALU.madd_74_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_83_LC_4_15_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_83_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_83_LC_4_15_3 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \ALU.mult_madd_83_LC_4_15_3  (
            .in0(N__19216),
            .in1(N__19171),
            .in2(N__19229),
            .in3(N__19199),
            .lcout(\ALU.madd_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBQJS3_6_LC_4_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNIBQJS3_6_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBQJS3_6_LC_4_15_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \ALU.d_RNIBQJS3_6_LC_4_15_4  (
            .in0(N__24263),
            .in1(N__26281),
            .in2(_gnd_net_),
            .in3(N__26715),
            .lcout(\ALU.N_219_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_79_0_LC_4_15_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_79_0_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_79_0_LC_4_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_79_0_LC_4_15_5  (
            .in0(N__19215),
            .in1(N__19198),
            .in2(_gnd_net_),
            .in3(N__19190),
            .lcout(\ALU.madd_79_0 ),
            .ltout(\ALU.madd_79_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_88_LC_4_15_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_88_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_88_LC_4_15_6 .LUT_INIT=16'b1101111001001000;
    LogicCell40 \ALU.mult_madd_88_LC_4_15_6  (
            .in0(N__19172),
            .in1(N__19149),
            .in2(N__19133),
            .in3(N__19130),
            .lcout(),
            .ltout(\ALU.madd_88_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_7_LC_4_15_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_7_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_7_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_axb_7_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__19306),
            .in2(N__19124),
            .in3(N__19121),
            .lcout(\ALU.madd_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_73_LC_4_16_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_73_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_73_LC_4_16_0 .LUT_INIT=16'b1111001000100000;
    LogicCell40 \ALU.mult_madd_73_LC_4_16_0  (
            .in0(N__37500),
            .in1(N__46449),
            .in2(N__19040),
            .in3(N__19115),
            .lcout(\ALU.madd_73 ),
            .ltout(\ALU.madd_73_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_113_LC_4_16_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_113_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_113_LC_4_16_1 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \ALU.mult_madd_113_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__19333),
            .in2(N__19109),
            .in3(N__21670),
            .lcout(\ALU.madd_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFCMC8_7_LC_4_16_2 .C_ON=1'b0;
    defparam \ALU.d_RNIFCMC8_7_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFCMC8_7_LC_4_16_2 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNIFCMC8_7_LC_4_16_2  (
            .in0(N__19853),
            .in1(N__19098),
            .in2(N__30059),
            .in3(N__37997),
            .lcout(\ALU.a0_b_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_154_LC_4_16_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_154_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_154_LC_4_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_154_LC_4_16_3  (
            .in0(N__19367),
            .in1(N__20347),
            .in2(_gnd_net_),
            .in3(N__19348),
            .lcout(\ALU.madd_154 ),
            .ltout(\ALU.madd_154_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_159_LC_4_16_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_159_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_159_LC_4_16_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.mult_madd_159_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19337),
            .in3(N__19269),
            .lcout(\ALU.madd_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_109_LC_4_16_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_109_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_109_LC_4_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_109_LC_4_16_5  (
            .in0(N__19334),
            .in1(N__21671),
            .in2(_gnd_net_),
            .in3(N__19313),
            .lcout(\ALU.madd_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_9_ma_LC_4_16_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_cry_9_ma_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_9_ma_LC_4_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_madd_cry_9_ma_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__19288),
            .in2(_gnd_net_),
            .in3(N__19270),
            .lcout(\ALU.madd_cry_9_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m271_ns_1_LC_4_16_7 .C_ON=1'b0;
    defparam \ALU.m271_ns_1_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m271_ns_1_LC_4_16_7 .LUT_INIT=16'b0000001110000000;
    LogicCell40 \ALU.m271_ns_1_LC_4_16_7  (
            .in0(N__24922),
            .in1(N__30215),
            .in2(N__26627),
            .in3(N__29753),
            .lcout(\ALU.m271_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_e_0_3_LC_5_1_0 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_e_0_3_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_e_0_3_LC_5_1_0 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \CONTROL.aluOperation_e_0_3_LC_5_1_0  (
            .in0(N__33317),
            .in1(N__33385),
            .in2(N__19256),
            .in3(N__19406),
            .lcout(aluOperation_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47622),
            .ce(N__33442),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m5s2_LC_5_1_1 .C_ON=1'b0;
    defparam \ALU.a_15_m5s2_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m5s2_LC_5_1_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALU.a_15_m5s2_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__20478),
            .in2(_gnd_net_),
            .in3(N__44029),
            .lcout(\ALU.a_15_sm3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m282_LC_5_1_2 .C_ON=1'b0;
    defparam \ALU.m282_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \ALU.m282_LC_5_1_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ALU.m282_LC_5_1_2  (
            .in0(N__22440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22573),
            .lcout(\ALU.N_283_0 ),
            .ltout(\ALU.N_283_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_e_0_4_LC_5_1_3 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_e_0_4_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_e_0_4_LC_5_1_3 .LUT_INIT=16'b1100000000100010;
    LogicCell40 \CONTROL.aluOperation_e_0_4_LC_5_1_3  (
            .in0(N__33384),
            .in1(N__19244),
            .in2(N__19232),
            .in3(N__33318),
            .lcout(aluOperation_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47622),
            .ce(N__33442),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_e_0_2_LC_5_1_4 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_e_0_2_LC_5_1_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_e_0_2_LC_5_1_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CONTROL.aluOperation_e_0_2_LC_5_1_4  (
            .in0(N__33316),
            .in1(N__19430),
            .in2(_gnd_net_),
            .in3(N__19418),
            .lcout(aluOperation_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47622),
            .ce(N__33442),
            .sr(_gnd_net_));
    defparam \ALU.m650_ns_1_LC_5_1_5 .C_ON=1'b0;
    defparam \ALU.m650_ns_1_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.m650_ns_1_LC_5_1_5 .LUT_INIT=16'b0011110100001010;
    LogicCell40 \ALU.m650_ns_1_LC_5_1_5  (
            .in0(N__45697),
            .in1(N__22441),
            .in2(N__22596),
            .in3(N__22724),
            .lcout(),
            .ltout(\ALU.m650_nsZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m650_ns_LC_5_1_6 .C_ON=1'b0;
    defparam \ALU.m650_ns_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m650_ns_LC_5_1_6 .LUT_INIT=16'b1001101000010010;
    LogicCell40 \ALU.m650_ns_LC_5_1_6  (
            .in0(N__22725),
            .in1(N__22299),
            .in2(N__19409),
            .in3(N__19405),
            .lcout(N_727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m14_LC_5_1_7 .C_ON=1'b0;
    defparam \ALU.m14_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m14_LC_5_1_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ALU.m14_LC_5_1_7  (
            .in0(N__22569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22439),
            .lcout(\ALU.N_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_1_LC_5_2_0 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_1_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperation_1_LC_5_2_0 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \CONTROL.aluOperation_1_LC_5_2_0  (
            .in0(N__33438),
            .in1(N__45698),
            .in2(N__33335),
            .in3(N__19397),
            .lcout(aluOperation_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47631),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINJ76G_13_LC_5_2_1 .C_ON=1'b0;
    defparam \ALU.c_RNINJ76G_13_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINJ76G_13_LC_5_2_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNINJ76G_13_LC_5_2_1  (
            .in0(N__38923),
            .in1(N__38755),
            .in2(_gnd_net_),
            .in3(N__38437),
            .lcout(),
            .ltout(\ALU.N_577_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIN1J811_11_LC_5_2_2 .C_ON=1'b0;
    defparam \ALU.c_RNIN1J811_11_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIN1J811_11_LC_5_2_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNIN1J811_11_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__38696),
            .in2(N__19391),
            .in3(N__20122),
            .lcout(\ALU.N_633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHDLLS_3_LC_5_2_3 .C_ON=1'b0;
    defparam \ALU.d_RNIHDLLS_3_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHDLLS_3_LC_5_2_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIHDLLS_3_LC_5_2_3  (
            .in0(N__38697),
            .in1(N__20147),
            .in2(_gnd_net_),
            .in3(N__22985),
            .lcout(),
            .ltout(\ALU.N_528_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8DL9U1_3_LC_5_2_4 .C_ON=1'b0;
    defparam \ALU.d_RNI8DL9U1_3_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8DL9U1_3_LC_5_2_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNI8DL9U1_3_LC_5_2_4  (
            .in0(N__44480),
            .in1(_gnd_net_),
            .in2(N__19388),
            .in3(N__19378),
            .lcout(),
            .ltout(\ALU.d_RNI8DL9U1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7AI932_0_LC_5_2_5 .C_ON=1'b0;
    defparam \ALU.d_RNI7AI932_0_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7AI932_0_LC_5_2_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNI7AI932_0_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(N__43097),
            .in2(N__19454),
            .in3(N__19601),
            .lcout(\ALU.a_15_m3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m713_LC_5_2_6 .C_ON=1'b0;
    defparam \ALU.m713_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m713_LC_5_2_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ALU.m713_LC_5_2_6  (
            .in0(N__44060),
            .in1(N__38922),
            .in2(_gnd_net_),
            .in3(N__43491),
            .lcout(\ALU.log_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID35S7_9_LC_5_3_0 .C_ON=1'b0;
    defparam \ALU.d_RNID35S7_9_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID35S7_9_LC_5_3_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ALU.d_RNID35S7_9_LC_5_3_0  (
            .in0(N__40070),
            .in1(_gnd_net_),
            .in2(N__39837),
            .in3(N__43511),
            .lcout(\ALU.N_221 ),
            .ltout(\ALU.N_221_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIDIAPG_11_LC_5_3_1 .C_ON=1'b0;
    defparam \ALU.c_RNIDIAPG_11_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIDIAPG_11_LC_5_3_1 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \ALU.c_RNIDIAPG_11_LC_5_3_1  (
            .in0(N__39044),
            .in1(N__22934),
            .in2(N__19451),
            .in3(_gnd_net_),
            .lcout(\ALU.N_253 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI30A98_13_LC_5_3_2 .C_ON=1'b0;
    defparam \ALU.c_RNI30A98_13_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI30A98_13_LC_5_3_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNI30A98_13_LC_5_3_2  (
            .in0(N__43545),
            .in1(N__40765),
            .in2(_gnd_net_),
            .in3(N__25340),
            .lcout(\ALU.N_588 ),
            .ltout(\ALU.N_588_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3FF6H_11_LC_5_3_3 .C_ON=1'b0;
    defparam \ALU.c_RNI3FF6H_11_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3FF6H_11_LC_5_3_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.c_RNI3FF6H_11_LC_5_3_3  (
            .in0(N__39045),
            .in1(_gnd_net_),
            .in2(N__19448),
            .in3(N__20720),
            .lcout(\ALU.N_575 ),
            .ltout(\ALU.N_575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIMVPEP_15_LC_5_3_4 .C_ON=1'b0;
    defparam \ALU.c_RNIMVPEP_15_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIMVPEP_15_LC_5_3_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ALU.c_RNIMVPEP_15_LC_5_3_4  (
            .in0(N__38436),
            .in1(N__38652),
            .in2(N__19439),
            .in3(N__39046),
            .lcout(\ALU.N_635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI1HUMG_11_LC_5_3_5 .C_ON=1'b0;
    defparam \ALU.c_RNI1HUMG_11_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI1HUMG_11_LC_5_3_5 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.c_RNI1HUMG_11_LC_5_3_5  (
            .in0(N__19436),
            .in1(N__39384),
            .in2(N__39080),
            .in3(N__27608),
            .lcout(\ALU.N_476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIURRD4_0_LC_5_3_6 .C_ON=1'b0;
    defparam \ALU.d_RNIURRD4_0_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIURRD4_0_LC_5_3_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ALU.d_RNIURRD4_0_LC_5_3_6  (
            .in0(N__39015),
            .in1(N__38653),
            .in2(N__43638),
            .in3(N__38028),
            .lcout(\ALU.N_415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIUS558_9_LC_5_3_7 .C_ON=1'b0;
    defparam \ALU.d_RNIUS558_9_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIUS558_9_LC_5_3_7 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.d_RNIUS558_9_LC_5_3_7  (
            .in0(N__43510),
            .in1(N__39795),
            .in2(N__39079),
            .in3(N__40069),
            .lcout(\ALU.rshift_3_ns_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBIR3G_13_LC_5_4_0 .C_ON=1'b0;
    defparam \ALU.c_RNIBIR3G_13_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBIR3G_13_LC_5_4_0 .LUT_INIT=16'b1110001100100011;
    LogicCell40 \ALU.c_RNIBIR3G_13_LC_5_4_0  (
            .in0(N__25343),
            .in1(N__19481),
            .in2(N__39077),
            .in3(N__40768),
            .lcout(\ALU.N_257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIQ3U41_14_LC_5_4_1 .C_ON=1'b0;
    defparam \ALU.a_RNIQ3U41_14_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIQ3U41_14_LC_5_4_1 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.a_RNIQ3U41_14_LC_5_4_1  (
            .in0(N__35912),
            .in1(N__30728),
            .in2(N__35587),
            .in3(N__31385),
            .lcout(\ALU.dout_3_ns_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIK6K78_14_LC_5_4_2 .C_ON=1'b0;
    defparam \ALU.c_RNIK6K78_14_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIK6K78_14_LC_5_4_2 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.c_RNIK6K78_14_LC_5_4_2  (
            .in0(N__43673),
            .in1(N__40614),
            .in2(N__39078),
            .in3(N__40766),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIQIGEG_11_LC_5_4_3 .C_ON=1'b0;
    defparam \ALU.c_RNIQIGEG_11_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIQIGEG_11_LC_5_4_3 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.c_RNIQIGEG_11_LC_5_4_3  (
            .in0(N__39387),
            .in1(N__39036),
            .in2(N__19466),
            .in3(N__25344),
            .lcout(\ALU.N_256 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI30A98_0_13_LC_5_4_4 .C_ON=1'b0;
    defparam \ALU.c_RNI30A98_0_13_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI30A98_0_13_LC_5_4_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ALU.c_RNI30A98_0_13_LC_5_4_4  (
            .in0(N__25342),
            .in1(_gnd_net_),
            .in2(N__43719),
            .in3(N__40767),
            .lcout(\ALU.N_225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIID898_0_11_LC_5_4_5 .C_ON=1'b0;
    defparam \ALU.c_RNIID898_0_11_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIID898_0_11_LC_5_4_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.c_RNIID898_0_11_LC_5_4_5  (
            .in0(N__39386),
            .in1(N__43669),
            .in2(_gnd_net_),
            .in3(N__25341),
            .lcout(),
            .ltout(\ALU.N_224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIO0TVG_11_LC_5_4_6 .C_ON=1'b0;
    defparam \ALU.c_RNIO0TVG_11_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIO0TVG_11_LC_5_4_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ALU.c_RNIO0TVG_11_LC_5_4_6  (
            .in0(N__19511),
            .in1(_gnd_net_),
            .in2(N__19457),
            .in3(N__39013),
            .lcout(\ALU.N_254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIG4C2T_1_LC_5_4_7 .C_ON=1'b0;
    defparam \ALU.d_RNIG4C2T_1_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIG4C2T_1_LC_5_4_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ALU.d_RNIG4C2T_1_LC_5_4_7  (
            .in0(N__23008),
            .in1(_gnd_net_),
            .in2(N__20819),
            .in3(N__38728),
            .lcout(\ALU.N_310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_1_LC_5_5_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_1_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_1_LC_5_5_0 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_484_1_LC_5_5_0  (
            .in0(N__42945),
            .in1(N__39586),
            .in2(N__40433),
            .in3(N__39463),
            .lcout(\ALU.madd_484_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINSF07_5_LC_5_5_1 .C_ON=1'b0;
    defparam \ALU.d_RNINSF07_5_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINSF07_5_LC_5_5_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNINSF07_5_LC_5_5_1  (
            .in0(N__43665),
            .in1(N__40423),
            .in2(_gnd_net_),
            .in3(N__42946),
            .lcout(\ALU.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIF7TU3_4_LC_5_5_2 .C_ON=1'b0;
    defparam \ALU.d_RNIF7TU3_4_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIF7TU3_4_LC_5_5_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \ALU.d_RNIF7TU3_4_LC_5_5_2  (
            .in0(N__42947),
            .in1(N__23468),
            .in2(_gnd_net_),
            .in3(N__29426),
            .lcout(\ALU.N_289_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC8LH7_7_LC_5_5_3 .C_ON=1'b0;
    defparam \ALU.d_RNIC8LH7_7_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC8LH7_7_LC_5_5_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNIC8LH7_7_LC_5_5_3  (
            .in0(N__46946),
            .in1(N__43666),
            .in2(_gnd_net_),
            .in3(N__40075),
            .lcout(\ALU.N_220 ),
            .ltout(\ALU.N_220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIR98G_7_LC_5_5_4 .C_ON=1'b0;
    defparam \ALU.d_RNIIR98G_7_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIR98G_7_LC_5_5_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIIR98G_7_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__39014),
            .in2(N__19514),
            .in3(N__19510),
            .lcout(\ALU.N_252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILPJD8_9_LC_5_5_5 .C_ON=1'b0;
    defparam \ALU.d_RNILPJD8_9_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILPJD8_9_LC_5_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNILPJD8_9_LC_5_5_5  (
            .in0(N__43664),
            .in1(N__39836),
            .in2(_gnd_net_),
            .in3(N__27603),
            .lcout(\ALU.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_4_LC_5_5_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_4_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_4_LC_5_5_6 .LUT_INIT=16'b1011010001000100;
    LogicCell40 \ALU.mult_madd_484_4_LC_5_5_6  (
            .in0(N__21488),
            .in1(N__46945),
            .in2(N__32670),
            .in3(N__38324),
            .lcout(\ALU.madd_484_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIDBD49_15_LC_5_5_7 .C_ON=1'b0;
    defparam \ALU.c_RNIDBD49_15_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIDBD49_15_LC_5_5_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.c_RNIDBD49_15_LC_5_5_7  (
            .in0(N__32604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32661),
            .lcout(\ALU.un9_addsub_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILBFG4_2_LC_5_6_0 .C_ON=1'b0;
    defparam \ALU.d_RNILBFG4_2_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILBFG4_2_LC_5_6_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \ALU.d_RNILBFG4_2_LC_5_6_0  (
            .in0(N__19487),
            .in1(N__29380),
            .in2(_gnd_net_),
            .in3(N__36980),
            .lcout(\ALU.d_RNILBFG4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m240_LC_5_6_1 .C_ON=1'b0;
    defparam \ALU.m240_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.m240_LC_5_6_1 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \ALU.m240_LC_5_6_1  (
            .in0(N__19639),
            .in1(N__19660),
            .in2(_gnd_net_),
            .in3(N__20290),
            .lcout(\ALU.N_241_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI59DJ3_2_LC_5_6_2 .C_ON=1'b0;
    defparam \ALU.d_RNI59DJ3_2_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI59DJ3_2_LC_5_6_2 .LUT_INIT=16'b0111000001111111;
    LogicCell40 \ALU.d_RNI59DJ3_2_LC_5_6_2  (
            .in0(N__20289),
            .in1(N__29378),
            .in2(N__26577),
            .in3(N__28730),
            .lcout(\ALU.N_240_0_i ),
            .ltout(\ALU.N_240_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEDJEA_2_LC_5_6_3 .C_ON=1'b0;
    defparam \ALU.d_RNIEDJEA_2_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEDJEA_2_LC_5_6_3 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \ALU.d_RNIEDJEA_2_LC_5_6_3  (
            .in0(N__36979),
            .in1(_gnd_net_),
            .in2(N__19664),
            .in3(N__37201),
            .lcout(\ALU.d_RNIEDJEAZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m10_LC_5_6_4 .C_ON=1'b0;
    defparam \ALU.m10_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m10_LC_5_6_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \ALU.m10_LC_5_6_4  (
            .in0(N__19661),
            .in1(N__19640),
            .in2(_gnd_net_),
            .in3(N__20944),
            .lcout(\ALU.N_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_6_LC_5_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_6_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_6_LC_5_6_5 .LUT_INIT=16'b1000001000100010;
    LogicCell40 \ALU.mult_madd_6_LC_5_6_5  (
            .in0(N__38024),
            .in1(N__41722),
            .in2(N__33148),
            .in3(N__37202),
            .lcout(\ALU.madd_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIUV3H4_0_LC_5_6_6 .C_ON=1'b0;
    defparam \ALU.d_RNIUV3H4_0_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIUV3H4_0_LC_5_6_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \ALU.d_RNIUV3H4_0_LC_5_6_6  (
            .in0(N__19613),
            .in1(N__29379),
            .in2(_gnd_net_),
            .in3(N__38025),
            .lcout(\ALU.d_RNIUV3H4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_0_LC_5_6_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_0_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_0_LC_5_6_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_0_LC_5_6_7  (
            .in0(N__38023),
            .in1(N__37200),
            .in2(N__37002),
            .in3(N__38274),
            .lcout(\ALU.madd_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILU4U8_12_LC_5_7_0 .C_ON=1'b0;
    defparam \ALU.d_RNILU4U8_12_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILU4U8_12_LC_5_7_0 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.d_RNILU4U8_12_LC_5_7_0  (
            .in0(N__20895),
            .in1(N__37981),
            .in2(N__24193),
            .in3(N__25452),
            .lcout(\ALU.a0_b_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_rep1_e_LC_5_7_1 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_rep1_e_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluReadBus_rep1_e_LC_5_7_1 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \CONTROL.aluReadBus_rep1_e_LC_5_7_1  (
            .in0(N__33355),
            .in1(N__19588),
            .in2(N__19562),
            .in3(N__22294),
            .lcout(aluReadBus_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47662),
            .ce(N__34691),
            .sr(_gnd_net_));
    defparam \CONTROL.aluReadBus_fast_e_LC_5_7_2 .C_ON=1'b0;
    defparam \CONTROL.aluReadBus_fast_e_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluReadBus_fast_e_LC_5_7_2 .LUT_INIT=16'b1100110000000101;
    LogicCell40 \CONTROL.aluReadBus_fast_e_LC_5_7_2  (
            .in0(N__22292),
            .in1(N__19558),
            .in2(N__19589),
            .in3(N__33357),
            .lcout(aluReadBus_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47662),
            .ce(N__34691),
            .sr(_gnd_net_));
    defparam \ALU.m246_LC_5_7_3 .C_ON=1'b0;
    defparam \ALU.m246_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m246_LC_5_7_3 .LUT_INIT=16'b1110111001111111;
    LogicCell40 \ALU.m246_LC_5_7_3  (
            .in0(N__30130),
            .in1(N__25122),
            .in2(N__21859),
            .in3(N__29679),
            .lcout(\ALU.N_247_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_e_0_2_LC_5_7_4 .C_ON=1'b0;
    defparam \CONTROL.busState_1_e_0_2_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.busState_1_e_0_2_LC_5_7_4 .LUT_INIT=16'b1100110001010000;
    LogicCell40 \CONTROL.busState_1_e_0_2_LC_5_7_4  (
            .in0(N__22291),
            .in1(N__19557),
            .in2(N__22595),
            .in3(N__33358),
            .lcout(busState_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47662),
            .ce(N__34691),
            .sr(_gnd_net_));
    defparam \CONTROL.busState_1_e_0_0_LC_5_7_5 .C_ON=1'b0;
    defparam \CONTROL.busState_1_e_0_0_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.busState_1_e_0_0_LC_5_7_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \CONTROL.busState_1_e_0_0_LC_5_7_5  (
            .in0(N__33356),
            .in1(N__22293),
            .in2(N__22736),
            .in3(N__19880),
            .lcout(busState_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47662),
            .ce(N__34691),
            .sr(_gnd_net_));
    defparam \ALU.m210_LC_5_7_6 .C_ON=1'b0;
    defparam \ALU.m210_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m210_LC_5_7_6 .LUT_INIT=16'b1011111111110101;
    LogicCell40 \ALU.m210_LC_5_7_6  (
            .in0(N__29678),
            .in1(N__19871),
            .in2(N__25165),
            .in3(N__30129),
            .lcout(\ALU.N_211_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m204_LC_5_7_7 .C_ON=1'b0;
    defparam \ALU.m204_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m204_LC_5_7_7 .LUT_INIT=16'b1110111001111111;
    LogicCell40 \ALU.m204_LC_5_7_7  (
            .in0(N__30131),
            .in1(N__25123),
            .in2(N__19757),
            .in3(N__29680),
            .lcout(\ALU.N_205_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_367_LC_5_8_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_367_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_367_LC_5_8_0 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_367_LC_5_8_0  (
            .in0(N__19697),
            .in1(N__42016),
            .in2(N__19718),
            .in3(N__39452),
            .lcout(\ALU.madd_367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRV558_13_LC_5_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNIRV558_13_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRV558_13_LC_5_8_1 .LUT_INIT=16'b0010101000100000;
    LogicCell40 \ALU.d_RNIRV558_13_LC_5_8_1  (
            .in0(N__37429),
            .in1(N__25060),
            .in2(N__29994),
            .in3(N__24999),
            .lcout(\ALU.d_RNIRV558Z0Z_13 ),
            .ltout(\ALU.d_RNIRV558Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_371_LC_5_8_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_371_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_371_LC_5_8_2 .LUT_INIT=16'b1110100010100000;
    LogicCell40 \ALU.mult_madd_371_LC_5_8_2  (
            .in0(N__19696),
            .in1(N__42017),
            .in2(N__19709),
            .in3(N__39453),
            .lcout(\ALU.madd_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBAHT8_12_LC_5_8_3 .C_ON=1'b0;
    defparam \ALU.d_RNIBAHT8_12_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBAHT8_12_LC_5_8_3 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \ALU.d_RNIBAHT8_12_LC_5_8_3  (
            .in0(N__20915),
            .in1(N__36981),
            .in2(N__29993),
            .in3(N__25453),
            .lcout(\ALU.a2_b_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_259_LC_5_8_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_259_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_259_LC_5_8_4 .LUT_INIT=16'b1110101010000000;
    LogicCell40 \ALU.mult_madd_259_LC_5_8_4  (
            .in0(N__19930),
            .in1(N__37769),
            .in2(N__39383),
            .in3(N__19937),
            .lcout(\ALU.madd_259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMIK85_11_LC_5_8_5 .C_ON=1'b0;
    defparam \ALU.d_RNIMIK85_11_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMIK85_11_LC_5_8_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ALU.d_RNIMIK85_11_LC_5_8_5  (
            .in0(N__24909),
            .in1(N__24134),
            .in2(N__31180),
            .in3(N__29310),
            .lcout(\ALU.N_186_0 ),
            .ltout(\ALU.N_186_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3JLT7_1_LC_5_8_6 .C_ON=1'b0;
    defparam \ALU.d_RNI3JLT7_1_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3JLT7_1_LC_5_8_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNI3JLT7_1_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19940),
            .in3(N__37428),
            .lcout(\ALU.a1_b_11 ),
            .ltout(\ALU.a1_b_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_255_LC_5_8_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_255_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_255_LC_5_8_7 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_255_LC_5_8_7  (
            .in0(N__37768),
            .in1(N__19931),
            .in2(N__19922),
            .in3(N__39341),
            .lcout(\ALU.madd_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIU5N11_8_LC_5_9_0 .C_ON=1'b0;
    defparam \ALU.e_RNIU5N11_8_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIU5N11_8_LC_5_9_0 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \ALU.e_RNIU5N11_8_LC_5_9_0  (
            .in0(N__31067),
            .in1(N__27349),
            .in2(N__30974),
            .in3(N__27134),
            .lcout(\ALU.dout_3_ns_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIIIOA1_8_LC_5_9_1 .C_ON=1'b0;
    defparam \ALU.f_RNIIIOA1_8_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIIIOA1_8_LC_5_9_1 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.f_RNIIIOA1_8_LC_5_9_1  (
            .in0(N__35989),
            .in1(N__47719),
            .in2(N__25654),
            .in3(N__35899),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI35CK1_8_LC_5_9_2 .C_ON=1'b0;
    defparam \ALU.d_RNI35CK1_8_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI35CK1_8_LC_5_9_2 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNI35CK1_8_LC_5_9_2  (
            .in0(N__25595),
            .in1(N__35366),
            .in2(N__19898),
            .in3(N__25628),
            .lcout(\ALU.N_755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNITF602_8_LC_5_9_3 .C_ON=1'b0;
    defparam \ALU.g_RNITF602_8_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNITF602_8_LC_5_9_3 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \ALU.g_RNITF602_8_LC_5_9_3  (
            .in0(N__30908),
            .in1(N__35737),
            .in2(N__30941),
            .in3(N__19895),
            .lcout(),
            .ltout(\ALU.N_707_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI40CO3_8_LC_5_9_4 .C_ON=1'b0;
    defparam \ALU.d_RNI40CO3_8_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI40CO3_8_LC_5_9_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNI40CO3_8_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__35231),
            .in2(N__19889),
            .in3(N__19886),
            .lcout(\ALU.aluOut_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_26_LC_5_10_0.C_ON=1'b0;
    defparam testWord_26_LC_5_10_0.SEQ_MODE=4'b1000;
    defparam testWord_26_LC_5_10_0.LUT_INIT=16'b1110001010101010;
    LogicCell40 testWord_26_LC_5_10_0 (
            .in0(N__20089),
            .in1(N__41501),
            .in2(N__41563),
            .in3(N__41230),
            .lcout(ctrlOut_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47678),
            .ce(N__41055),
            .sr(_gnd_net_));
    defparam \ALU.m272_ns_1_LC_5_10_1 .C_ON=1'b0;
    defparam \ALU.m272_ns_1_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.m272_ns_1_LC_5_10_1 .LUT_INIT=16'b0000010110000000;
    LogicCell40 \ALU.m272_ns_1_LC_5_10_1  (
            .in0(N__30172),
            .in1(N__20087),
            .in2(N__26651),
            .in3(N__29704),
            .lcout(),
            .ltout(\ALU.m272_nsZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIEUU85_10_LC_5_10_2 .C_ON=1'b0;
    defparam \ALU.c_RNIEUU85_10_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIEUU85_10_LC_5_10_2 .LUT_INIT=16'b0000111101110111;
    LogicCell40 \ALU.c_RNIEUU85_10_LC_5_10_2  (
            .in0(N__20088),
            .in1(N__29367),
            .in2(N__20111),
            .in3(N__27540),
            .lcout(\ALU.N_273_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g0_7_a3_0_0_LC_5_10_3 .C_ON=1'b0;
    defparam \ALU.g0_7_a3_0_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.g0_7_a3_0_0_LC_5_10_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \ALU.g0_7_a3_0_0_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__20082),
            .in2(_gnd_net_),
            .in3(N__29701),
            .lcout(\ALU.g0_7_a3_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g0_6_LC_5_10_4 .C_ON=1'b0;
    defparam \ALU.g0_6_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.g0_6_LC_5_10_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ALU.g0_6_LC_5_10_4  (
            .in0(N__29703),
            .in1(N__30021),
            .in2(N__20090),
            .in3(N__30171),
            .lcout(\ALU.N_191_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m190_LC_5_10_5 .C_ON=1'b0;
    defparam \ALU.m190_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.m190_LC_5_10_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ALU.m190_LC_5_10_5  (
            .in0(N__30170),
            .in1(N__20083),
            .in2(N__24235),
            .in3(N__29702),
            .lcout(\ALU.N_191_0 ),
            .ltout(\ALU.N_191_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBRVD8_10_LC_5_10_6 .C_ON=1'b0;
    defparam \ALU.d_RNIBRVD8_10_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBRVD8_10_LC_5_10_6 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \ALU.d_RNIBRVD8_10_LC_5_10_6  (
            .in0(N__30026),
            .in1(N__37391),
            .in2(N__20027),
            .in3(N__20013),
            .lcout(\ALU.a1_b_10 ),
            .ltout(\ALU.a1_b_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_203_LC_5_10_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_203_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_203_LC_5_10_7 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_203_LC_5_10_7  (
            .in0(N__39334),
            .in1(N__19954),
            .in2(N__19985),
            .in3(N__38213),
            .lcout(\ALU.madd_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFO567_9_LC_5_11_0 .C_ON=1'b0;
    defparam \ALU.d_RNIFO567_9_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFO567_9_LC_5_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIFO567_9_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__39752),
            .in2(_gnd_net_),
            .in3(N__37145),
            .lcout(\ALU.a9_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI08N11_9_LC_5_11_1 .C_ON=1'b0;
    defparam \ALU.e_RNI08N11_9_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI08N11_9_LC_5_11_1 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \ALU.e_RNI08N11_9_LC_5_11_1  (
            .in0(N__38405),
            .in1(N__38375),
            .in2(N__27353),
            .in3(N__27133),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNI1K602_9_LC_5_11_2 .C_ON=1'b0;
    defparam \ALU.g_RNI1K602_9_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNI1K602_9_LC_5_11_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.g_RNI1K602_9_LC_5_11_2  (
            .in0(N__35748),
            .in1(N__36131),
            .in2(N__19943),
            .in3(N__32720),
            .lcout(),
            .ltout(\ALU.N_708_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC8CO3_9_LC_5_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIC8CO3_9_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC8CO3_9_LC_5_11_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIC8CO3_9_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__35230),
            .in2(N__20171),
            .in3(N__20165),
            .lcout(\ALU.aluOut_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIKKOA1_9_LC_5_11_4 .C_ON=1'b0;
    defparam \ALU.f_RNIKKOA1_9_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIKKOA1_9_LC_5_11_4 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \ALU.f_RNIKKOA1_9_LC_5_11_4  (
            .in0(N__28160),
            .in1(N__28133),
            .in2(N__36004),
            .in3(N__35897),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI79CK1_9_LC_5_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNI79CK1_9_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI79CK1_9_LC_5_11_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI79CK1_9_LC_5_11_5  (
            .in0(N__35367),
            .in1(N__32839),
            .in2(N__20168),
            .in3(N__32797),
            .lcout(\ALU.N_756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHBIK1_4_LC_5_12_0 .C_ON=1'b0;
    defparam \ALU.d_RNIHBIK1_4_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHBIK1_4_LC_5_12_0 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.d_RNIHBIK1_4_LC_5_12_0  (
            .in0(N__27287),
            .in1(N__36542),
            .in2(N__35754),
            .in3(N__28997),
            .lcout(),
            .ltout(\ALU.N_751_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHB2E3_4_LC_5_12_1 .C_ON=1'b0;
    defparam \ALU.d_RNIHB2E3_4_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHB2E3_4_LC_5_12_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.d_RNIHB2E3_4_LC_5_12_1  (
            .in0(N__35232),
            .in1(_gnd_net_),
            .in2(N__20159),
            .in3(N__20156),
            .lcout(\ALU.aluOut_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNISKML1_4_LC_5_12_2 .C_ON=1'b0;
    defparam \ALU.g_RNISKML1_4_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNISKML1_4_LC_5_12_2 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.g_RNISKML1_4_LC_5_12_2  (
            .in0(N__26975),
            .in1(N__31862),
            .in2(N__35753),
            .in3(N__29051),
            .lcout(\ALU.N_703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8MG97_5_LC_5_12_3 .C_ON=1'b0;
    defparam \ALU.d_RNI8MG97_5_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8MG97_5_LC_5_12_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.d_RNI8MG97_5_LC_5_12_3  (
            .in0(N__43762),
            .in1(N__40427),
            .in2(N__39139),
            .in3(N__42821),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI609EE_6_LC_5_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNI609EE_6_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI609EE_6_LC_5_12_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \ALU.d_RNI609EE_6_LC_5_12_4  (
            .in0(N__46657),
            .in1(N__46837),
            .in2(N__20150),
            .in3(N__39105),
            .lcout(\ALU.N_472 ),
            .ltout(\ALU.N_472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6EKGV_6_LC_5_12_5 .C_ON=1'b0;
    defparam \ALU.d_RNI6EKGV_6_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6EKGV_6_LC_5_12_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNI6EKGV_6_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__38743),
            .in2(N__20135),
            .in3(N__20132),
            .lcout(\ALU.N_532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_N_1700_i_LC_5_12_7 .C_ON=1'b0;
    defparam \ALU.mult_N_1700_i_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_N_1700_i_LC_5_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ALU.mult_N_1700_i_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38178),
            .lcout(\ALU.N_1700_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNI81NL1_7_LC_5_13_0 .C_ON=1'b0;
    defparam \ALU.g_RNI81NL1_7_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNI81NL1_7_LC_5_13_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.g_RNI81NL1_7_LC_5_13_0  (
            .in0(N__31814),
            .in1(N__31694),
            .in2(N__35738),
            .in3(N__21599),
            .lcout(),
            .ltout(\ALU.N_706_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBDSD3_7_LC_5_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIBDSD3_7_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBDSD3_7_LC_5_13_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIBDSD3_7_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__35220),
            .in2(N__20213),
            .in3(N__20210),
            .lcout(\ALU.aluOut_7 ),
            .ltout(\ALU.aluOut_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIE5297_6_LC_5_13_2 .C_ON=1'b0;
    defparam \ALU.d_RNIE5297_6_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIE5297_6_LC_5_13_2 .LUT_INIT=16'b0111000000100000;
    LogicCell40 \ALU.d_RNIE5297_6_LC_5_13_2  (
            .in0(N__26595),
            .in1(N__26280),
            .in2(N__20204),
            .in3(N__26711),
            .lcout(\ALU.a7_b_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIP6PD3_1_LC_5_13_3 .C_ON=1'b0;
    defparam \ALU.d_RNIP6PD3_1_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIP6PD3_1_LC_5_13_3 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ALU.d_RNIP6PD3_1_LC_5_13_3  (
            .in0(N__25169),
            .in1(N__23336),
            .in2(_gnd_net_),
            .in3(N__23290),
            .lcout(\ALU.N_249_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI64QK7_4_LC_5_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNI64QK7_4_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI64QK7_4_LC_5_13_4 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNI64QK7_4_LC_5_13_4  (
            .in0(N__23485),
            .in1(N__23566),
            .in2(N__26626),
            .in3(N__37894),
            .lcout(\ALU.a0_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIP0RR6_3_LC_5_13_7 .C_ON=1'b0;
    defparam \ALU.d_RNIP0RR6_3_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIP0RR6_3_LC_5_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIP0RR6_3_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__41926),
            .in2(_gnd_net_),
            .in3(N__38177),
            .lcout(\ALU.a3_b_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIAE1U4_11_LC_5_14_0 .C_ON=1'b0;
    defparam \ALU.c_RNIAE1U4_11_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIAE1U4_11_LC_5_14_0 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \ALU.c_RNIAE1U4_11_LC_5_14_0  (
            .in0(N__24926),
            .in1(N__39382),
            .in2(N__20186),
            .in3(N__29309),
            .lcout(\ALU.N_272_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_89_0_LC_5_14_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_89_0_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_89_0_LC_5_14_1 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_89_0_LC_5_14_1  (
            .in0(N__38176),
            .in1(N__40098),
            .in2(N__37156),
            .in3(N__46658),
            .lcout(\ALU.madd_89_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_20_0_LC_5_14_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_20_0_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_20_0_LC_5_14_2 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_20_0_LC_5_14_2  (
            .in0(N__41883),
            .in1(N__37098),
            .in2(N__38273),
            .in3(N__40277),
            .lcout(),
            .ltout(\ALU.madd_20_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_20_LC_5_14_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_20_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_20_LC_5_14_3 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \ALU.mult_madd_20_LC_5_14_3  (
            .in0(N__42823),
            .in1(_gnd_net_),
            .in2(N__20306),
            .in3(N__37627),
            .lcout(\ALU.madd_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC6QK6_5_LC_5_14_4 .C_ON=1'b0;
    defparam \ALU.d_RNIC6QK6_5_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC6QK6_5_LC_5_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIC6QK6_5_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__40276),
            .in2(_gnd_net_),
            .in3(N__37094),
            .lcout(\ALU.a5_b_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m4_LC_5_14_5 .C_ON=1'b0;
    defparam \ALU.m4_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.m4_LC_5_14_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ALU.m4_LC_5_14_5  (
            .in0(N__30196),
            .in1(N__25215),
            .in2(_gnd_net_),
            .in3(N__29735),
            .lcout(\ALU.N_5_0 ),
            .ltout(\ALU.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3GPD3_2_LC_5_14_6 .C_ON=1'b0;
    defparam \ALU.d_RNI3GPD3_2_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3GPD3_2_LC_5_14_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ALU.d_RNI3GPD3_2_LC_5_14_6  (
            .in0(N__25170),
            .in1(N__20291),
            .in2(N__20252),
            .in3(N__28726),
            .lcout(\ALU.N_240_0 ),
            .ltout(\ALU.N_240_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_24_0_tz_LC_5_14_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_24_0_tz_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_24_0_tz_LC_5_14_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ALU.mult_madd_24_0_tz_LC_5_14_7  (
            .in0(N__42822),
            .in1(N__41882),
            .in2(N__20249),
            .in3(N__37626),
            .lcout(\ALU.madd_24_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_66_LC_5_15_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_66_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_66_LC_5_15_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALU.mult_madd_66_LC_5_15_0  (
            .in0(N__36938),
            .in1(N__41704),
            .in2(N__42969),
            .in3(N__28068),
            .lcout(\ALU.madd_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_8_0_LC_5_15_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_8_0_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_8_0_LC_5_15_1 .LUT_INIT=16'b0111100010001000;
    LogicCell40 \ALU.mult_madd_8_0_LC_5_15_1  (
            .in0(N__38192),
            .in1(N__42916),
            .in2(N__37158),
            .in3(N__36940),
            .lcout(\ALU.madd_8_0 ),
            .ltout(\ALU.madd_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_18_LC_5_15_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_18_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_18_LC_5_15_2 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ALU.mult_madd_18_LC_5_15_2  (
            .in0(N__37656),
            .in1(N__20228),
            .in2(N__20216),
            .in3(N__41973),
            .lcout(\ALU.madd_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_128_0_tz_LC_5_15_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_128_0_tz_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_128_0_tz_LC_5_15_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ALU.mult_madd_128_0_tz_LC_5_15_3  (
            .in0(N__40044),
            .in1(N__46839),
            .in2(N__37157),
            .in3(N__37654),
            .lcout(\ALU.madd_128_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_68_0_tz_LC_5_15_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_68_0_tz_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_68_0_tz_LC_5_15_4 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \ALU.mult_madd_68_0_tz_LC_5_15_4  (
            .in0(N__36939),
            .in1(N__41705),
            .in2(N__42970),
            .in3(N__28069),
            .lcout(\ALU.madd_68_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRALR6_7_LC_5_15_5 .C_ON=1'b0;
    defparam \ALU.d_RNIRALR6_7_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRALR6_7_LC_5_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALU.d_RNIRALR6_7_LC_5_15_5  (
            .in0(N__38191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46838),
            .lcout(\ALU.a7_b_0 ),
            .ltout(\ALU.a7_b_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_59_LC_5_15_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_59_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_59_LC_5_15_6 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \ALU.mult_madd_59_LC_5_15_6  (
            .in0(N__37655),
            .in1(N__46638),
            .in2(N__20417),
            .in3(N__24526),
            .lcout(\ALU.madd_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_5_LC_5_15_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_5_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_5_LC_5_15_7 .LUT_INIT=16'b0010001011010010;
    LogicCell40 \ALU.mult_madd_484_5_LC_5_15_7  (
            .in0(N__40045),
            .in1(N__47067),
            .in2(N__39852),
            .in3(N__46444),
            .lcout(\ALU.madd_484_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_26_LC_5_16_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_26_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_26_LC_5_16_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ALU.mult_g0_26_LC_5_16_0  (
            .in0(N__40046),
            .in1(N__46876),
            .in2(N__37203),
            .in3(N__37657),
            .lcout(\ALU.madd_128_0_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_104_LC_5_16_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_104_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_104_LC_5_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_104_LC_5_16_1  (
            .in0(N__20573),
            .in1(N__20588),
            .in2(N__24515),
            .in3(N__20594),
            .lcout(\ALU.madd_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_149_LC_5_16_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_149_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_149_LC_5_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_149_LC_5_16_2  (
            .in0(N__20541),
            .in1(N__21948),
            .in2(_gnd_net_),
            .in3(N__20554),
            .lcout(\ALU.madd_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_128_0_LC_5_16_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_128_0_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_128_0_LC_5_16_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ALU.mult_madd_128_0_LC_5_16_3  (
            .in0(N__38272),
            .in1(N__39825),
            .in2(_gnd_net_),
            .in3(N__20336),
            .lcout(\ALU.madd_128_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_m3_LC_5_16_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_m3_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_m3_LC_5_16_4 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \ALU.mult_madd_m3_LC_5_16_4  (
            .in0(N__20543),
            .in1(N__21950),
            .in2(_gnd_net_),
            .in3(N__20555),
            .lcout(\ALU.madd_N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_68_LC_5_16_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_68_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_68_LC_5_16_5 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \ALU.mult_madd_68_LC_5_16_5  (
            .in0(N__41993),
            .in1(N__20606),
            .in2(N__42698),
            .in3(N__20600),
            .lcout(\ALU.madd_68 ),
            .ltout(\ALU.madd_68_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_108_LC_5_16_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_108_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_108_LC_5_16_6 .LUT_INIT=16'b1101010011101000;
    LogicCell40 \ALU.mult_madd_108_LC_5_16_6  (
            .in0(N__20587),
            .in1(N__24511),
            .in2(N__20576),
            .in3(N__20572),
            .lcout(\ALU.madd_108 ),
            .ltout(\ALU.madd_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_153_LC_5_16_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_153_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_153_LC_5_16_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \ALU.mult_madd_153_LC_5_16_7  (
            .in0(N__21949),
            .in1(_gnd_net_),
            .in2(N__20546),
            .in3(N__20542),
            .lcout(\ALU.madd_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXready_LC_6_1_0 .C_ON=1'b0;
    defparam \FTDI.RXready_LC_6_1_0 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXready_LC_6_1_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \FTDI.RXready_LC_6_1_0  (
            .in0(N__24767),
            .in1(N__20668),
            .in2(N__24661),
            .in3(N__24742),
            .lcout(RXready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXreadyC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.gap_RNI29TH_2_LC_6_1_1 .C_ON=1'b0;
    defparam \FTDI.gap_RNI29TH_2_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.gap_RNI29TH_2_LC_6_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FTDI.gap_RNI29TH_2_LC_6_1_1  (
            .in0(_gnd_net_),
            .in1(N__29249),
            .in2(_gnd_net_),
            .in3(N__24652),
            .lcout(\FTDI.N_201_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_2_LC_6_1_2 .C_ON=1'b0;
    defparam \FTDI.RXstate_2_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_2_LC_6_1_2 .LUT_INIT=16'b0110000010100000;
    LogicCell40 \FTDI.RXstate_2_LC_6_1_2  (
            .in0(N__24768),
            .in1(N__20669),
            .in2(N__24662),
            .in3(N__24743),
            .lcout(\FTDI.RXstateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.RXreadyC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m681_1_LC_6_1_3 .C_ON=1'b0;
    defparam \ALU.m681_1_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m681_1_LC_6_1_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALU.m681_1_LC_6_1_3  (
            .in0(N__43090),
            .in1(N__20479),
            .in2(N__48054),
            .in3(N__44028),
            .lcout(),
            .ltout(\ALU.m681Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m681_LC_6_1_4 .C_ON=1'b0;
    defparam \ALU.m681_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m681_LC_6_1_4 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \ALU.m681_LC_6_1_4  (
            .in0(N__33173),
            .in1(N__45699),
            .in2(N__20462),
            .in3(N__26649),
            .lcout(\ALU.N_730_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m57_LC_6_1_5 .C_ON=1'b0;
    defparam \ALU.m57_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \ALU.m57_LC_6_1_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.m57_LC_6_1_5  (
            .in0(_gnd_net_),
            .in1(N__30285),
            .in2(_gnd_net_),
            .in3(N__21883),
            .lcout(\ALU.N_58_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNI67DS1_0_LC_6_1_6 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNI67DS1_0_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNI67DS1_0_LC_6_1_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \FTDI.RXstate_RNI67DS1_0_LC_6_1_6  (
            .in0(N__24766),
            .in1(N__24741),
            .in2(N__24660),
            .in3(N__24688),
            .lcout(\FTDI.gap8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNIV5TH_0_LC_6_1_7 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNIV5TH_0_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNIV5TH_0_LC_6_1_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \FTDI.RXstate_RNIV5TH_0_LC_6_1_7  (
            .in0(N__24689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29250),
            .lcout(\FTDI.N_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEN0V7_0_LC_6_2_0 .C_ON=1'b0;
    defparam \ALU.d_RNIEN0V7_0_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEN0V7_0_LC_6_2_0 .LUT_INIT=16'b0000111101011010;
    LogicCell40 \ALU.d_RNIEN0V7_0_LC_6_2_0  (
            .in0(N__38306),
            .in1(_gnd_net_),
            .in2(N__38045),
            .in3(N__43859),
            .lcout(\ALU.a_15_m1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID9RV5_0_LC_6_2_1 .C_ON=1'b0;
    defparam \ALU.d_RNID9RV5_0_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID9RV5_0_LC_6_2_1 .LUT_INIT=16'b0010011100100010;
    LogicCell40 \ALU.d_RNID9RV5_0_LC_6_2_1  (
            .in0(N__44037),
            .in1(N__47230),
            .in2(N__44524),
            .in3(N__20755),
            .lcout(),
            .ltout(\ALU.a_15_m4_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINPK3M_0_LC_6_2_2 .C_ON=1'b0;
    defparam \ALU.d_RNINPK3M_0_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINPK3M_0_LC_6_2_2 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \ALU.d_RNINPK3M_0_LC_6_2_2  (
            .in0(N__44159),
            .in1(N__20660),
            .in2(N__20654),
            .in3(N__20624),
            .lcout(),
            .ltout(\ALU.a_15_m4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITQOAQ2_0_LC_6_2_3 .C_ON=1'b0;
    defparam \ALU.d_RNITQOAQ2_0_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITQOAQ2_0_LC_6_2_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNITQOAQ2_0_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(N__46310),
            .in2(N__20651),
            .in3(N__20648),
            .lcout(\ALU.a_15_m5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m4_bm_1_8_LC_6_2_4 .C_ON=1'b0;
    defparam \ALU.a_15_m4_bm_1_8_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m4_bm_1_8_LC_6_2_4 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \ALU.a_15_m4_bm_1_8_LC_6_2_4  (
            .in0(N__47229),
            .in1(_gnd_net_),
            .in2(N__43881),
            .in3(N__24579),
            .lcout(\ALU.a_15_m4_bm_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITTVL7_0_LC_6_2_5 .C_ON=1'b0;
    defparam \ALU.d_RNITTVL7_0_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITTVL7_0_LC_6_2_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \ALU.d_RNITTVL7_0_LC_6_2_5  (
            .in0(N__24580),
            .in1(N__38022),
            .in2(_gnd_net_),
            .in3(N__38307),
            .lcout(\ALU.a_15_m0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_0_LC_6_2_6 .C_ON=1'b0;
    defparam \CONTROL.aluParams_0_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluParams_0_LC_6_2_6 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \CONTROL.aluParams_0_LC_6_2_6  (
            .in0(N__22137),
            .in1(N__20618),
            .in2(_gnd_net_),
            .in3(N__43583),
            .lcout(aluParams_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47623),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPD997_6_LC_6_2_7 .C_ON=1'b0;
    defparam \ALU.d_RNIPD997_6_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPD997_6_LC_6_2_7 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.d_RNIPD997_6_LC_6_2_7  (
            .in0(N__43582),
            .in1(N__40424),
            .in2(N__38968),
            .in3(N__46734),
            .lcout(\ALU.rshift_3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI5PUHV_10_LC_6_3_0 .C_ON=1'b0;
    defparam \ALU.c_RNI5PUHV_10_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI5PUHV_10_LC_6_3_0 .LUT_INIT=16'b0000100000111011;
    LogicCell40 \ALU.c_RNI5PUHV_10_LC_6_3_0  (
            .in0(N__20702),
            .in1(N__43139),
            .in2(N__44449),
            .in3(N__20735),
            .lcout(\ALU.a_15_m3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFL4K8_11_LC_6_3_1 .C_ON=1'b0;
    defparam \ALU.c_RNIFL4K8_11_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFL4K8_11_LC_6_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIFL4K8_11_LC_6_3_1  (
            .in0(N__43674),
            .in1(N__39385),
            .in2(_gnd_net_),
            .in3(N__27589),
            .lcout(\ALU.N_461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3BB3U_5_LC_6_3_2 .C_ON=1'b0;
    defparam \ALU.d_RNI3BB3U_5_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3BB3U_5_LC_6_3_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNI3BB3U_5_LC_6_3_2  (
            .in0(N__38559),
            .in1(N__24818),
            .in2(_gnd_net_),
            .in3(N__20714),
            .lcout(),
            .ltout(\ALU.N_530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIP8ITN1_5_LC_6_3_3 .C_ON=1'b0;
    defparam \ALU.d_RNIP8ITN1_5_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIP8ITN1_5_LC_6_3_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIP8ITN1_5_LC_6_3_3  (
            .in0(_gnd_net_),
            .in1(N__44393),
            .in2(N__20705),
            .in3(N__20701),
            .lcout(),
            .ltout(\ALU.d_RNIP8ITN1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFHQSS1_2_LC_6_3_4 .C_ON=1'b0;
    defparam \ALU.d_RNIFHQSS1_2_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFHQSS1_2_LC_6_3_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIFHQSS1_2_LC_6_3_4  (
            .in0(_gnd_net_),
            .in1(N__43140),
            .in2(N__20693),
            .in3(N__20690),
            .lcout(),
            .ltout(\ALU.a_15_m3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDVDOJ2_2_LC_6_3_5 .C_ON=1'b0;
    defparam \ALU.d_RNIDVDOJ2_2_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDVDOJ2_2_LC_6_3_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIDVDOJ2_2_LC_6_3_5  (
            .in0(_gnd_net_),
            .in1(N__46311),
            .in2(N__20681),
            .in3(N__20675),
            .lcout(\ALU.a_15_m5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIE937B_0_LC_6_3_6 .C_ON=1'b0;
    defparam \ALU.d_RNIE937B_0_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIE937B_0_LC_6_3_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.d_RNIE937B_0_LC_6_3_6  (
            .in0(N__38560),
            .in1(N__44422),
            .in2(_gnd_net_),
            .in3(N__39180),
            .lcout(),
            .ltout(\ALU.d_RNIE937BZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVM1UL_2_LC_6_3_7 .C_ON=1'b0;
    defparam \ALU.d_RNIVM1UL_2_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVM1UL_2_LC_6_3_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIVM1UL_2_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(N__44139),
            .in2(N__20678),
            .in3(N__24830),
            .lcout(\ALU.a_15_m4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI75NNF_6_LC_6_4_0 .C_ON=1'b0;
    defparam \ALU.d_RNI75NNF_6_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI75NNF_6_LC_6_4_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.d_RNI75NNF_6_LC_6_4_0  (
            .in0(N__38966),
            .in1(N__22915),
            .in2(N__38603),
            .in3(N__22894),
            .lcout(\ALU.lshift_7_ns_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINVVJ11_13_LC_6_4_1 .C_ON=1'b0;
    defparam \ALU.c_RNINVVJ11_13_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINVVJ11_13_LC_6_4_1 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.c_RNINVVJ11_13_LC_6_4_1  (
            .in0(N__38593),
            .in1(N__20777),
            .in2(N__44492),
            .in3(N__20767),
            .lcout(\ALU.lshift_15_ns_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNII1LGE_5_LC_6_4_2 .C_ON=1'b0;
    defparam \ALU.d_RNII1LGE_5_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNII1LGE_5_LC_6_4_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNII1LGE_5_LC_6_4_2  (
            .in0(N__38967),
            .in1(N__22810),
            .in2(_gnd_net_),
            .in3(N__22895),
            .lcout(\ALU.N_249 ),
            .ltout(\ALU.N_249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIUGCLV_11_LC_6_4_3 .C_ON=1'b0;
    defparam \ALU.c_RNIUGCLV_11_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIUGCLV_11_LC_6_4_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNIUGCLV_11_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(N__38528),
            .in2(N__20771),
            .in3(N__20768),
            .lcout(),
            .ltout(\ALU.c_RNIUGCLVZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILTHAE1_1_LC_6_4_4 .C_ON=1'b0;
    defparam \ALU.d_RNILTHAE1_1_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILTHAE1_1_LC_6_4_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNILTHAE1_1_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(N__44443),
            .in2(N__20759),
            .in3(N__22823),
            .lcout(\ALU.lshift_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEUKR11_0_LC_6_4_5 .C_ON=1'b0;
    defparam \ALU.d_RNIEUKR11_0_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEUKR11_0_LC_6_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIEUKR11_0_LC_6_4_5  (
            .in0(N__44442),
            .in1(N__20756),
            .in2(_gnd_net_),
            .in3(N__20744),
            .lcout(\ALU.d_RNIEUKR11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI83IG7_3_LC_6_4_6 .C_ON=1'b0;
    defparam \ALU.d_RNI83IG7_3_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI83IG7_3_LC_6_4_6 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.d_RNI83IG7_3_LC_6_4_6  (
            .in0(N__43620),
            .in1(N__41995),
            .in2(N__42997),
            .in3(N__39141),
            .lcout(),
            .ltout(\ALU.lshift_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICH0SD_1_LC_6_4_7 .C_ON=1'b0;
    defparam \ALU.d_RNICH0SD_1_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICH0SD_1_LC_6_4_7 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.d_RNICH0SD_1_LC_6_4_7  (
            .in0(N__36957),
            .in1(N__38965),
            .in2(N__20738),
            .in3(N__37426),
            .lcout(\ALU.N_246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFL4K8_0_11_LC_6_5_0 .C_ON=1'b0;
    defparam \ALU.c_RNIFL4K8_0_11_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFL4K8_0_11_LC_6_5_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.c_RNIFL4K8_0_11_LC_6_5_0  (
            .in0(N__27558),
            .in1(N__43586),
            .in2(_gnd_net_),
            .in3(N__39389),
            .lcout(\ALU.N_223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5MUQE_6_LC_6_5_1 .C_ON=1'b0;
    defparam \ALU.d_RNI5MUQE_6_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5MUQE_6_LC_6_5_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNI5MUQE_6_LC_6_5_1  (
            .in0(N__39142),
            .in1(N__20825),
            .in2(_gnd_net_),
            .in3(N__20801),
            .lcout(\ALU.N_250 ),
            .ltout(\ALU.N_250_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNISJ8601_11_LC_6_5_2 .C_ON=1'b0;
    defparam \ALU.c_RNISJ8601_11_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNISJ8601_11_LC_6_5_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.c_RNISJ8601_11_LC_6_5_2  (
            .in0(N__38722),
            .in1(_gnd_net_),
            .in2(N__20810),
            .in3(N__20807),
            .lcout(\ALU.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIVUE24_0_LC_6_5_3 .C_ON=1'b0;
    defparam \ALU.d_RNIVUE24_0_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIVUE24_0_LC_6_5_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.d_RNIVUE24_0_LC_6_5_3  (
            .in0(N__43587),
            .in1(N__39144),
            .in2(_gnd_net_),
            .in3(N__37962),
            .lcout(\ALU.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIK8CGE_5_LC_6_5_4 .C_ON=1'b0;
    defparam \ALU.d_RNIK8CGE_5_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIK8CGE_5_LC_6_5_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNIK8CGE_5_LC_6_5_4  (
            .in0(N__39145),
            .in1(N__22803),
            .in2(_gnd_net_),
            .in3(N__23043),
            .lcout(\ALU.N_247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8K807_6_LC_6_5_5 .C_ON=1'b0;
    defparam \ALU.d_RNI8K807_6_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8K807_6_LC_6_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNI8K807_6_LC_6_5_5  (
            .in0(N__43585),
            .in1(N__40402),
            .in2(_gnd_net_),
            .in3(N__46720),
            .lcout(\ALU.N_218 ),
            .ltout(\ALU.N_218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGNQGE_3_LC_6_5_6 .C_ON=1'b0;
    defparam \ALU.d_RNIGNQGE_3_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGNQGE_3_LC_6_5_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIGNQGE_3_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(N__39143),
            .in2(N__20795),
            .in3(N__23024),
            .lcout(\ALU.N_361 ),
            .ltout(\ALU.N_361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1GH4V_7_LC_6_5_7 .C_ON=1'b0;
    defparam \ALU.d_RNI1GH4V_7_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1GH4V_7_LC_6_5_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNI1GH4V_7_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(N__38723),
            .in2(N__20792),
            .in3(N__20788),
            .lcout(\ALU.d_RNI1GH4VZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_28_LC_6_6_0.C_ON=1'b0;
    defparam testWord_28_LC_6_6_0.SEQ_MODE=4'b1000;
    defparam testWord_28_LC_6_6_0.LUT_INIT=16'b1011100011110000;
    LogicCell40 testWord_28_LC_6_6_0 (
            .in0(N__32293),
            .in1(N__41159),
            .in2(N__20972),
            .in3(N__41474),
            .lcout(ctrlOut_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47650),
            .ce(N__41060),
            .sr(_gnd_net_));
    defparam \ALU.m270_ns_1_LC_6_6_1 .C_ON=1'b0;
    defparam \ALU.m270_ns_1_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.m270_ns_1_LC_6_6_1 .LUT_INIT=16'b0001000110000000;
    LogicCell40 \ALU.m270_ns_1_LC_6_6_1  (
            .in0(N__30193),
            .in1(N__26637),
            .in2(N__20971),
            .in3(N__29692),
            .lcout(),
            .ltout(\ALU.m270_nsZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNILQ2U4_12_LC_6_6_2 .C_ON=1'b0;
    defparam \ALU.c_RNILQ2U4_12_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNILQ2U4_12_LC_6_6_2 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.c_RNILQ2U4_12_LC_6_6_2  (
            .in0(N__25348),
            .in1(N__20966),
            .in2(N__20975),
            .in3(N__29403),
            .lcout(\ALU.N_271_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m178_LC_6_6_3 .C_ON=1'b0;
    defparam \ALU.m178_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.m178_LC_6_6_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ALU.m178_LC_6_6_3  (
            .in0(N__30192),
            .in1(N__25139),
            .in2(N__20970),
            .in3(N__29691),
            .lcout(\ALU.N_179_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIM75G5_15_LC_6_6_4 .C_ON=1'b0;
    defparam \ALU.d_RNIM75G5_15_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIM75G5_15_LC_6_6_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ALU.d_RNIM75G5_15_LC_6_6_4  (
            .in0(N__24149),
            .in1(N__29402),
            .in2(N__20945),
            .in3(N__31322),
            .lcout(\ALU.N_7_0 ),
            .ltout(\ALU.N_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_0_LC_6_6_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_0_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_0_LC_6_6_5 .LUT_INIT=16'b0110101011000000;
    LogicCell40 \ALU.mult_madd_484_0_LC_6_6_5  (
            .in0(N__41976),
            .in1(N__37961),
            .in2(N__20921),
            .in3(N__40826),
            .lcout(\ALU.madd_484_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4K3G5_12_LC_6_6_6 .C_ON=1'b0;
    defparam \ALU.d_RNI4K3G5_12_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4K3G5_12_LC_6_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNI4K3G5_12_LC_6_6_6  (
            .in0(N__24148),
            .in1(N__20894),
            .in2(_gnd_net_),
            .in3(N__25442),
            .lcout(\ALU.N_180_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_13_LC_6_7_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_13_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_13_LC_6_7_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \ALU.a_15_m2_ns_1_13_LC_6_7_0  (
            .in0(N__47233),
            .in1(N__24588),
            .in2(_gnd_net_),
            .in3(N__43861),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNID22SC_13_LC_6_7_1 .C_ON=1'b0;
    defparam \ALU.c_RNID22SC_13_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNID22SC_13_LC_6_7_1 .LUT_INIT=16'b1001010100101011;
    LogicCell40 \ALU.c_RNID22SC_13_LC_6_7_1  (
            .in0(N__40746),
            .in1(N__24969),
            .in2(N__20873),
            .in3(N__47234),
            .lcout(\ALU.a_15_m2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m714_LC_6_7_2 .C_ON=1'b0;
    defparam \ALU.m714_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.m714_LC_6_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.m714_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__44133),
            .in2(_gnd_net_),
            .in3(N__43584),
            .lcout(\ALU.log_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_3_LC_6_7_3 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_3_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_3_LC_6_7_3 .LUT_INIT=16'b1011010001000100;
    LogicCell40 \ALU.mult_madd_484_3_LC_6_7_3  (
            .in0(N__22002),
            .in1(N__46729),
            .in2(N__40764),
            .in3(N__37231),
            .lcout(\ALU.madd_484_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIG6C84_9_LC_6_7_4 .C_ON=1'b0;
    defparam \ALU.d_RNIG6C84_9_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIG6C84_9_LC_6_7_4 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \ALU.d_RNIG6C84_9_LC_6_7_4  (
            .in0(N__32990),
            .in1(N__28109),
            .in2(N__24449),
            .in3(N__32849),
            .lcout(\ALU.operand2_9 ),
            .ltout(\ALU.operand2_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHIKU4_9_LC_6_7_5 .C_ON=1'b0;
    defparam \ALU.d_RNIHIKU4_9_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHIKU4_9_LC_6_7_5 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \ALU.d_RNIHIKU4_9_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__21057),
            .in2(N__21032),
            .in3(N__24144),
            .lcout(\ALU.N_207_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_9_LC_6_7_6 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_9_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_9_LC_6_7_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \ALU.a_15_m2_ns_1_9_LC_6_7_6  (
            .in0(N__47231),
            .in1(N__24587),
            .in2(_gnd_net_),
            .in3(N__43860),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6904C_9_LC_6_7_7 .C_ON=1'b0;
    defparam \ALU.d_RNI6904C_9_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6904C_9_LC_6_7_7 .LUT_INIT=16'b1001001101001101;
    LogicCell40 \ALU.d_RNI6904C_9_LC_6_7_7  (
            .in0(N__22003),
            .in1(N__47232),
            .in2(N__21029),
            .in3(N__39832),
            .lcout(\ALU.a_15_m2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_13_LC_6_8_0 .C_ON=1'b0;
    defparam \ALU.h_13_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_13_LC_6_8_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.h_13_LC_6_8_0  (
            .in0(N__48598),
            .in1(N__33940),
            .in2(N__45873),
            .in3(N__33881),
            .lcout(\ALU.hZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(N__45489),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO7LU_13_LC_6_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNIO7LU_13_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO7LU_13_LC_6_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIO7LU_13_LC_6_8_1  (
            .in0(N__45334),
            .in1(N__35446),
            .in2(_gnd_net_),
            .in3(N__35435),
            .lcout(),
            .ltout(\ALU.d_RNIO7LUZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8DRP4_0_13_LC_6_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNI8DRP4_0_13_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8DRP4_0_13_LC_6_8_2 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \ALU.d_RNI8DRP4_0_13_LC_6_8_2  (
            .in0(N__28439),
            .in1(N__32994),
            .in2(N__21026),
            .in3(N__31103),
            .lcout(\ALU.operand2_13 ),
            .ltout(\ALU.operand2_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDT3G5_13_LC_6_8_3 .C_ON=1'b0;
    defparam \ALU.d_RNIDT3G5_13_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDT3G5_13_LC_6_8_3 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \ALU.d_RNIDT3G5_13_LC_6_8_3  (
            .in0(N__25053),
            .in1(_gnd_net_),
            .in2(N__21023),
            .in3(N__24153),
            .lcout(\ALU.N_177_0 ),
            .ltout(\ALU.N_177_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_2_LC_6_8_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_2_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_2_LC_6_8_4 .LUT_INIT=16'b0000110010100110;
    LogicCell40 \ALU.mult_madd_484_2_LC_6_8_4  (
            .in0(N__37376),
            .in1(N__36878),
            .in2(N__21020),
            .in3(N__21313),
            .lcout(),
            .ltout(\ALU.madd_484_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_12_LC_6_8_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_12_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_12_LC_6_8_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \ALU.mult_madd_484_12_LC_6_8_5  (
            .in0(N__21017),
            .in1(N__21008),
            .in2(N__20996),
            .in3(N__20993),
            .lcout(\ALU.madd_484_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7TLM8_0_LC_6_9_0 .C_ON=1'b1;
    defparam \ALU.d_RNI7TLM8_0_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7TLM8_0_LC_6_9_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \ALU.d_RNI7TLM8_0_LC_6_9_0  (
            .in0(N__39440),
            .in1(N__37968),
            .in2(N__36325),
            .in3(_gnd_net_),
            .lcout(\ALU.a0_b_11 ),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\ALU.un2_addsub_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_0_c_RNI5MA0E_LC_6_9_1 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_0_c_RNI5MA0E_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_0_c_RNI5MA0E_LC_6_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_0_c_RNI5MA0E_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__23351),
            .in2(N__23279),
            .in3(N__21215),
            .lcout(\ALU.un2_addsub_cry_0_c_RNI5MA0EZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_0 ),
            .carryout(\ALU.un2_addsub_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_1_c_RNI966GE_LC_6_9_2 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_1_c_RNI966GE_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_1_c_RNI966GE_LC_6_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_1_c_RNI966GE_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__21212),
            .in2(N__21197),
            .in3(N__21179),
            .lcout(\ALU.un2_addsub_cry_1_c_RNI966GEZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_1 ),
            .carryout(\ALU.un2_addsub_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_2_c_RNI5IV5F_LC_6_9_3 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_2_c_RNI5IV5F_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_2_c_RNI5IV5F_LC_6_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_2_c_RNI5IV5F_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__41719),
            .in2(N__23846),
            .in3(N__21176),
            .lcout(\ALU.un2_addsub_cry_2_c_RNI5IV5FZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_2 ),
            .carryout(\ALU.un2_addsub_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_3_c_RNIOGGJG_LC_6_9_4 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_3_c_RNIOGGJG_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_3_c_RNIOGGJG_LC_6_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_3_c_RNIOGGJG_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__42683),
            .in2(N__21800),
            .in3(N__21173),
            .lcout(\ALU.un2_addsub_cry_3_c_RNIOGGJGZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_3 ),
            .carryout(\ALU.un2_addsub_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_4_c_RNI284VE_LC_6_9_5 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_4_c_RNI284VE_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_4_c_RNI284VE_LC_6_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_4_c_RNI284VE_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__28090),
            .in2(N__21170),
            .in3(N__21152),
            .lcout(\ALU.un2_addsub_cry_4_c_RNI284VEZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_4 ),
            .carryout(\ALU.un2_addsub_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_5_c_RNIL7IGF_LC_6_9_6 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_5_c_RNIL7IGF_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_5_c_RNIL7IGF_LC_6_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_5_c_RNIL7IGF_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(N__46474),
            .in2(N__21149),
            .in3(N__21128),
            .lcout(\ALU.un2_addsub_cry_5_c_RNIL7IGFZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_5 ),
            .carryout(\ALU.un2_addsub_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_6_c_RNIL4LMI_LC_6_9_7 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_6_c_RNIL4LMI_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_6_c_RNIL4LMI_LC_6_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_6_c_RNIL4LMI_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(N__47101),
            .in2(N__21125),
            .in3(N__21101),
            .lcout(\ALU.un2_addsub_cry_6_c_RNIL4LMIZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_6 ),
            .carryout(\ALU.un2_addsub_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_7_c_RNIL8JHG_LC_6_10_0 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_7_c_RNIL8JHG_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_7_c_RNIL8JHG_LC_6_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_7_c_RNIL8JHG_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__21471),
            .in2(N__21404),
            .in3(N__21386),
            .lcout(\ALU.un2_addsub_cry_7_c_RNIL8JHGZ0 ),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\ALU.un2_addsub_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_8_c_RNIKR81J_LC_6_10_1 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_8_c_RNIKR81J_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_8_c_RNIKR81J_LC_6_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_8_c_RNIKR81J_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__22057),
            .in2(N__21383),
            .in3(N__21368),
            .lcout(\ALU.un2_addsub_cry_8_c_RNIKR81JZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_8 ),
            .carryout(\ALU.un2_addsub_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_9_c_RNIVCOFA_LC_6_10_2 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_9_c_RNIVCOFA_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_9_c_RNIVCOFA_LC_6_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_9_c_RNIVCOFA_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__27511),
            .in2(N__21365),
            .in3(N__21347),
            .lcout(\ALU.un2_addsub_cry_9_c_RNIVCOFAZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_9 ),
            .carryout(\ALU.un2_addsub_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_10_c_RNIUS1OJ_LC_6_10_3 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_10_c_RNIUS1OJ_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_10_c_RNIUS1OJ_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_10_c_RNIUS1OJ_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__25571),
            .in2(N__24848),
            .in3(N__21344),
            .lcout(\ALU.un2_addsub_cry_10_c_RNIUS1OJZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_10 ),
            .carryout(\ALU.un2_addsub_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_11_c_RNII7OF9_LC_6_10_4 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_11_c_RNII7OF9_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_11_c_RNII7OF9_LC_6_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_11_c_RNII7OF9_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__25379),
            .in2(N__21341),
            .in3(N__21320),
            .lcout(\ALU.un2_addsub_cry_11_c_RNII7OFZ0Z9 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_11 ),
            .carryout(\ALU.un2_addsub_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_12_c_RNIUL1GK_LC_6_10_5 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_12_c_RNIUL1GK_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_12_c_RNIUL1GK_LC_6_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_12_c_RNIUL1GK_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__24973),
            .in2(N__24947),
            .in3(N__21317),
            .lcout(\ALU.un2_addsub_cry_12_c_RNIUL1GKZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_12 ),
            .carryout(\ALU.un2_addsub_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_13_c_RNINVE5K_LC_6_10_6 .C_ON=1'b1;
    defparam \ALU.un2_addsub_cry_13_c_RNINVE5K_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_13_c_RNINVE5K_LC_6_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un2_addsub_cry_13_c_RNINVE5K_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__21314),
            .in2(N__21263),
            .in3(N__21245),
            .lcout(\ALU.un2_addsub_cry_13_c_RNINVE5KZ0 ),
            .ltout(),
            .carryin(\ALU.un2_addsub_cry_13 ),
            .carryout(\ALU.un2_addsub_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_14_c_RNINOK69_LC_6_10_7 .C_ON=1'b0;
    defparam \ALU.un2_addsub_cry_14_c_RNINOK69_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_14_c_RNINOK69_LC_6_10_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \ALU.un2_addsub_cry_14_c_RNINOK69_LC_6_10_7  (
            .in0(N__32608),
            .in1(N__32675),
            .in2(_gnd_net_),
            .in3(N__21242),
            .lcout(\ALU.un2_addsub_cry_14_c_RNINOKZ0Z69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_10_LC_6_11_0 .C_ON=1'b0;
    defparam \ALU.h_10_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_10_LC_6_11_0 .LUT_INIT=16'b0101010111010001;
    LogicCell40 \ALU.h_10_LC_6_11_0  (
            .in0(N__34326),
            .in1(N__45842),
            .in2(N__34415),
            .in3(N__48251),
            .lcout(\ALU.hZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47679),
            .ce(N__45586),
            .sr(_gnd_net_));
    defparam \ALU.g0_2_1_LC_6_11_1 .C_ON=1'b0;
    defparam \ALU.g0_2_1_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.g0_2_1_LC_6_11_1 .LUT_INIT=16'b0001110111011101;
    LogicCell40 \ALU.g0_2_1_LC_6_11_1  (
            .in0(N__31260),
            .in1(N__25213),
            .in2(N__30216),
            .in3(N__21518),
            .lcout(\ALU.g0_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIPN2P1_10_LC_6_11_2 .C_ON=1'b0;
    defparam \ALU.a_RNIPN2P1_10_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIPN2P1_10_LC_6_11_2 .LUT_INIT=16'b0000110011111010;
    LogicCell40 \ALU.a_RNIPN2P1_10_LC_6_11_2  (
            .in0(N__28600),
            .in1(N__23707),
            .in2(N__34514),
            .in3(N__34814),
            .lcout(),
            .ltout(\ALU.N_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIULHV4_10_LC_6_11_3 .C_ON=1'b0;
    defparam \ALU.a_RNIULHV4_10_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIULHV4_10_LC_6_11_3 .LUT_INIT=16'b0101000011101110;
    LogicCell40 \ALU.a_RNIULHV4_10_LC_6_11_3  (
            .in0(N__25214),
            .in1(N__21500),
            .in2(N__21512),
            .in3(N__21509),
            .lcout(\ALU.N_192_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGNUR_10_LC_6_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNIGNUR_10_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGNUR_10_LC_6_11_4 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \ALU.d_RNIGNUR_10_LC_6_11_4  (
            .in0(N__28422),
            .in1(N__35026),
            .in2(N__24427),
            .in3(N__34901),
            .lcout(),
            .ltout(\ALU.g0_7_m4_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIT7R92_10_LC_6_11_5 .C_ON=1'b0;
    defparam \ALU.b_RNIT7R92_10_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIT7R92_10_LC_6_11_5 .LUT_INIT=16'b0000111111001010;
    LogicCell40 \ALU.b_RNIT7R92_10_LC_6_11_5  (
            .in0(N__26827),
            .in1(N__28525),
            .in2(N__21503),
            .in3(N__34508),
            .lcout(\ALU.N_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNITA7N_0_LC_6_12_0 .C_ON=1'b0;
    defparam \ALU.e_RNITA7N_0_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNITA7N_0_LC_6_12_0 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \ALU.e_RNITA7N_0_LC_6_12_0  (
            .in0(N__28933),
            .in1(N__27124),
            .in2(N__27040),
            .in3(N__28952),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIC4ML1_0_LC_6_12_1 .C_ON=1'b0;
    defparam \ALU.g_RNIC4ML1_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIC4ML1_0_LC_6_12_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.g_RNIC4ML1_0_LC_6_12_1  (
            .in0(N__35707),
            .in1(N__31943),
            .in2(N__21494),
            .in3(N__29138),
            .lcout(\ALU.N_699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIGRS31_0_LC_6_12_2 .C_ON=1'b0;
    defparam \ALU.f_RNIGRS31_0_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIGRS31_0_LC_6_12_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.f_RNIGRS31_0_LC_6_12_2  (
            .in0(N__27126),
            .in1(N__27325),
            .in2(N__36299),
            .in3(N__35051),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1RHK1_0_LC_6_12_3 .C_ON=1'b0;
    defparam \ALU.d_RNI1RHK1_0_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1RHK1_0_LC_6_12_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI1RHK1_0_LC_6_12_3  (
            .in0(N__35708),
            .in1(N__21536),
            .in2(N__21491),
            .in3(N__42194),
            .lcout(\ALU.N_747 ),
            .ltout(\ALU.N_747_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHA1E3_0_LC_6_12_4 .C_ON=1'b0;
    defparam \ALU.d_RNIHA1E3_0_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHA1E3_0_LC_6_12_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.d_RNIHA1E3_0_LC_6_12_4  (
            .in0(N__35206),
            .in1(_gnd_net_),
            .in2(N__21623),
            .in3(N__27256),
            .lcout(\ALU.aluOut_0 ),
            .ltout(\ALU.aluOut_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_N_2L1_LC_6_12_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_N_2L1_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_N_2L1_LC_6_12_5 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \ALU.mult_g0_0_0_N_2L1_LC_6_12_5  (
            .in0(N__39531),
            .in1(_gnd_net_),
            .in2(N__21620),
            .in3(_gnd_net_),
            .lcout(\ALU.g0_0_0_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIBP7N_7_LC_6_12_6 .C_ON=1'b0;
    defparam \ALU.e_RNIBP7N_7_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIBP7N_7_LC_6_12_6 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \ALU.e_RNIBP7N_7_LC_6_12_6  (
            .in0(N__28798),
            .in1(N__27870),
            .in2(N__27041),
            .in3(N__27125),
            .lcout(\ALU.dout_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9BO713_0_LC_6_13_0 .C_ON=1'b0;
    defparam \ALU.d_RNI9BO713_0_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9BO713_0_LC_6_13_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ALU.d_RNI9BO713_0_LC_6_13_0  (
            .in0(N__37933),
            .in1(N__46041),
            .in2(N__21593),
            .in3(N__38190),
            .lcout(\ALU.d_RNI9BO713Z0Z_0 ),
            .ltout(\ALU.d_RNI9BO713Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_0_LC_6_13_1 .C_ON=1'b0;
    defparam \ALU.h_0_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \ALU.h_0_LC_6_13_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.h_0_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__48433),
            .in2(N__21581),
            .in3(N__42326),
            .lcout(\ALU.hZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47687),
            .ce(N__45587),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIHCSL1_0_LC_6_13_2 .C_ON=1'b0;
    defparam \ALU.e_RNIHCSL1_0_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIHCSL1_0_LC_6_13_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.e_RNIHCSL1_0_LC_6_13_2  (
            .in0(N__31041),
            .in1(N__31597),
            .in2(N__28904),
            .in3(N__28850),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPDJU2_0_LC_6_13_3 .C_ON=1'b0;
    defparam \ALU.d_RNIPDJU2_0_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPDJU2_0_LC_6_13_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIPDJU2_0_LC_6_13_3  (
            .in0(N__31262),
            .in1(N__21524),
            .in2(N__21578),
            .in3(N__31607),
            .lcout(),
            .ltout(\ALU.operand2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGTOD3_0_LC_6_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNIGTOD3_0_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGTOD3_0_LC_6_13_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ALU.d_RNIGTOD3_0_LC_6_13_4  (
            .in0(N__21575),
            .in1(N__29292),
            .in2(N__21539),
            .in3(N__25220),
            .lcout(\ALU.N_252_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIE4R7_0_LC_6_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNIE4R7_0_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIE4R7_0_LC_6_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIE4R7_0_LC_6_13_5  (
            .in0(N__21535),
            .in1(N__42193),
            .in2(_gnd_net_),
            .in3(N__32068),
            .lcout(\ALU.d_RNIE4R7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIT0CO_1_LC_6_14_0 .C_ON=1'b0;
    defparam \ALU.g_RNIT0CO_1_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIT0CO_1_LC_6_14_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.g_RNIT0CO_1_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__34884),
            .in2(N__31922),
            .in3(N__29117),
            .lcout(),
            .ltout(\ALU.g_RNIT0COZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNILGSL1_1_LC_6_14_1 .C_ON=1'b0;
    defparam \ALU.e_RNILGSL1_1_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNILGSL1_1_LC_6_14_1 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \ALU.e_RNILGSL1_1_LC_6_14_1  (
            .in0(N__31046),
            .in1(N__31598),
            .in2(N__21659),
            .in3(N__21653),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1MJU2_1_LC_6_14_2 .C_ON=1'b0;
    defparam \ALU.d_RNI1MJU2_1_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1MJU2_1_LC_6_14_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI1MJU2_1_LC_6_14_2  (
            .in0(N__31265),
            .in1(N__28838),
            .in2(N__21656),
            .in3(N__31709),
            .lcout(\ALU.operand2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIPKVJ_1_LC_6_14_3 .C_ON=1'b0;
    defparam \ALU.e_RNIPKVJ_1_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIPKVJ_1_LC_6_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.e_RNIPKVJ_1_LC_6_14_3  (
            .in0(N__34883),
            .in1(N__44596),
            .in2(_gnd_net_),
            .in3(N__26933),
            .lcout(\ALU.e_RNIPKVJZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_11_LC_6_14_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_11_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_11_LC_6_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALU.mult_madd_11_LC_6_14_4  (
            .in0(N__41863),
            .in1(N__37118),
            .in2(N__36945),
            .in3(N__37647),
            .lcout(\ALU.madd_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMH5R6_2_LC_6_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNIMH5R6_2_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMH5R6_2_LC_6_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.d_RNIMH5R6_2_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(N__36861),
            .in2(_gnd_net_),
            .in3(N__38179),
            .lcout(\ALU.a2_b_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_12_0_tz_LC_6_14_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_12_0_tz_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_12_0_tz_LC_6_14_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \ALU.mult_madd_12_0_tz_LC_6_14_6  (
            .in0(N__41862),
            .in1(N__37117),
            .in2(N__36944),
            .in3(N__37646),
            .lcout(\ALU.madd_12_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIVFBD1_15_LC_6_15_0 .C_ON=1'b0;
    defparam \ALU.b_RNIVFBD1_15_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIVFBD1_15_LC_6_15_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.b_RNIVFBD1_15_LC_6_15_0  (
            .in0(N__28496),
            .in1(N__35699),
            .in2(N__25916),
            .in3(N__35576),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC5K02_15_LC_6_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIC5K02_15_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC5K02_15_LC_6_15_1 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.d_RNIC5K02_15_LC_6_15_1  (
            .in0(N__33476),
            .in1(N__35376),
            .in2(N__21626),
            .in3(N__33500),
            .lcout(\ALU.N_762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_1_rep2_e_LC_6_15_2 .C_ON=1'b0;
    defparam \CONTROL.operand1_1_rep2_e_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_1_rep2_e_LC_6_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.operand1_1_rep2_e_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26881),
            .lcout(aluOperand1_1_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47689),
            .ce(N__27727),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5IGD1_5_LC_6_15_3 .C_ON=1'b0;
    defparam \ALU.d_RNI5IGD1_5_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5IGD1_5_LC_6_15_3 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.d_RNI5IGD1_5_LC_6_15_3  (
            .in0(N__31406),
            .in1(N__43400),
            .in2(N__35384),
            .in3(N__23663),
            .lcout(),
            .ltout(\ALU.N_752_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9M073_5_LC_6_15_4 .C_ON=1'b0;
    defparam \ALU.d_RNI9M073_5_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9M073_5_LC_6_15_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNI9M073_5_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__35183),
            .in2(N__21815),
            .in3(N__21809),
            .lcout(\ALU.aluOut_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_fast_e_1_LC_6_15_5 .C_ON=1'b0;
    defparam \CONTROL.operand1_fast_e_1_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_fast_e_1_LC_6_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.operand1_fast_e_1_LC_6_15_5  (
            .in0(N__26882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(aluOperand1_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47689),
            .ce(N__27727),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI7L7N_5_LC_6_15_6 .C_ON=1'b0;
    defparam \ALU.e_RNI7L7N_5_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI7L7N_5_LC_6_15_6 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \ALU.e_RNI7L7N_5_LC_6_15_6  (
            .in0(N__27108),
            .in1(N__44641),
            .in2(N__27039),
            .in3(N__28868),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNI0PML1_5_LC_6_15_7 .C_ON=1'b0;
    defparam \ALU.g_RNI0PML1_5_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNI0PML1_5_LC_6_15_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.g_RNI0PML1_5_LC_6_15_7  (
            .in0(N__35698),
            .in1(N__31835),
            .in2(N__21812),
            .in3(N__29030),
            .lcout(\ALU.N_704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI65RK7_4_LC_6_16_0 .C_ON=1'b0;
    defparam \ALU.d_RNI65RK7_4_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI65RK7_4_LC_6_16_0 .LUT_INIT=16'b0110101001011001;
    LogicCell40 \ALU.d_RNI65RK7_4_LC_6_16_0  (
            .in0(N__42904),
            .in1(N__26605),
            .in2(N__23500),
            .in3(N__23559),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI312TB_4_LC_6_16_1 .C_ON=1'b0;
    defparam \ALU.d_RNI312TB_4_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI312TB_4_LC_6_16_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNI312TB_4_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21803),
            .in3(N__42696),
            .lcout(\ALU.d_RNI312TBZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITKRB7_5_LC_6_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNITKRB7_5_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITKRB7_5_LC_6_16_3 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNITKRB7_5_LC_6_16_3  (
            .in0(N__21788),
            .in1(N__41864),
            .in2(N__24340),
            .in3(N__21724),
            .lcout(\ALU.a3_b_5 ),
            .ltout(\ALU.a3_b_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_94_LC_6_16_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_94_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_94_LC_6_16_4 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \ALU.mult_madd_94_LC_6_16_4  (
            .in0(N__40292),
            .in1(N__22100),
            .in2(N__21674),
            .in3(N__41695),
            .lcout(\ALU.madd_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIE79M7_4_LC_6_16_5 .C_ON=1'b0;
    defparam \ALU.d_RNIE79M7_4_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIE79M7_4_LC_6_16_5 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \ALU.d_RNIE79M7_4_LC_6_16_5  (
            .in0(N__23558),
            .in1(N__23493),
            .in2(N__24341),
            .in3(N__42903),
            .lcout(\ALU.a4_b_4 ),
            .ltout(\ALU.a4_b_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_98_LC_6_16_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_98_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_98_LC_6_16_6 .LUT_INIT=16'b1100000011101000;
    LogicCell40 \ALU.mult_madd_98_LC_6_16_6  (
            .in0(N__40291),
            .in1(N__22094),
            .in2(N__22088),
            .in3(N__41694),
            .lcout(\ALU.madd_98 ),
            .ltout(\ALU.madd_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_139_LC_6_16_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_139_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_139_LC_6_16_7 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \ALU.mult_madd_139_LC_6_16_7  (
            .in0(N__22068),
            .in1(N__38034),
            .in2(N__21980),
            .in3(N__21973),
            .lcout(\ALU.madd_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNO_0_3_LC_7_1_5 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNO_0_3_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNO_0_3_LC_7_1_5 .LUT_INIT=16'b0100010011001101;
    LogicCell40 \FTDI.RXstate_RNO_0_3_LC_7_1_5  (
            .in0(N__24740),
            .in1(N__24659),
            .in2(N__21934),
            .in3(N__24772),
            .lcout(\FTDI.m13_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_1_LC_7_1_6.C_ON=1'b0;
    defparam testState_1_LC_7_1_6.SEQ_MODE=4'b1000;
    defparam testState_1_LC_7_1_6.LUT_INIT=16'b0001001111100000;
    LogicCell40 testState_1_LC_7_1_6 (
            .in0(N__21888),
            .in1(N__30805),
            .in2(N__30302),
            .in3(N__41293),
            .lcout(testStateZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47612),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_0_LC_7_1_7.C_ON=1'b0;
    defparam testState_0_LC_7_1_7.SEQ_MODE=4'b1000;
    defparam testState_0_LC_7_1_7.LUT_INIT=16'b0000001101011100;
    LogicCell40 testState_0_LC_7_1_7 (
            .in0(N__41292),
            .in1(N__21887),
            .in2(N__30809),
            .in3(N__30289),
            .lcout(testStateZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47612),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m40_LC_7_2_0 .C_ON=1'b0;
    defparam \ALU.m40_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \ALU.m40_LC_7_2_0 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \ALU.m40_LC_7_2_0  (
            .in0(N__22581),
            .in1(N__22723),
            .in2(N__21860),
            .in3(N__22436),
            .lcout(),
            .ltout(\ALU.N_41_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_e_0_1_LC_7_2_1 .C_ON=1'b0;
    defparam \CONTROL.aluParams_e_0_1_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluParams_e_0_1_LC_7_2_1 .LUT_INIT=16'b0111011111000000;
    LogicCell40 \CONTROL.aluParams_e_0_1_LC_7_2_1  (
            .in0(N__22437),
            .in1(N__33331),
            .in2(N__21824),
            .in3(N__22742),
            .lcout(aluParams_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47618),
            .ce(N__22139),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPKIOE_7_LC_7_2_2 .C_ON=1'b0;
    defparam \ALU.d_RNIPKIOE_7_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPKIOE_7_LC_7_2_2 .LUT_INIT=16'b1110010101000101;
    LogicCell40 \ALU.d_RNIPKIOE_7_LC_7_2_2  (
            .in0(N__21821),
            .in1(N__40111),
            .in2(N__38972),
            .in3(N__46974),
            .lcout(\ALU.N_473 ),
            .ltout(\ALU.N_473_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4HG101_7_LC_7_2_3 .C_ON=1'b0;
    defparam \ALU.d_RNI4HG101_7_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4HG101_7_LC_7_2_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNI4HG101_7_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(N__38540),
            .in2(N__22745),
            .in3(N__31767),
            .lcout(\ALU.d_RNI4HG101Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m42_ns_1_LC_7_2_4 .C_ON=1'b0;
    defparam \ALU.m42_ns_1_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m42_ns_1_LC_7_2_4 .LUT_INIT=16'b0101010101001100;
    LogicCell40 \ALU.m42_ns_1_LC_7_2_4  (
            .in0(N__22297),
            .in1(N__38888),
            .in2(N__22598),
            .in3(N__33330),
            .lcout(\ALU.m42_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINEO9E_1_LC_7_2_5 .C_ON=1'b0;
    defparam \ALU.d_RNINEO9E_1_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINEO9E_1_LC_7_2_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.d_RNINEO9E_1_LC_7_2_5  (
            .in0(N__38887),
            .in1(N__23144),
            .in2(N__38678),
            .in3(N__23054),
            .lcout(\ALU.lshift_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m286_am_LC_7_2_6 .C_ON=1'b0;
    defparam \ALU.m286_am_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \ALU.m286_am_LC_7_2_6 .LUT_INIT=16'b1000011010000010;
    LogicCell40 \ALU.m286_am_LC_7_2_6  (
            .in0(N__22295),
            .in1(N__22432),
            .in2(N__22597),
            .in3(N__22721),
            .lcout(\ALU.m286_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m286_bm_LC_7_2_7 .C_ON=1'b0;
    defparam \ALU.m286_bm_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m286_bm_LC_7_2_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALU.m286_bm_LC_7_2_7  (
            .in0(N__22722),
            .in1(N__22574),
            .in2(N__22442),
            .in3(N__22296),
            .lcout(\ALU.m286_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICH0SD_3_LC_7_3_0 .C_ON=1'b0;
    defparam \ALU.d_RNICH0SD_3_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICH0SD_3_LC_7_3_0 .LUT_INIT=16'b1101010110000101;
    LogicCell40 \ALU.d_RNICH0SD_3_LC_7_3_0  (
            .in0(N__22829),
            .in1(N__42015),
            .in2(N__38971),
            .in3(N__42996),
            .lcout(),
            .ltout(\ALU.N_469_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI41DBT_3_LC_7_3_1 .C_ON=1'b0;
    defparam \ALU.d_RNI41DBT_3_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI41DBT_3_LC_7_3_1 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.d_RNI41DBT_3_LC_7_3_1  (
            .in0(N__44420),
            .in1(N__38591),
            .in2(N__22166),
            .in3(N__22163),
            .lcout(),
            .ltout(\ALU.rshift_15_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIO3KRQ1_15_LC_7_3_2 .C_ON=1'b0;
    defparam \ALU.c_RNIO3KRQ1_15_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIO3KRQ1_15_LC_7_3_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNIO3KRQ1_15_LC_7_3_2  (
            .in0(N__44421),
            .in1(N__31790),
            .in2(N__22157),
            .in3(N__31771),
            .lcout(\ALU.rshift_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluParams_2_LC_7_3_3 .C_ON=1'b0;
    defparam \CONTROL.aluParams_2_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluParams_2_LC_7_3_3 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \CONTROL.aluParams_2_LC_7_3_3  (
            .in0(N__22154),
            .in1(N__22138),
            .in2(_gnd_net_),
            .in3(N__38592),
            .lcout(aluParams_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47624),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6JKM8_9_LC_7_3_4 .C_ON=1'b0;
    defparam \ALU.d_RNI6JKM8_9_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6JKM8_9_LC_7_3_4 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.d_RNI6JKM8_9_LC_7_3_4  (
            .in0(N__43621),
            .in1(N__39855),
            .in2(N__38969),
            .in3(N__27588),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNICVGTG_11_LC_7_3_5 .C_ON=1'b0;
    defparam \ALU.c_RNICVGTG_11_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNICVGTG_11_LC_7_3_5 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.c_RNICVGTG_11_LC_7_3_5  (
            .in0(N__39012),
            .in1(N__39286),
            .in2(N__22832),
            .in3(N__25370),
            .lcout(\ALU.N_477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI19RM6_1_LC_7_3_6 .C_ON=1'b0;
    defparam \ALU.d_RNI19RM6_1_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI19RM6_1_LC_7_3_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.d_RNI19RM6_1_LC_7_3_6  (
            .in0(N__43622),
            .in1(N__36993),
            .in2(N__38970),
            .in3(N__37427),
            .lcout(\ALU.rshift_3_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINEO9E_0_1_LC_7_4_0 .C_ON=1'b0;
    defparam \ALU.d_RNINEO9E_0_1_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINEO9E_0_1_LC_7_4_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \ALU.d_RNINEO9E_0_1_LC_7_4_0  (
            .in0(N__23053),
            .in1(N__39029),
            .in2(N__38677),
            .in3(N__23143),
            .lcout(\ALU.d_RNINEO9E_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJ1PCQ_1_LC_7_4_1 .C_ON=1'b0;
    defparam \ALU.d_RNIJ1PCQ_1_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJ1PCQ_1_LC_7_4_1 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \ALU.d_RNIJ1PCQ_1_LC_7_4_1  (
            .in0(N__44149),
            .in1(N__23639),
            .in2(N__44521),
            .in3(N__22841),
            .lcout(\ALU.d_RNIJ1PCQZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9HFAU_5_LC_7_4_2 .C_ON=1'b0;
    defparam \ALU.d_RNI9HFAU_5_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9HFAU_5_LC_7_4_2 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.d_RNI9HFAU_5_LC_7_4_2  (
            .in0(N__23052),
            .in1(N__22814),
            .in2(N__38676),
            .in3(N__22787),
            .lcout(),
            .ltout(\ALU.N_311_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKBPO51_5_LC_7_4_3 .C_ON=1'b0;
    defparam \ALU.d_RNIKBPO51_5_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKBPO51_5_LC_7_4_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIKBPO51_5_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(N__44438),
            .in2(N__22781),
            .in3(N__22840),
            .lcout(),
            .ltout(\ALU.lshift_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPFIBI1_9_LC_7_4_4 .C_ON=1'b0;
    defparam \ALU.d_RNIPFIBI1_9_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPFIBI1_9_LC_7_4_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIPFIBI1_9_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__44148),
            .in2(N__22778),
            .in3(N__22775),
            .lcout(\ALU.d_RNIPFIBI1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA28GU1_1_LC_7_4_6 .C_ON=1'b0;
    defparam \ALU.d_RNIA28GU1_1_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA28GU1_1_LC_7_4_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \ALU.d_RNIA28GU1_1_LC_7_4_6  (
            .in0(N__43149),
            .in1(N__22763),
            .in2(_gnd_net_),
            .in3(N__22751),
            .lcout(),
            .ltout(\ALU.d_RNIA28GU1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISQIQP2_1_LC_7_4_7 .C_ON=1'b0;
    defparam \ALU.d_RNISQIQP2_1_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISQIQP2_1_LC_7_4_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNISQIQP2_1_LC_7_4_7  (
            .in0(N__46326),
            .in1(_gnd_net_),
            .in2(N__22955),
            .in3(N__22952),
            .lcout(\ALU.a_15_m5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI2CSHH_13_LC_7_5_0 .C_ON=1'b0;
    defparam \ALU.c_RNI2CSHH_13_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI2CSHH_13_LC_7_5_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.c_RNI2CSHH_13_LC_7_5_0  (
            .in0(N__39150),
            .in1(N__22946),
            .in2(N__38727),
            .in3(N__22933),
            .lcout(),
            .ltout(\ALU.lshift_7_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIONI011_6_LC_7_5_1 .C_ON=1'b0;
    defparam \ALU.d_RNIONI011_6_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIONI011_6_LC_7_5_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.d_RNIONI011_6_LC_7_5_1  (
            .in0(N__38689),
            .in1(N__22919),
            .in2(N__22898),
            .in3(N__22893),
            .lcout(),
            .ltout(\ALU.N_315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINQ8VM1_6_LC_7_5_2 .C_ON=1'b0;
    defparam \ALU.d_RNINQ8VM1_6_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINQ8VM1_6_LC_7_5_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNINQ8VM1_6_LC_7_5_2  (
            .in0(N__44487),
            .in1(_gnd_net_),
            .in2(N__22871),
            .in3(N__27958),
            .lcout(),
            .ltout(\ALU.lshift_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3O3A42_13_LC_7_5_3 .C_ON=1'b0;
    defparam \ALU.c_RNI3O3A42_13_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3O3A42_13_LC_7_5_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.c_RNI3O3A42_13_LC_7_5_3  (
            .in0(N__44150),
            .in1(_gnd_net_),
            .in2(N__22868),
            .in3(N__22865),
            .lcout(),
            .ltout(\ALU.a_15_m4_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI88B4N2_13_LC_7_5_4 .C_ON=1'b0;
    defparam \ALU.c_RNI88B4N2_13_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI88B4N2_13_LC_7_5_4 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \ALU.c_RNI88B4N2_13_LC_7_5_4  (
            .in0(N__46330),
            .in1(_gnd_net_),
            .in2(N__22856),
            .in3(N__24791),
            .lcout(c_RNI88B4N2_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIV49JL_1_LC_7_5_5 .C_ON=1'b0;
    defparam \ALU.d_RNIV49JL_1_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIV49JL_1_LC_7_5_5 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ALU.d_RNIV49JL_1_LC_7_5_5  (
            .in0(N__39037),
            .in1(N__23142),
            .in2(N__38729),
            .in3(N__22853),
            .lcout(\ALU.N_420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI1HDEU1_13_LC_7_5_6 .C_ON=1'b0;
    defparam \ALU.c_RNI1HDEU1_13_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI1HDEU1_13_LC_7_5_6 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \ALU.c_RNI1HDEU1_13_LC_7_5_6  (
            .in0(N__23104),
            .in1(N__23089),
            .in2(N__44522),
            .in3(N__22847),
            .lcout(\ALU.lshift_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBSS27_1_LC_7_5_7 .C_ON=1'b0;
    defparam \ALU.d_RNIBSS27_1_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBSS27_1_LC_7_5_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ALU.d_RNIBSS27_1_LC_7_5_7  (
            .in0(N__38685),
            .in1(N__39149),
            .in2(_gnd_net_),
            .in3(N__23141),
            .lcout(\ALU.N_416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICIR67_3_LC_7_6_0 .C_ON=1'b0;
    defparam \ALU.d_RNICIR67_3_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICIR67_3_LC_7_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNICIR67_3_LC_7_6_0  (
            .in0(N__43714),
            .in1(N__36953),
            .in2(_gnd_net_),
            .in3(N__41977),
            .lcout(\ALU.N_377 ),
            .ltout(\ALU.N_377_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIOHBUD_1_LC_7_6_1 .C_ON=1'b0;
    defparam \ALU.d_RNIOHBUD_1_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIOHBUD_1_LC_7_6_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIOHBUD_1_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__39147),
            .in2(N__23027),
            .in3(N__23137),
            .lcout(\ALU.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIN9H77_3_LC_7_6_2 .C_ON=1'b0;
    defparam \ALU.d_RNIN9H77_3_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIN9H77_3_LC_7_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIN9H77_3_LC_7_6_2  (
            .in0(N__43715),
            .in1(N__41978),
            .in2(_gnd_net_),
            .in3(N__42980),
            .lcout(\ALU.N_216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIADS9I_0_LC_7_6_3 .C_ON=1'b0;
    defparam \ALU.d_RNIADS9I_0_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIADS9I_0_LC_7_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIADS9I_0_LC_7_6_3  (
            .in0(N__38724),
            .in1(N__23018),
            .in2(_gnd_net_),
            .in3(N__23012),
            .lcout(\ALU.N_419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGFQD6_1_LC_7_6_4 .C_ON=1'b0;
    defparam \ALU.d_RNIGFQD6_1_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGFQD6_1_LC_7_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNIGFQD6_1_LC_7_6_4  (
            .in0(N__43713),
            .in1(N__36952),
            .in2(_gnd_net_),
            .in3(N__37419),
            .lcout(\ALU.N_376 ),
            .ltout(\ALU.N_376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEBMRA_0_LC_7_6_5 .C_ON=1'b0;
    defparam \ALU.d_RNIEBMRA_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEBMRA_0_LC_7_6_5 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ALU.d_RNIEBMRA_0_LC_7_6_5  (
            .in0(N__38725),
            .in1(N__39148),
            .in2(N__22997),
            .in3(N__27245),
            .lcout(),
            .ltout(\ALU.d_RNIEBMRAZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFPKBA1_0_LC_7_6_6 .C_ON=1'b0;
    defparam \ALU.d_RNIFPKBA1_0_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFPKBA1_0_LC_7_6_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIFPKBA1_0_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__44444),
            .in2(N__22994),
            .in3(N__22991),
            .lcout(\ALU.lshift_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICGVRD_3_LC_7_6_7 .C_ON=1'b0;
    defparam \ALU.d_RNICGVRD_3_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICGVRD_3_LC_7_6_7 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \ALU.d_RNICGVRD_3_LC_7_6_7  (
            .in0(N__41979),
            .in1(N__39146),
            .in2(N__36997),
            .in3(N__23111),
            .lcout(\ALU.N_468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIG5BH6_3_LC_7_7_0 .C_ON=1'b0;
    defparam \ALU.d_RNIG5BH6_3_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIG5BH6_3_LC_7_7_0 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIG5BH6_3_LC_7_7_0  (
            .in0(N__23917),
            .in1(N__37371),
            .in2(N__26598),
            .in3(N__24014),
            .lcout(\ALU.a1_b_3 ),
            .ltout(\ALU.a1_b_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_13_LC_7_7_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_13_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_13_LC_7_7_1 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ALU.mult_madd_13_LC_7_7_1  (
            .in0(N__23219),
            .in1(N__23158),
            .in2(N__23192),
            .in3(N__23189),
            .lcout(\ALU.madd_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKFBA7_3_LC_7_7_2 .C_ON=1'b0;
    defparam \ALU.d_RNIKFBA7_3_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKFBA7_3_LC_7_7_2 .LUT_INIT=16'b0101110000000000;
    LogicCell40 \ALU.d_RNIKFBA7_3_LC_7_7_2  (
            .in0(N__23918),
            .in1(N__24013),
            .in2(N__26599),
            .in3(N__37994),
            .lcout(\ALU.a0_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIR5FE6_1_LC_7_7_3 .C_ON=1'b0;
    defparam \ALU.d_RNIR5FE6_1_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIR5FE6_1_LC_7_7_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \ALU.d_RNIR5FE6_1_LC_7_7_3  (
            .in0(N__37995),
            .in1(_gnd_net_),
            .in2(N__37425),
            .in3(N__43684),
            .lcout(\ALU.N_375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILPO64_4_LC_7_7_4 .C_ON=1'b0;
    defparam \ALU.d_RNILPO64_4_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILPO64_4_LC_7_7_4 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \ALU.d_RNILPO64_4_LC_7_7_4  (
            .in0(N__23456),
            .in1(_gnd_net_),
            .in2(N__26600),
            .in3(N__23568),
            .lcout(\ALU.N_231_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI35AS3_3_LC_7_7_5 .C_ON=1'b0;
    defparam \ALU.d_RNI35AS3_3_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI35AS3_3_LC_7_7_5 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ALU.d_RNI35AS3_3_LC_7_7_5  (
            .in0(N__24015),
            .in1(N__26549),
            .in2(_gnd_net_),
            .in3(N__23919),
            .lcout(\ALU.N_237_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNICVFN6_1_LC_7_7_6 .C_ON=1'b0;
    defparam \ALU.d_RNICVFN6_1_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNICVFN6_1_LC_7_7_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.d_RNICVFN6_1_LC_7_7_6  (
            .in0(N__43683),
            .in1(N__37372),
            .in2(N__39140),
            .in3(N__37996),
            .lcout(\ALU.rshift_3_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9GDQS_1_LC_7_7_7 .C_ON=1'b0;
    defparam \ALU.d_RNI9GDQS_1_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9GDQS_1_LC_7_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNI9GDQS_1_LC_7_7_7  (
            .in0(N__38726),
            .in1(N__23105),
            .in2(_gnd_net_),
            .in3(N__23090),
            .lcout(\ALU.N_422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI1FPGN1_10_LC_7_8_0 .C_ON=1'b0;
    defparam \ALU.a_RNI1FPGN1_10_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI1FPGN1_10_LC_7_8_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ALU.a_RNI1FPGN1_10_LC_7_8_0  (
            .in0(N__23078),
            .in1(_gnd_net_),
            .in2(N__44218),
            .in3(N__23258),
            .lcout(),
            .ltout(\ALU.a_15_m4_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI5V90O2_10_LC_7_8_1 .C_ON=1'b0;
    defparam \ALU.c_RNI5V90O2_10_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI5V90O2_10_LC_7_8_1 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \ALU.c_RNI5V90O2_10_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__23069),
            .in2(N__23057),
            .in3(N__46382),
            .lcout(c_RNI5V90O2_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIJQBMC_10_LC_7_8_2 .C_ON=1'b0;
    defparam \ALU.a_RNIJQBMC_10_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIJQBMC_10_LC_7_8_2 .LUT_INIT=16'b0011100111010100;
    LogicCell40 \ALU.a_RNIJQBMC_10_LC_7_8_2  (
            .in0(N__23252),
            .in1(N__27550),
            .in2(N__39606),
            .in3(N__47279),
            .lcout(\ALU.a_15_m2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_10_LC_7_8_3 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_10_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_10_LC_7_8_3 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.a_15_m2_ns_1_10_LC_7_8_3  (
            .in0(N__47278),
            .in1(N__44188),
            .in2(N__43938),
            .in3(N__43729),
            .lcout(\ALU.a_15_m2_ns_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_9_c_RNI8H83V_LC_7_8_4 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_9_c_RNI8H83V_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_9_c_RNI8H83V_LC_7_8_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ALU.un9_addsub_cry_9_c_RNI8H83V_LC_7_8_4  (
            .in0(N__42522),
            .in1(N__39488),
            .in2(_gnd_net_),
            .in3(N__23246),
            .lcout(),
            .ltout(un9_addsub_cry_9_c_RNI8H83V_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_RNINNN4N3_0_LC_7_8_5 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_RNINNN4N3_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_RNINNN4N3_0_LC_7_8_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \CONTROL.aluOperation_RNINNN4N3_0_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__48329),
            .in2(N__23237),
            .in3(N__23234),
            .lcout(aluOperation_RNINNN4N3_0),
            .ltout(aluOperation_RNINNN4N3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_10_LC_7_8_6 .C_ON=1'b0;
    defparam \ALU.a_10_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \ALU.a_10_LC_7_8_6 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.a_10_LC_7_8_6  (
            .in0(N__48330),
            .in1(N__45967),
            .in2(N__23228),
            .in3(N__34411),
            .lcout(\ALU.aZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47656),
            .ce(N__44837),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIM5AD1_11_LC_7_9_0 .C_ON=1'b0;
    defparam \ALU.b_RNIM5AD1_11_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIM5AD1_11_LC_7_9_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.b_RNIM5AD1_11_LC_7_9_0  (
            .in0(N__35906),
            .in1(N__28475),
            .in2(N__35582),
            .in3(N__28457),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRII02_11_LC_7_9_1 .C_ON=1'b0;
    defparam \ALU.d_RNIRII02_11_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRII02_11_LC_7_9_1 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNIRII02_11_LC_7_9_1  (
            .in0(N__31136),
            .in1(N__35374),
            .in2(N__23225),
            .in3(N__31157),
            .lcout(\ALU.N_758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI41LF1_11_LC_7_9_2 .C_ON=1'b0;
    defparam \ALU.a_RNI41LF1_11_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI41LF1_11_LC_7_9_2 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \ALU.a_RNI41LF1_11_LC_7_9_2  (
            .in0(N__30830),
            .in1(N__35996),
            .in2(N__35911),
            .in3(N__32489),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI76HQ1_11_LC_7_9_3 .C_ON=1'b0;
    defparam \ALU.c_RNI76HQ1_11_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI76HQ1_11_LC_7_9_3 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.c_RNI76HQ1_11_LC_7_9_3  (
            .in0(N__34112),
            .in1(N__35375),
            .in2(N__23222),
            .in3(N__31307),
            .lcout(),
            .ltout(\ALU.N_710_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI64TU3_11_LC_7_9_4 .C_ON=1'b0;
    defparam \ALU.c_RNI64TU3_11_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI64TU3_11_LC_7_9_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.c_RNI64TU3_11_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__23378),
            .in2(N__23372),
            .in3(N__35222),
            .lcout(\ALU.aluOut_11 ),
            .ltout(\ALU.aluOut_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_484_6_LC_7_9_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_484_6_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_484_6_LC_7_9_5 .LUT_INIT=16'b0010001011010010;
    LogicCell40 \ALU.mult_madd_484_6_LC_7_9_5  (
            .in0(N__27499),
            .in1(N__28089),
            .in2(N__23369),
            .in3(N__42644),
            .lcout(\ALU.madd_484_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJM067_1_LC_7_10_0 .C_ON=1'b0;
    defparam \ALU.d_RNIJM067_1_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJM067_1_LC_7_10_0 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \ALU.d_RNIJM067_1_LC_7_10_0  (
            .in0(N__37348),
            .in1(N__43933),
            .in2(_gnd_net_),
            .in3(N__37716),
            .lcout(\ALU.d_RNIJM067Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI80E86_1_LC_7_10_1 .C_ON=1'b0;
    defparam \ALU.d_RNI80E86_1_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI80E86_1_LC_7_10_1 .LUT_INIT=16'b0110110001100011;
    LogicCell40 \ALU.d_RNI80E86_1_LC_7_10_1  (
            .in0(N__23338),
            .in1(N__37347),
            .in2(N__26642),
            .in3(N__23300),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC4AT9_1_LC_7_10_2 .C_ON=1'b0;
    defparam \ALU.d_RNIC4AT9_1_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC4AT9_1_LC_7_10_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNIC4AT9_1_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23354),
            .in3(N__23278),
            .lcout(\ALU.d_RNIC4AT9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI5NDI1_1_LC_7_10_3 .C_ON=1'b0;
    defparam \ALU.e_RNI5NDI1_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI5NDI1_1_LC_7_10_3 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \ALU.e_RNI5NDI1_1_LC_7_10_3  (
            .in0(N__27377),
            .in1(N__35224),
            .in2(N__35385),
            .in3(N__26945),
            .lcout(),
            .ltout(\ALU.dout_7_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID01L2_1_LC_7_10_4 .C_ON=1'b0;
    defparam \ALU.d_RNID01L2_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID01L2_1_LC_7_10_4 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNID01L2_1_LC_7_10_4  (
            .in0(N__28826),
            .in1(N__35225),
            .in2(N__23345),
            .in3(N__31724),
            .lcout(\ALU.aluOut_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI44SK3_1_LC_7_10_5 .C_ON=1'b0;
    defparam \ALU.d_RNI44SK3_1_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI44SK3_1_LC_7_10_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \ALU.d_RNI44SK3_1_LC_7_10_5  (
            .in0(N__30049),
            .in1(N__23337),
            .in2(_gnd_net_),
            .in3(N__23299),
            .lcout(\ALU.N_249_0 ),
            .ltout(\ALU.N_249_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI61SHA_1_LC_7_10_6 .C_ON=1'b0;
    defparam \ALU.d_RNI61SHA_1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI61SHA_1_LC_7_10_6 .LUT_INIT=16'b1010111010001100;
    LogicCell40 \ALU.d_RNI61SHA_1_LC_7_10_6  (
            .in0(N__37349),
            .in1(N__24594),
            .in2(N__23261),
            .in3(N__37717),
            .lcout(),
            .ltout(\ALU.d_RNI61SHAZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9CMFI_1_LC_7_10_7 .C_ON=1'b0;
    defparam \ALU.d_RNI9CMFI_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9CMFI_1_LC_7_10_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNI9CMFI_1_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__47277),
            .in2(N__23648),
            .in3(N__23645),
            .lcout(\ALU.a_15_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIK6LL_4_LC_7_11_0 .C_ON=1'b0;
    defparam \ALU.g_RNIK6LL_4_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIK6LL_4_LC_7_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_RNIK6LL_4_LC_7_11_0  (
            .in0(N__32081),
            .in1(N__31861),
            .in2(_gnd_net_),
            .in3(N__29047),
            .lcout(),
            .ltout(\ALU.g_RNIK6LLZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI5F2S1_4_LC_7_11_1 .C_ON=1'b0;
    defparam \ALU.e_RNI5F2S1_4_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI5F2S1_4_LC_7_11_1 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \ALU.e_RNI5F2S1_4_LC_7_11_1  (
            .in0(N__31261),
            .in1(N__35027),
            .in2(N__23627),
            .in3(N__23624),
            .lcout(\ALU.operand2_7_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIGQ8H_4_LC_7_11_2 .C_ON=1'b0;
    defparam \ALU.e_RNIGQ8H_4_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIGQ8H_4_LC_7_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.e_RNIGQ8H_4_LC_7_11_2  (
            .in0(N__32080),
            .in1(N__27941),
            .in2(_gnd_net_),
            .in3(N__26963),
            .lcout(\ALU.e_RNIGQ8HZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAS7T6_4_LC_7_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIAS7T6_4_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAS7T6_4_LC_7_11_3 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIAS7T6_4_LC_7_11_3  (
            .in0(N__23487),
            .in1(N__37318),
            .in2(N__24290),
            .in3(N__23523),
            .lcout(\ALU.a1_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3GJL7_4_LC_7_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNI3GJL7_4_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3GJL7_4_LC_7_11_4 .LUT_INIT=16'b0010111000000000;
    LogicCell40 \ALU.d_RNI3GJL7_4_LC_7_11_4  (
            .in0(N__23524),
            .in1(N__24253),
            .in2(N__23489),
            .in3(N__36813),
            .lcout(\ALU.a2_b_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1LUH3_4_LC_7_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNI1LUH3_4_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1LUH3_4_LC_7_11_5 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.d_RNI1LUH3_4_LC_7_11_5  (
            .in0(N__24389),
            .in1(N__45389),
            .in2(N__33104),
            .in3(N__23579),
            .lcout(\ALU.operand2_4 ),
            .ltout(\ALU.operand2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITR684_4_LC_7_11_6 .C_ON=1'b0;
    defparam \ALU.d_RNITR684_4_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITR684_4_LC_7_11_6 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \ALU.d_RNITR684_4_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__23488),
            .in2(N__23396),
            .in3(N__24249),
            .lcout(\ALU.N_231_0 ),
            .ltout(\ALU.N_231_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_168_LC_7_11_7 .C_ON=1'b0;
    defparam \ALU.mult_madd_168_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_168_LC_7_11_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ALU.mult_madd_168_LC_7_11_7  (
            .in0(N__39751),
            .in1(N__46648),
            .in2(N__23393),
            .in3(N__37715),
            .lcout(\ALU.madd_93_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIGOP81_10_LC_7_12_0 .C_ON=1'b0;
    defparam \ALU.a_RNIGOP81_10_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIGOP81_10_LC_7_12_0 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \ALU.a_RNIGOP81_10_LC_7_12_0  (
            .in0(N__28593),
            .in1(N__23706),
            .in2(N__27337),
            .in3(N__27129),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI1PNQ1_10_LC_7_12_1 .C_ON=1'b0;
    defparam \ALU.c_RNI1PNQ1_10_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI1PNQ1_10_LC_7_12_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNI1PNQ1_10_LC_7_12_1  (
            .in0(N__35709),
            .in1(N__34283),
            .in2(N__23678),
            .in3(N__34933),
            .lcout(\ALU.N_709 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNI471O1_10_LC_7_12_2 .C_ON=1'b0;
    defparam \ALU.b_RNI471O1_10_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNI471O1_10_LC_7_12_2 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \ALU.b_RNI471O1_10_LC_7_12_2  (
            .in0(N__26828),
            .in1(N__28526),
            .in2(N__35985),
            .in3(N__35876),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7I9B2_10_LC_7_12_3 .C_ON=1'b0;
    defparam \ALU.d_RNI7I9B2_10_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7I9B2_10_LC_7_12_3 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.d_RNI7I9B2_10_LC_7_12_3  (
            .in0(N__28426),
            .in1(N__35352),
            .in2(N__23675),
            .in3(N__24423),
            .lcout(),
            .ltout(\ALU.N_757_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNICMQ94_10_LC_7_12_4 .C_ON=1'b0;
    defparam \ALU.c_RNICMQ94_10_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNICMQ94_10_LC_7_12_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.c_RNICMQ94_10_LC_7_12_4  (
            .in0(N__35207),
            .in1(_gnd_net_),
            .in2(N__23672),
            .in3(N__23669),
            .lcout(\ALU.aluOut_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_2_rep1_e_LC_7_12_5 .C_ON=1'b0;
    defparam \CONTROL.operand1_2_rep1_e_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_2_rep1_e_LC_7_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.operand1_2_rep1_e_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27185),
            .lcout(aluOperand1_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47680),
            .ce(N__27697),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIQ5T31_5_LC_7_12_6 .C_ON=1'b0;
    defparam \ALU.f_RNIQ5T31_5_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIQ5T31_5_LC_7_12_6 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.f_RNIQ5T31_5_LC_7_12_6  (
            .in0(N__27321),
            .in1(N__48965),
            .in2(N__36440),
            .in3(N__27128),
            .lcout(\ALU.dout_6_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGUO51_6_LC_7_13_0 .C_ON=1'b0;
    defparam \ALU.d_RNIGUO51_6_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGUO51_6_LC_7_13_0 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \ALU.d_RNIGUO51_6_LC_7_13_0  (
            .in0(N__35013),
            .in1(N__43373),
            .in2(N__45622),
            .in3(N__23720),
            .lcout(),
            .ltout(\ALU.N_865_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDHB63_6_LC_7_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIDHB63_6_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDHB63_6_LC_7_13_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIDHB63_6_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__32995),
            .in2(N__23651),
            .in3(N__23789),
            .lcout(\ALU.operand2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIKC1M_6_LC_7_13_2 .C_ON=1'b0;
    defparam \ALU.e_RNIKC1M_6_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIKC1M_6_LC_7_13_2 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \ALU.e_RNIKC1M_6_LC_7_13_2  (
            .in0(N__27897),
            .in1(N__28622),
            .in2(N__31044),
            .in3(N__32049),
            .lcout(),
            .ltout(\ALU.operand2_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIBICH1_6_LC_7_13_3 .C_ON=1'b0;
    defparam \ALU.g_RNIBICH1_6_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIBICH1_6_LC_7_13_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.g_RNIBICH1_6_LC_7_13_3  (
            .in0(N__28975),
            .in1(N__29015),
            .in2(N__23792),
            .in3(N__35012),
            .lcout(\ALU.N_817 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDTEA7_6_LC_7_13_4 .C_ON=1'b0;
    defparam \ALU.d_RNIDTEA7_6_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDTEA7_6_LC_7_13_4 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \ALU.d_RNIDTEA7_6_LC_7_13_4  (
            .in0(N__26690),
            .in1(N__26279),
            .in2(N__24315),
            .in3(N__46622),
            .lcout(\ALU.a6_b_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKTLA7_6_LC_7_13_5 .C_ON=1'b0;
    defparam \ALU.d_RNIKTLA7_6_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKTLA7_6_LC_7_13_5 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIKTLA7_6_LC_7_13_5  (
            .in0(N__26278),
            .in1(N__41809),
            .in2(N__24313),
            .in3(N__26689),
            .lcout(\ALU.a3_b_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNINI7O_6_LC_7_13_6 .C_ON=1'b0;
    defparam \ALU.f_RNINI7O_6_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNINI7O_6_LC_7_13_6 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \ALU.f_RNINI7O_6_LC_7_13_6  (
            .in0(N__36419),
            .in1(N__45129),
            .in2(N__31045),
            .in3(N__48815),
            .lcout(\ALU.operand2_6_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNII4LL_3_LC_7_14_0 .C_ON=1'b0;
    defparam \ALU.g_RNII4LL_3_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNII4LL_3_LC_7_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.g_RNII4LL_3_LC_7_14_0  (
            .in0(N__29072),
            .in1(N__31879),
            .in2(_gnd_net_),
            .in3(N__32069),
            .lcout(\ALU.g_RNII4LLZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID7IK1_3_LC_7_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNID7IK1_3_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID7IK1_3_LC_7_14_1 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \ALU.d_RNID7IK1_3_LC_7_14_1  (
            .in0(N__35671),
            .in1(N__45158),
            .in2(N__45185),
            .in3(N__27365),
            .lcout(),
            .ltout(\ALU.N_750_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI932E3_3_LC_7_14_2 .C_ON=1'b0;
    defparam \ALU.d_RNI932E3_3_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI932E3_3_LC_7_14_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.d_RNI932E3_3_LC_7_14_2  (
            .in0(N__23825),
            .in1(_gnd_net_),
            .in2(N__23714),
            .in3(N__35221),
            .lcout(\ALU.aluOut_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7PG73_3_LC_7_14_3 .C_ON=1'b0;
    defparam \ALU.d_RNI7PG73_3_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7PG73_3_LC_7_14_3 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \ALU.d_RNI7PG73_3_LC_7_14_3  (
            .in0(N__44987),
            .in1(N__43247),
            .in2(N__33103),
            .in3(N__23810),
            .lcout(\ALU.operand2_3 ),
            .ltout(\ALU.operand2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI1CMM3_3_LC_7_14_4 .C_ON=1'b0;
    defparam \ALU.d_RNI1CMM3_3_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI1CMM3_3_LC_7_14_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \ALU.d_RNI1CMM3_3_LC_7_14_4  (
            .in0(N__23938),
            .in1(_gnd_net_),
            .in2(N__23711),
            .in3(N__25221),
            .lcout(\ALU.N_237_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKAQB7_3_LC_7_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNIKAQB7_3_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKAQB7_3_LC_7_14_5 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \ALU.d_RNIKAQB7_3_LC_7_14_5  (
            .in0(N__23974),
            .in1(N__23940),
            .in2(N__24316),
            .in3(N__41861),
            .lcout(\ALU.a3_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHR4B7_3_LC_7_14_6 .C_ON=1'b0;
    defparam \ALU.d_RNIHR4B7_3_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHR4B7_3_LC_7_14_6 .LUT_INIT=16'b0100110001000000;
    LogicCell40 \ALU.d_RNIHR4B7_3_LC_7_14_6  (
            .in0(N__23937),
            .in1(N__36844),
            .in2(N__24314),
            .in3(N__23972),
            .lcout(\ALU.a2_b_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC8CA7_3_LC_7_14_7 .C_ON=1'b0;
    defparam \ALU.d_RNIC8CA7_3_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC8CA7_3_LC_7_14_7 .LUT_INIT=16'b0011101011000101;
    LogicCell40 \ALU.d_RNIC8CA7_3_LC_7_14_7  (
            .in0(N__23973),
            .in1(N__23939),
            .in2(N__26641),
            .in3(N__41860),
            .lcout(\ALU.un2_addsub_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIDK21B_3_LC_7_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIDK21B_3_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIDK21B_3_LC_7_15_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ALU.d_RNIDK21B_3_LC_7_15_1  (
            .in0(N__23852),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41667),
            .lcout(\ALU.d_RNIDK21BZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI3H7N_3_LC_7_15_2 .C_ON=1'b0;
    defparam \ALU.e_RNI3H7N_3_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI3H7N_3_LC_7_15_2 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \ALU.e_RNI3H7N_3_LC_7_15_2  (
            .in0(N__44908),
            .in1(N__27029),
            .in2(N__27120),
            .in3(N__28637),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIOGML1_3_LC_7_15_3 .C_ON=1'b0;
    defparam \ALU.g_RNIOGML1_3_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIOGML1_3_LC_7_15_3 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.g_RNIOGML1_3_LC_7_15_3  (
            .in0(N__31883),
            .in1(N__35706),
            .in2(N__23828),
            .in3(N__29071),
            .lcout(\ALU.N_702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNITOVJ_3_LC_7_15_4 .C_ON=1'b0;
    defparam \ALU.e_RNITOVJ_3_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNITOVJ_3_LC_7_15_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.e_RNITOVJ_3_LC_7_15_4  (
            .in0(N__44907),
            .in1(N__28636),
            .in2(_gnd_net_),
            .in3(N__34891),
            .lcout(),
            .ltout(\ALU.e_RNITOVJZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIGBPU1_3_LC_7_15_5 .C_ON=1'b0;
    defparam \ALU.e_RNIGBPU1_3_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIGBPU1_3_LC_7_15_5 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \ALU.e_RNIGBPU1_3_LC_7_15_5  (
            .in0(N__31264),
            .in1(N__23819),
            .in2(N__23813),
            .in3(N__35028),
            .lcout(\ALU.operand2_7_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_6_c_RNIUKMKR_LC_7_15_6 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_6_c_RNIUKMKR_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_6_c_RNIUKMKR_LC_7_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.un9_addsub_cry_6_c_RNIUKMKR_LC_7_15_6  (
            .in0(N__42530),
            .in1(N__40145),
            .in2(_gnd_net_),
            .in3(N__23804),
            .lcout(\ALU.un9_addsub_cry_6_c_RNIUKMKRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_63_LC_7_16_0 .C_ON=1'b0;
    defparam \ALU.mult_madd_63_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_63_LC_7_16_0 .LUT_INIT=16'b1110100010001000;
    LogicCell40 \ALU.mult_madd_63_LC_7_16_0  (
            .in0(N__24545),
            .in1(N__24533),
            .in2(N__46682),
            .in3(N__37718),
            .lcout(\ALU.madd_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_2_l_fx_LC_7_16_1 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_2_l_fx_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_2_l_fx_LC_7_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ALU.mult_madd_axb_2_l_fx_LC_7_16_1  (
            .in0(N__24500),
            .in1(N__24488),
            .in2(N__25838),
            .in3(N__24470),
            .lcout(\ALU.madd_axb_2_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_9_LC_7_16_2 .C_ON=1'b0;
    defparam \ALU.h_9_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \ALU.h_9_LC_7_16_2 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.h_9_LC_7_16_2  (
            .in0(N__48597),
            .in1(N__36275),
            .in2(N__46162),
            .in3(N__36205),
            .lcout(\ALU.hZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47690),
            .ce(N__45574),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI2B0L_9_LC_7_16_3 .C_ON=1'b0;
    defparam \ALU.d_RNI2B0L_9_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI2B0L_9_LC_7_16_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNI2B0L_9_LC_7_16_3  (
            .in0(N__32817),
            .in1(N__32798),
            .in2(_gnd_net_),
            .in3(N__45338),
            .lcout(\ALU.d_RNI2B0LZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIORSD1_15_LC_7_16_4 .C_ON=1'b0;
    defparam \ALU.b_RNIORSD1_15_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIORSD1_15_LC_7_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.b_RNIORSD1_15_LC_7_16_4  (
            .in0(N__25912),
            .in1(N__28495),
            .in2(_gnd_net_),
            .in3(N__45337),
            .lcout(\ALU.b_RNIORSD1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNII1LU_10_LC_7_16_5 .C_ON=1'b0;
    defparam \ALU.d_RNII1LU_10_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNII1LU_10_LC_7_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNII1LU_10_LC_7_16_5  (
            .in0(N__45336),
            .in1(N__24431),
            .in2(_gnd_net_),
            .in3(N__28427),
            .lcout(\ALU.d_RNII1LUZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO00L_4_LC_7_16_6 .C_ON=1'b0;
    defparam \ALU.d_RNIO00L_4_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO00L_4_LC_7_16_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNIO00L_4_LC_7_16_6  (
            .in0(N__36535),
            .in1(N__45335),
            .in2(_gnd_net_),
            .in3(N__28990),
            .lcout(\ALU.d_RNIO00LZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_8_LC_9_1_0 .C_ON=1'b0;
    defparam \ALU.d_8_LC_9_1_0 .SEQ_MODE=4'b1000;
    defparam \ALU.d_8_LC_9_1_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_8_LC_9_1_0  (
            .in0(N__48105),
            .in1(N__47888),
            .in2(_gnd_net_),
            .in3(N__47778),
            .lcout(\ALU.dZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47606),
            .ce(N__43324),
            .sr(_gnd_net_));
    defparam \FTDI.gap_0_LC_9_2_0 .C_ON=1'b0;
    defparam \FTDI.gap_0_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \FTDI.gap_0_LC_9_2_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \FTDI.gap_0_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(N__29206),
            .in2(_gnd_net_),
            .in3(N__29195),
            .lcout(\FTDI.gapZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_2_LC_9_2_1 .C_ON=1'b0;
    defparam \FTDI.baudAcc_2_LC_9_2_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_2_LC_9_2_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \FTDI.baudAcc_2_LC_9_2_1  (
            .in0(N__29570),
            .in1(N__29587),
            .in2(_gnd_net_),
            .in3(N__30422),
            .lcout(\FTDI.baudAccZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_RNO_0_0_LC_9_2_2 .C_ON=1'b0;
    defparam \FTDI.RXstate_RNO_0_0_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \FTDI.RXstate_RNO_0_0_LC_9_2_2 .LUT_INIT=16'b0111010111110100;
    LogicCell40 \FTDI.RXstate_RNO_0_0_LC_9_2_2  (
            .in0(N__24627),
            .in1(N__24776),
            .in2(N__29266),
            .in3(N__24722),
            .lcout(),
            .ltout(\FTDI.N_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_0_LC_9_2_3 .C_ON=1'b0;
    defparam \FTDI.RXstate_0_LC_9_2_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_0_LC_9_2_3 .LUT_INIT=16'b0000111110001000;
    LogicCell40 \FTDI.RXstate_0_LC_9_2_3  (
            .in0(N__29262),
            .in1(N__24632),
            .in2(N__24746),
            .in3(N__24681),
            .lcout(\FTDI.RXstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_1_LC_9_2_4 .C_ON=1'b0;
    defparam \FTDI.RXstate_1_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_1_LC_9_2_4 .LUT_INIT=16'b0111000010000000;
    LogicCell40 \FTDI.RXstate_1_LC_9_2_4  (
            .in0(N__24682),
            .in1(N__29261),
            .in2(N__24645),
            .in3(N__24723),
            .lcout(\FTDI.RXstateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.RXstate_3_LC_9_2_7 .C_ON=1'b0;
    defparam \FTDI.RXstate_3_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.RXstate_3_LC_9_2_7 .LUT_INIT=16'b1000110011101110;
    LogicCell40 \FTDI.RXstate_3_LC_9_2_7  (
            .in0(N__24701),
            .in1(N__24631),
            .in2(N__29267),
            .in3(N__24680),
            .lcout(\FTDI.RXstateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2s2_LC_9_3_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2s2_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2s2_LC_9_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.a_15_m2s2_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__38973),
            .in2(_gnd_net_),
            .in3(N__44121),
            .lcout(\ALU.a_15_sm0 ),
            .ltout(\ALU.a_15_sm0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_12_LC_9_3_1 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_12_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_12_LC_9_3_1 .LUT_INIT=16'b0000010111110101;
    LogicCell40 \ALU.a_15_m2_ns_1_12_LC_9_3_1  (
            .in0(N__24596),
            .in1(_gnd_net_),
            .in2(N__24602),
            .in3(N__43900),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNISG1SC_12_LC_9_3_2 .C_ON=1'b0;
    defparam \ALU.c_RNISG1SC_12_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNISG1SC_12_LC_9_3_2 .LUT_INIT=16'b0110011110000110;
    LogicCell40 \ALU.c_RNISG1SC_12_LC_9_3_2  (
            .in0(N__25378),
            .in1(N__47220),
            .in2(N__24599),
            .in3(N__40849),
            .lcout(\ALU.a_15_m2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m4_bm_1_2_LC_9_3_3 .C_ON=1'b0;
    defparam \ALU.a_15_m4_bm_1_2_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m4_bm_1_2_LC_9_3_3 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \ALU.a_15_m4_bm_1_2_LC_9_3_3  (
            .in0(N__24595),
            .in1(N__47210),
            .in2(_gnd_net_),
            .in3(N__43899),
            .lcout(),
            .ltout(\ALU.a_15_m4_bm_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIII58A_2_LC_9_3_4 .C_ON=1'b0;
    defparam \ALU.d_RNIII58A_2_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIII58A_2_LC_9_3_4 .LUT_INIT=16'b0110011110000110;
    LogicCell40 \ALU.d_RNIII58A_2_LC_9_3_4  (
            .in0(N__47211),
            .in1(N__36937),
            .in2(N__24833),
            .in3(N__37256),
            .lcout(\ALU.d_RNIII58AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNITBSF7_3_LC_9_3_5 .C_ON=1'b0;
    defparam \ALU.d_RNITBSF7_3_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNITBSF7_3_LC_9_3_5 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \ALU.d_RNITBSF7_3_LC_9_3_5  (
            .in0(N__36936),
            .in1(N__39005),
            .in2(N__43727),
            .in3(N__42014),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI870EE_5_LC_9_3_6 .C_ON=1'b0;
    defparam \ALU.d_RNI870EE_5_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI870EE_5_LC_9_3_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI870EE_5_LC_9_3_6  (
            .in0(N__39006),
            .in1(N__40429),
            .in2(N__24821),
            .in3(N__42998),
            .lcout(\ALU.N_470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIFE9GA_0_LC_9_3_7 .C_ON=1'b0;
    defparam \ALU.d_RNIFE9GA_0_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIFE9GA_0_LC_9_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIFE9GA_0_LC_9_3_7  (
            .in0(N__38974),
            .in1(N__27235),
            .in2(_gnd_net_),
            .in3(N__24809),
            .lcout(\ALU.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI3DJU7_14_LC_9_4_0 .C_ON=1'b0;
    defparam \ALU.c_RNI3DJU7_14_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI3DJU7_14_LC_9_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNI3DJU7_14_LC_9_4_0  (
            .in0(N__43676),
            .in1(N__40627),
            .in2(_gnd_net_),
            .in3(N__40747),
            .lcout(\ALU.N_589 ),
            .ltout(\ALU.N_589_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI72MIC_0_15_LC_9_4_1 .C_ON=1'b0;
    defparam \ALU.c_RNI72MIC_0_15_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI72MIC_0_15_LC_9_4_1 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ALU.c_RNI72MIC_0_15_LC_9_4_1  (
            .in0(N__39017),
            .in1(N__38730),
            .in2(N__24797),
            .in3(N__30478),
            .lcout(),
            .ltout(\ALU.rshift_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI6PLSH_13_LC_9_4_2 .C_ON=1'b0;
    defparam \ALU.c_RNI6PLSH_13_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI6PLSH_13_LC_9_4_2 .LUT_INIT=16'b0001000111010001;
    LogicCell40 \ALU.c_RNI6PLSH_13_LC_9_4_2  (
            .in0(N__25235),
            .in1(N__43150),
            .in2(N__24794),
            .in3(N__44518),
            .lcout(\ALU.a_15_m3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI6KSGG_11_LC_9_4_3 .C_ON=1'b0;
    defparam \ALU.c_RNI6KSGG_11_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI6KSGG_11_LC_9_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNI6KSGG_11_LC_9_4_3  (
            .in0(N__39016),
            .in1(N__30495),
            .in2(_gnd_net_),
            .in3(N__25241),
            .lcout(\ALU.N_576 ),
            .ltout(\ALU.N_576_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIA9V4L_0_15_LC_9_4_4 .C_ON=1'b0;
    defparam \ALU.c_RNIA9V4L_0_15_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIA9V4L_0_15_LC_9_4_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ALU.c_RNIA9V4L_0_15_LC_9_4_4  (
            .in0(N__30479),
            .in1(N__38731),
            .in2(N__24779),
            .in3(N__39018),
            .lcout(),
            .ltout(\ALU.N_636_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNILI6TQ_11_LC_9_4_5 .C_ON=1'b0;
    defparam \ALU.c_RNILI6TQ_11_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNILI6TQ_11_LC_9_4_5 .LUT_INIT=16'b0100000001110011;
    LogicCell40 \ALU.c_RNILI6TQ_11_LC_9_4_5  (
            .in0(N__44519),
            .in1(N__43151),
            .in2(N__25418),
            .in3(N__25415),
            .lcout(\ALU.a_15_m3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIT87FA1_7_LC_9_4_6 .C_ON=1'b0;
    defparam \ALU.d_RNIT87FA1_7_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIT87FA1_7_LC_9_4_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \ALU.d_RNIT87FA1_7_LC_9_4_6  (
            .in0(N__43152),
            .in1(N__27383),
            .in2(_gnd_net_),
            .in3(N__25394),
            .lcout(\ALU.d_RNIT87FA1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIID898_11_LC_9_4_7 .C_ON=1'b0;
    defparam \ALU.c_RNIID898_11_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIID898_11_LC_9_4_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.c_RNIID898_11_LC_9_4_7  (
            .in0(N__43707),
            .in1(N__39390),
            .in2(_gnd_net_),
            .in3(N__25377),
            .lcout(\ALU.N_462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI5RLE5_13_LC_9_5_0 .C_ON=1'b0;
    defparam \ALU.d_RNI5RLE5_13_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI5RLE5_13_LC_9_5_0 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \ALU.d_RNI5RLE5_13_LC_9_5_0  (
            .in0(N__25010),
            .in1(_gnd_net_),
            .in2(N__26601),
            .in3(N__25039),
            .lcout(\ALU.N_177_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIURPF4_13_LC_9_5_1 .C_ON=1'b0;
    defparam \ALU.c_RNIURPF4_13_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIURPF4_13_LC_9_5_1 .LUT_INIT=16'b1111000011110101;
    LogicCell40 \ALU.c_RNIURPF4_13_LC_9_5_1  (
            .in0(N__40752),
            .in1(_gnd_net_),
            .in2(N__25052),
            .in3(N__29412),
            .lcout(\ALU.N_270_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m174_LC_9_5_2 .C_ON=1'b0;
    defparam \ALU.m174_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.m174_LC_9_5_2 .LUT_INIT=16'b1110111001111111;
    LogicCell40 \ALU.m174_LC_9_5_2  (
            .in0(N__30211),
            .in1(N__25204),
            .in2(N__30238),
            .in3(N__29741),
            .lcout(\ALU.N_175_0 ),
            .ltout(\ALU.N_175_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISHKD9_13_LC_9_5_3 .C_ON=1'b0;
    defparam \ALU.d_RNISHKD9_13_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISHKD9_13_LC_9_5_3 .LUT_INIT=16'b0110101001011001;
    LogicCell40 \ALU.d_RNISHKD9_13_LC_9_5_3  (
            .in0(N__40751),
            .in1(N__26553),
            .in2(N__25013),
            .in3(N__25009),
            .lcout(),
            .ltout(\ALU.un2_addsub_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9FOTE_13_LC_9_5_4 .C_ON=1'b0;
    defparam \ALU.d_RNI9FOTE_13_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9FOTE_13_LC_9_5_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \ALU.d_RNI9FOTE_13_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24980),
            .in3(N__24977),
            .lcout(\ALU.d_RNI9FOTEZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEG675_11_LC_9_5_5 .C_ON=1'b0;
    defparam \ALU.d_RNIEG675_11_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEG675_11_LC_9_5_5 .LUT_INIT=16'b0101111100110011;
    LogicCell40 \ALU.d_RNIEG675_11_LC_9_5_5  (
            .in0(N__24905),
            .in1(N__31181),
            .in2(N__29438),
            .in3(N__26554),
            .lcout(\ALU.N_186_0_i ),
            .ltout(\ALU.N_186_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIA7OEE_11_LC_9_5_6 .C_ON=1'b0;
    defparam \ALU.c_RNIA7OEE_11_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIA7OEE_11_LC_9_5_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \ALU.c_RNIA7OEE_11_LC_9_5_6  (
            .in0(N__39388),
            .in1(_gnd_net_),
            .in2(N__25574),
            .in3(N__39472),
            .lcout(\ALU.c_RNIA7OEEZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_29_LC_9_5_7.C_ON=1'b0;
    defparam testWord_29_LC_9_5_7.SEQ_MODE=4'b1000;
    defparam testWord_29_LC_9_5_7.LUT_INIT=16'b1111011110000000;
    LogicCell40 testWord_29_LC_9_5_7 (
            .in0(N__41359),
            .in1(N__41214),
            .in2(N__25556),
            .in3(N__30234),
            .lcout(ctrlOut_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47625),
            .ce(N__41062),
            .sr(_gnd_net_));
    defparam \ALU.h_12_LC_9_6_0 .C_ON=1'b0;
    defparam \ALU.h_12_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_12_LC_9_6_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.h_12_LC_9_6_0  (
            .in0(N__48436),
            .in1(N__34076),
            .in2(N__45991),
            .in3(N__34030),
            .lcout(\ALU.hZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47632),
            .ce(N__45498),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIFPBO_12_LC_9_6_1 .C_ON=1'b0;
    defparam \ALU.a_RNIFPBO_12_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIFPBO_12_LC_9_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_RNIFPBO_12_LC_9_6_1  (
            .in0(N__45126),
            .in1(N__28561),
            .in2(_gnd_net_),
            .in3(N__28207),
            .lcout(\ALU.a_RNIFPBOZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIM5LU_12_LC_9_6_2 .C_ON=1'b0;
    defparam \ALU.d_RNIM5LU_12_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIM5LU_12_LC_9_6_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNIM5LU_12_LC_9_6_2  (
            .in0(N__25492),
            .in1(N__45333),
            .in2(_gnd_net_),
            .in3(N__28390),
            .lcout(\ALU.d_RNIM5LUZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJ949_12_LC_9_6_3 .C_ON=1'b0;
    defparam \ALU.c_RNIJ949_12_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJ949_12_LC_9_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIJ949_12_LC_9_6_3  (
            .in0(N__45127),
            .in1(N__33958),
            .in2(_gnd_net_),
            .in3(N__31282),
            .lcout(),
            .ltout(\ALU.c_RNIJ949Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI693U1_12_LC_9_6_4 .C_ON=1'b0;
    defparam \ALU.c_RNI693U1_12_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI693U1_12_LC_9_6_4 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \ALU.c_RNI693U1_12_LC_9_6_4  (
            .in0(N__33084),
            .in1(N__34494),
            .in2(N__25481),
            .in3(N__25478),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI05RP4_12_LC_9_6_5 .C_ON=1'b0;
    defparam \ALU.d_RNI05RP4_12_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI05RP4_12_LC_9_6_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNI05RP4_12_LC_9_6_5  (
            .in0(N__32991),
            .in1(N__25472),
            .in2(N__25466),
            .in3(N__28328),
            .lcout(\ALU.operand2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7GCMD22_8_LC_9_7_0 .C_ON=1'b0;
    defparam \ALU.d_RNI7GCMD22_8_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7GCMD22_8_LC_9_7_0 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ALU.d_RNI7GCMD22_8_LC_9_7_0  (
            .in0(N__25664),
            .in1(N__26108),
            .in2(N__45989),
            .in3(N__26132),
            .lcout(\ALU.d_RNI7GCMD22Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPCSJD1_8_LC_9_7_1 .C_ON=1'b0;
    defparam \ALU.d_RNIPCSJD1_8_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPCSJD1_8_LC_9_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIPCSJD1_8_LC_9_7_1  (
            .in0(N__44187),
            .in1(N__25712),
            .in2(_gnd_net_),
            .in3(N__25697),
            .lcout(),
            .ltout(\ALU.a_15_m4_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIM0ETK2_8_LC_9_7_2 .C_ON=1'b0;
    defparam \ALU.d_RNIM0ETK2_8_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIM0ETK2_8_LC_9_7_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.d_RNIM0ETK2_8_LC_9_7_2  (
            .in0(N__25685),
            .in1(_gnd_net_),
            .in2(N__25667),
            .in3(N__46394),
            .lcout(\ALU.a_15_m5_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIRM7O_8_LC_9_7_3 .C_ON=1'b0;
    defparam \ALU.f_RNIRM7O_8_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIRM7O_8_LC_9_7_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.f_RNIRM7O_8_LC_9_7_3  (
            .in0(N__47720),
            .in1(N__31043),
            .in2(N__25658),
            .in3(N__45122),
            .lcout(),
            .ltout(\ALU.operand2_6_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQU7D1_8_LC_9_7_4 .C_ON=1'b0;
    defparam \ALU.d_RNIQU7D1_8_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQU7D1_8_LC_9_7_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIQU7D1_8_LC_9_7_4  (
            .in0(N__25585),
            .in1(N__25627),
            .in2(N__25607),
            .in3(N__34496),
            .lcout(\ALU.N_867 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_8_LC_9_7_5 .C_ON=1'b0;
    defparam \ALU.h_8_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \ALU.h_8_LC_9_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.h_8_LC_9_7_5  (
            .in0(N__48434),
            .in1(N__47864),
            .in2(_gnd_net_),
            .in3(N__47756),
            .lcout(\ALU.hZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47638),
            .ce(N__45525),
            .sr(_gnd_net_));
    defparam \ALU.f_10_LC_9_8_0 .C_ON=1'b0;
    defparam \ALU.f_10_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \ALU.f_10_LC_9_8_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.f_10_LC_9_8_0  (
            .in0(N__48635),
            .in1(N__34310),
            .in2(N__46076),
            .in3(N__34404),
            .lcout(\ALU.fZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__36376),
            .sr(_gnd_net_));
    defparam \ALU.f_11_LC_9_8_1 .C_ON=1'b0;
    defparam \ALU.f_11_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \ALU.f_11_LC_9_8_1 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.f_11_LC_9_8_1  (
            .in0(N__48638),
            .in1(N__34245),
            .in2(N__46080),
            .in3(N__34174),
            .lcout(\ALU.fZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__36376),
            .sr(_gnd_net_));
    defparam \ALU.f_12_LC_9_8_2 .C_ON=1'b0;
    defparam \ALU.f_12_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \ALU.f_12_LC_9_8_2 .LUT_INIT=16'b0111010101000101;
    LogicCell40 \ALU.f_12_LC_9_8_2  (
            .in0(N__34086),
            .in1(N__48641),
            .in2(N__46077),
            .in3(N__34021),
            .lcout(\ALU.fZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__36376),
            .sr(_gnd_net_));
    defparam \ALU.f_14_LC_9_8_3 .C_ON=1'b0;
    defparam \ALU.f_14_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \ALU.f_14_LC_9_8_3 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.f_14_LC_9_8_3  (
            .in0(N__48640),
            .in1(N__33816),
            .in2(N__46082),
            .in3(N__33749),
            .lcout(\ALU.fZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__36376),
            .sr(_gnd_net_));
    defparam \ALU.f_15_LC_9_8_4 .C_ON=1'b0;
    defparam \ALU.f_15_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \ALU.f_15_LC_9_8_4 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \ALU.f_15_LC_9_8_4  (
            .in0(N__48636),
            .in1(N__33655),
            .in2(N__46078),
            .in3(N__33602),
            .lcout(\ALU.fZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__36376),
            .sr(_gnd_net_));
    defparam \ALU.f_13_LC_9_8_5 .C_ON=1'b0;
    defparam \ALU.f_13_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \ALU.f_13_LC_9_8_5 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.f_13_LC_9_8_5  (
            .in0(N__48639),
            .in1(N__33935),
            .in2(N__46081),
            .in3(N__33873),
            .lcout(\ALU.fZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__36376),
            .sr(_gnd_net_));
    defparam \ALU.f_9_LC_9_8_6 .C_ON=1'b0;
    defparam \ALU.f_9_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \ALU.f_9_LC_9_8_6 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.f_9_LC_9_8_6  (
            .in0(N__48637),
            .in1(N__36268),
            .in2(N__46079),
            .in3(N__36194),
            .lcout(\ALU.fZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__36376),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_0_0_c_LC_9_9_0 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_0_0_c_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_0_0_c_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU.mult_madd_cry_0_0_c_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__25892),
            .in2(N__36662),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\ALU.madd_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_1_0_s_LC_9_9_1 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_1_0_s_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_1_0_s_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_1_0_s_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__33113),
            .in2(N__25877),
            .in3(N__25856),
            .lcout(\ALU.mult_2 ),
            .ltout(),
            .carryin(\ALU.madd_cry_0 ),
            .carryout(\ALU.madd_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_2_s_LC_9_9_2 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_2_s_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_2_s_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_2_s_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__25853),
            .in2(N__25831),
            .in3(N__25796),
            .lcout(\ALU.mult_3 ),
            .ltout(),
            .carryin(\ALU.madd_cry_1 ),
            .carryout(\ALU.madd_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_3_s_LC_9_9_3 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_3_s_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_3_s_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_3_s_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__25793),
            .in2(N__25781),
            .in3(N__25760),
            .lcout(\ALU.mult_4 ),
            .ltout(),
            .carryin(\ALU.madd_cry_2 ),
            .carryout(\ALU.madd_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_4_s_LC_9_9_4 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_4_s_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_4_s_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_4_s_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__25757),
            .in2(N__25742),
            .in3(N__25715),
            .lcout(\ALU.mult_5 ),
            .ltout(),
            .carryin(\ALU.madd_cry_3 ),
            .carryout(\ALU.madd_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_5_s_LC_9_9_5 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_5_s_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_5_s_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_5_s_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__26179),
            .in2(N__26159),
            .in3(N__26138),
            .lcout(\ALU.mult_6 ),
            .ltout(),
            .carryin(\ALU.madd_cry_4 ),
            .carryout(\ALU.madd_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_5_THRU_LUT4_0_LC_9_9_6 .C_ON=1'b1;
    defparam \ALU.madd_cry_5_THRU_LUT4_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_5_THRU_LUT4_0_LC_9_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_5_THRU_LUT4_0_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__42349),
            .in2(_gnd_net_),
            .in3(N__26135),
            .lcout(\ALU.madd_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ALU.madd_cry_5 ),
            .carryout(\ALU.madd_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.madd_cry_6_THRU_LUT4_0_LC_9_9_7 .C_ON=1'b1;
    defparam \ALU.madd_cry_6_THRU_LUT4_0_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.madd_cry_6_THRU_LUT4_0_LC_9_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ALU.madd_cry_6_THRU_LUT4_0_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__26128),
            .in2(_gnd_net_),
            .in3(N__26099),
            .lcout(\ALU.madd_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ALU.madd_cry_6 ),
            .carryout(\ALU.madd_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_8_s_LC_9_10_0 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_8_s_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_8_s_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_8_s_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__26096),
            .in2(N__26078),
            .in3(N__26054),
            .lcout(\ALU.mult_9 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\ALU.madd_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_9_0_s_LC_9_10_1 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_9_0_s_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_9_0_s_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_9_0_s_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__26051),
            .in2(N__26039),
            .in3(N__26018),
            .lcout(\ALU.mult_10 ),
            .ltout(),
            .carryin(\ALU.madd_cry_8 ),
            .carryout(\ALU.madd_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_10_0_s_LC_9_10_2 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_10_0_s_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_10_0_s_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_10_0_s_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__26015),
            .in2(N__25997),
            .in3(N__25982),
            .lcout(\ALU.mult_11 ),
            .ltout(),
            .carryin(\ALU.madd_cry_9 ),
            .carryout(\ALU.madd_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_11_s_LC_9_10_3 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_11_s_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_11_s_LC_9_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ALU.mult_madd_cry_11_s_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25979),
            .in3(N__25964),
            .lcout(\ALU.mult_12 ),
            .ltout(),
            .carryin(\ALU.madd_cry_10 ),
            .carryout(\ALU.madd_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_12_s_LC_9_10_4 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_12_s_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_12_s_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_12_s_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__25961),
            .in2(N__25943),
            .in3(N__25919),
            .lcout(\ALU.mult_13 ),
            .ltout(),
            .carryin(\ALU.madd_cry_11 ),
            .carryout(\ALU.madd_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_cry_13_0_s_LC_9_10_5 .C_ON=1'b1;
    defparam \ALU.mult_madd_cry_13_0_s_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_cry_13_0_s_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.mult_madd_cry_13_0_s_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__26786),
            .in2(N__26771),
            .in3(N__26753),
            .lcout(\ALU.mult_14 ),
            .ltout(),
            .carryin(\ALU.madd_cry_12 ),
            .carryout(\ALU.madd_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_s_14_LC_9_10_6 .C_ON=1'b0;
    defparam \ALU.mult_madd_s_14_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_s_14_LC_9_10_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALU.mult_madd_s_14_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__26750),
            .in2(_gnd_net_),
            .in3(N__26735),
            .lcout(\ALU.mult_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3O5R3_6_LC_9_10_7 .C_ON=1'b0;
    defparam \ALU.d_RNI3O5R3_6_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3O5R3_6_LC_9_10_7 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ALU.d_RNI3O5R3_6_LC_9_10_7  (
            .in0(N__26728),
            .in1(N__26650),
            .in2(_gnd_net_),
            .in3(N__26253),
            .lcout(\ALU.N_219_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIS5U41_15_LC_9_11_0 .C_ON=1'b0;
    defparam \ALU.a_RNIS5U41_15_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIS5U41_15_LC_9_11_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.a_RNIS5U41_15_LC_9_11_0  (
            .in0(N__35871),
            .in1(N__31361),
            .in2(N__35554),
            .in3(N__31745),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI7JQF1_15_LC_9_11_1 .C_ON=1'b0;
    defparam \ALU.c_RNI7JQF1_15_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI7JQF1_15_LC_9_11_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.c_RNI7JQF1_15_LC_9_11_1  (
            .in0(N__35299),
            .in1(N__33539),
            .in2(N__26192),
            .in3(N__31523),
            .lcout(\ALU.N_714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_e_0_2_LC_9_11_2 .C_ON=1'b0;
    defparam \CONTROL.operand1_e_0_2_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_e_0_2_LC_9_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.operand1_e_0_2_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27195),
            .lcout(aluOperand1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47664),
            .ce(N__27723),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIM2101_2_LC_9_11_3 .C_ON=1'b0;
    defparam \ALU.f_RNIM2101_2_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIM2101_2_LC_9_11_3 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \ALU.f_RNIM2101_2_LC_9_11_3  (
            .in0(N__31963),
            .in1(N__35870),
            .in2(N__35531),
            .in3(N__36458),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIR8K91_2_LC_9_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNIR8K91_2_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIR8K91_2_LC_9_11_4 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \ALU.d_RNIR8K91_2_LC_9_11_4  (
            .in0(N__31427),
            .in1(N__35298),
            .in2(N__26189),
            .in3(N__42038),
            .lcout(),
            .ltout(\ALU.N_749_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6KCD3_2_LC_9_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNI6KCD3_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6KCD3_2_LC_9_11_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNI6KCD3_2_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__35202),
            .in2(N__26186),
            .in3(N__26918),
            .lcout(\ALU.aluOut_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNI70VV1_2_LC_9_11_6 .C_ON=1'b0;
    defparam \ALU.g_RNI70VV1_2_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNI70VV1_2_LC_9_11_6 .LUT_INIT=16'b1110010001010101;
    LogicCell40 \ALU.g_RNI70VV1_2_LC_9_11_6  (
            .in0(N__26912),
            .in1(N__31901),
            .in2(N__29096),
            .in3(N__35297),
            .lcout(\ALU.N_701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI40I81_2_LC_9_12_0 .C_ON=1'b0;
    defparam \ALU.e_RNI40I81_2_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI40I81_2_LC_9_12_0 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \ALU.e_RNI40I81_2_LC_9_12_0  (
            .in0(N__35853),
            .in1(N__28758),
            .in2(N__35966),
            .in3(N__28781),
            .lcout(\ALU.dout_3_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_2_rep2_e_LC_9_12_1 .C_ON=1'b0;
    defparam \CONTROL.operand1_2_rep2_e_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_2_rep2_e_LC_9_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.operand1_2_rep2_e_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27196),
            .lcout(aluOperand1_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47671),
            .ce(N__27719),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIGGOA1_7_LC_9_12_2 .C_ON=1'b0;
    defparam \ALU.f_RNIGGOA1_7_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIGGOA1_7_LC_9_12_2 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.f_RNIGGOA1_7_LC_9_12_2  (
            .in0(N__35852),
            .in1(N__36391),
            .in2(N__35965),
            .in3(N__48655),
            .lcout(\ALU.dout_6_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_1_rep1_e_LC_9_12_3 .C_ON=1'b0;
    defparam \CONTROL.operand1_1_rep1_e_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_1_rep1_e_LC_9_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \CONTROL.operand1_1_rep1_e_LC_9_12_3  (
            .in0(N__26879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(aluOperand1_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47671),
            .ce(N__27719),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIDCNA1_6_LC_9_12_4 .C_ON=1'b0;
    defparam \ALU.f_RNIDCNA1_6_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIDCNA1_6_LC_9_12_4 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.f_RNIDCNA1_6_LC_9_12_4  (
            .in0(N__27336),
            .in1(N__36415),
            .in2(N__35875),
            .in3(N__48811),
            .lcout(\ALU.dout_6_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIQQJ01_7_LC_9_12_5 .C_ON=1'b0;
    defparam \ALU.f_RNIQQJ01_7_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIQQJ01_7_LC_9_12_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.f_RNIQQJ01_7_LC_9_12_5  (
            .in0(N__48656),
            .in1(_gnd_net_),
            .in2(N__36395),
            .in3(N__45313),
            .lcout(\ALU.f_RNIQQJ01Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_e_0_1_LC_9_12_6 .C_ON=1'b0;
    defparam \CONTROL.operand1_e_0_1_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_e_0_1_LC_9_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.operand1_e_0_1_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26880),
            .lcout(aluOperand1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47671),
            .ce(N__27719),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIEHSD1_10_LC_9_12_7 .C_ON=1'b0;
    defparam \ALU.b_RNIEHSD1_10_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIEHSD1_10_LC_9_12_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.b_RNIEHSD1_10_LC_9_12_7  (
            .in0(N__26826),
            .in1(N__28518),
            .in2(_gnd_net_),
            .in3(N__45314),
            .lcout(\ALU.b_RNIEHSD1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_0_LC_9_13_0 .C_ON=1'b0;
    defparam \ALU.a_0_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \ALU.a_0_LC_9_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_0_LC_9_13_0  (
            .in0(N__48618),
            .in1(N__42311),
            .in2(_gnd_net_),
            .in3(N__42233),
            .lcout(a_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__44870),
            .sr(_gnd_net_));
    defparam \ALU.a_1_LC_9_13_1 .C_ON=1'b0;
    defparam \ALU.a_1_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \ALU.a_1_LC_9_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_1_LC_9_13_1  (
            .in0(N__48615),
            .in1(N__40994),
            .in2(_gnd_net_),
            .in3(N__36605),
            .lcout(a_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__44870),
            .sr(_gnd_net_));
    defparam \ALU.a_2_LC_9_13_2 .C_ON=1'b0;
    defparam \ALU.a_2_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.a_2_LC_9_13_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.a_2_LC_9_13_2  (
            .in0(N__42163),
            .in1(N__48616),
            .in2(_gnd_net_),
            .in3(N__42079),
            .lcout(a_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__44870),
            .sr(_gnd_net_));
    defparam \ALU.a_4_LC_9_13_4 .C_ON=1'b0;
    defparam \ALU.a_4_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \ALU.a_4_LC_9_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.a_4_LC_9_13_4  (
            .in0(N__49281),
            .in1(N__49220),
            .in2(_gnd_net_),
            .in3(N__48617),
            .lcout(a_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__44870),
            .sr(_gnd_net_));
    defparam \ALU.a_5_LC_9_13_5 .C_ON=1'b0;
    defparam \ALU.a_5_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \ALU.a_5_LC_9_13_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.a_5_LC_9_13_5  (
            .in0(N__49101),
            .in1(N__48620),
            .in2(_gnd_net_),
            .in3(N__49046),
            .lcout(a_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__44870),
            .sr(_gnd_net_));
    defparam \ALU.a_6_LC_9_13_6 .C_ON=1'b0;
    defparam \ALU.a_6_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \ALU.a_6_LC_9_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_6_LC_9_13_6  (
            .in0(N__48619),
            .in1(N__48891),
            .in2(_gnd_net_),
            .in3(N__48942),
            .lcout(a_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__44870),
            .sr(_gnd_net_));
    defparam \ALU.a_7_LC_9_13_7 .C_ON=1'b0;
    defparam \ALU.a_7_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \ALU.a_7_LC_9_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.a_7_LC_9_13_7  (
            .in0(N__48770),
            .in1(N__48716),
            .in2(_gnd_net_),
            .in3(N__48621),
            .lcout(a_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__44870),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI5J7N_4_LC_9_14_0 .C_ON=1'b0;
    defparam \ALU.e_RNI5J7N_4_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI5J7N_4_LC_9_14_0 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \ALU.e_RNI5J7N_4_LC_9_14_0  (
            .in0(N__27131),
            .in1(N__27924),
            .in2(N__27028),
            .in3(N__26959),
            .lcout(\ALU.dout_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_4_LC_9_14_1 .C_ON=1'b0;
    defparam \ALU.e_4_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.e_4_LC_9_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_4_LC_9_14_1  (
            .in0(N__48420),
            .in1(N__49286),
            .in2(_gnd_net_),
            .in3(N__49217),
            .lcout(\ALU.eZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47681),
            .ce(N__32444),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIS97J_1_LC_9_14_2 .C_ON=1'b0;
    defparam \ALU.e_RNIS97J_1_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIS97J_1_LC_9_14_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.e_RNIS97J_1_LC_9_14_2  (
            .in0(N__27011),
            .in1(N__44586),
            .in2(_gnd_net_),
            .in3(N__26932),
            .lcout(\ALU.e_RNIS97JZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_1_LC_9_14_3 .C_ON=1'b0;
    defparam \ALU.e_1_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.e_1_LC_9_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_1_LC_9_14_3  (
            .in0(N__48419),
            .in1(N__40998),
            .in2(_gnd_net_),
            .in3(N__36614),
            .lcout(\ALU.eZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47681),
            .ce(N__32444),
            .sr(_gnd_net_));
    defparam \ALU.g_RNI0MJN_1_LC_9_14_4 .C_ON=1'b0;
    defparam \ALU.g_RNI0MJN_1_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNI0MJN_1_LC_9_14_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ALU.g_RNI0MJN_1_LC_9_14_4  (
            .in0(N__29110),
            .in1(_gnd_net_),
            .in2(N__27027),
            .in3(N__31921),
            .lcout(\ALU.g_RNI0MJNZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIM1T31_3_LC_9_14_5 .C_ON=1'b0;
    defparam \ALU.f_RNIM1T31_3_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIM1T31_3_LC_9_14_5 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.f_RNIM1T31_3_LC_9_14_5  (
            .in0(N__27338),
            .in1(N__49310),
            .in2(N__43268),
            .in3(N__27130),
            .lcout(\ALU.dout_6_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIO3T31_4_LC_9_14_7 .C_ON=1'b0;
    defparam \ALU.f_RNIO3T31_4_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIO3T31_4_LC_9_14_7 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \ALU.f_RNIO3T31_4_LC_9_14_7  (
            .in0(N__27132),
            .in1(N__45410),
            .in2(N__27348),
            .in3(N__49151),
            .lcout(\ALU.dout_6_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIE5EP3_0_LC_9_15_0 .C_ON=1'b0;
    defparam \ALU.d_RNIE5EP3_0_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIE5EP3_0_LC_9_15_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \ALU.d_RNIE5EP3_0_LC_9_15_0  (
            .in0(N__27275),
            .in1(N__35135),
            .in2(N__43769),
            .in3(N__27263),
            .lcout(\ALU.N_404_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQQAK1_6_LC_9_15_1 .C_ON=1'b0;
    defparam \ALU.d_RNIQQAK1_6_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQQAK1_6_LC_9_15_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNIQQAK1_6_LC_9_15_1  (
            .in0(N__45623),
            .in1(N__43372),
            .in2(N__27212),
            .in3(N__35356),
            .lcout(),
            .ltout(\ALU.N_753_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI23RD3_6_LC_9_15_2 .C_ON=1'b0;
    defparam \ALU.d_RNI23RD3_6_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI23RD3_6_LC_9_15_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNI23RD3_6_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__35134),
            .in2(N__27200),
            .in3(N__27764),
            .lcout(\ALU.aluOut_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_fast_e_2_LC_9_15_3 .C_ON=1'b0;
    defparam \CONTROL.operand1_fast_e_2_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_fast_e_2_LC_9_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.operand1_fast_e_2_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27197),
            .lcout(aluOperand1_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47684),
            .ce(N__27728),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI9N7N_6_LC_9_15_4 .C_ON=1'b0;
    defparam \ALU.e_RNI9N7N_6_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI9N7N_6_LC_9_15_4 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \ALU.e_RNI9N7N_6_LC_9_15_4  (
            .in0(N__28621),
            .in1(N__27127),
            .in2(N__27026),
            .in3(N__27898),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNI4TML1_6_LC_9_15_5 .C_ON=1'b0;
    defparam \ALU.g_RNI4TML1_6_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNI4TML1_6_LC_9_15_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.g_RNI4TML1_6_LC_9_15_5  (
            .in0(N__35713),
            .in1(N__28976),
            .in2(N__27767),
            .in3(N__29011),
            .lcout(\ALU.N_705 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand1_e_0_0_LC_9_15_6 .C_ON=1'b0;
    defparam \CONTROL.operand1_e_0_0_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand1_e_0_0_LC_9_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \CONTROL.operand1_e_0_0_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27758),
            .lcout(aluOperand1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47684),
            .ce(N__27728),
            .sr(_gnd_net_));
    defparam \ALU.c_8_LC_10_1_0 .C_ON=1'b0;
    defparam \ALU.c_8_LC_10_1_0 .SEQ_MODE=4'b1000;
    defparam \ALU.c_8_LC_10_1_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_8_LC_10_1_0  (
            .in0(N__48074),
            .in1(N__47887),
            .in2(_gnd_net_),
            .in3(N__47798),
            .lcout(\ALU.cZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47600),
            .ce(N__31498),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_0_LC_10_2_2 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_0_LC_10_2_2 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_0_LC_10_2_2 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \FTDI.TXstate_RNO_0_0_LC_10_2_2  (
            .in0(N__29522),
            .in1(_gnd_net_),
            .in2(N__44749),
            .in3(N__30380),
            .lcout(\FTDI.TXstate_e_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI72MIC_15_LC_10_2_4 .C_ON=1'b0;
    defparam \ALU.c_RNI72MIC_15_LC_10_2_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI72MIC_15_LC_10_2_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \ALU.c_RNI72MIC_15_LC_10_2_4  (
            .in0(N__39022),
            .in1(N__30477),
            .in2(N__38734),
            .in3(N__30503),
            .lcout(),
            .ltout(\ALU.c_RNI72MICZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIBHJVC1_15_LC_10_2_5 .C_ON=1'b0;
    defparam \ALU.c_RNIBHJVC1_15_LC_10_2_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIBHJVC1_15_LC_10_2_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNIBHJVC1_15_LC_10_2_5  (
            .in0(_gnd_net_),
            .in1(N__44479),
            .in2(N__27620),
            .in3(N__27617),
            .lcout(\ALU.rshift_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_0_LC_10_2_6 .C_ON=1'b0;
    defparam \FTDI.baudAcc_0_LC_10_2_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_0_LC_10_2_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \FTDI.baudAcc_0_LC_10_2_6  (
            .in0(_gnd_net_),
            .in1(N__29586),
            .in2(_gnd_net_),
            .in3(N__30418),
            .lcout(\FTDI.baudAccZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6QT5G_9_LC_10_3_0 .C_ON=1'b0;
    defparam \ALU.d_RNI6QT5G_9_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6QT5G_9_LC_10_3_0 .LUT_INIT=16'b1101010110000101;
    LogicCell40 \ALU.d_RNI6QT5G_9_LC_10_3_0  (
            .in0(N__27809),
            .in1(N__39860),
            .in2(N__39084),
            .in3(N__27607),
            .lcout(\ALU.N_475 ),
            .ltout(\ALU.N_475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIGVM161_15_LC_10_3_1 .C_ON=1'b0;
    defparam \ALU.c_RNIGVM161_15_LC_10_3_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIGVM161_15_LC_10_3_1 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \ALU.c_RNIGVM161_15_LC_10_3_1  (
            .in0(N__44395),
            .in1(N__27827),
            .in2(N__27386),
            .in3(N__27803),
            .lcout(\ALU.rshift_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI4JFV4_15_LC_10_3_2 .C_ON=1'b0;
    defparam \ALU.c_RNI4JFV4_15_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI4JFV4_15_LC_10_3_2 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \ALU.c_RNI4JFV4_15_LC_10_3_2  (
            .in0(N__30469),
            .in1(N__44394),
            .in2(N__38714),
            .in3(N__39011),
            .lcout(\ALU.rshift_15_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI83IG7_0_3_LC_10_3_3 .C_ON=1'b0;
    defparam \ALU.d_RNI83IG7_0_3_LC_10_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI83IG7_0_3_LC_10_3_3 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \ALU.d_RNI83IG7_0_3_LC_10_3_3  (
            .in0(N__43690),
            .in1(N__42013),
            .in2(N__39069),
            .in3(N__42991),
            .lcout(),
            .ltout(\ALU.rshift_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4MEEE_6_LC_10_3_4 .C_ON=1'b0;
    defparam \ALU.d_RNI4MEEE_6_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4MEEE_6_LC_10_3_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \ALU.d_RNI4MEEE_6_LC_10_3_4  (
            .in0(N__39061),
            .in1(N__40428),
            .in2(N__27821),
            .in3(N__46716),
            .lcout(),
            .ltout(\ALU.N_471_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI9DPVU_6_LC_10_3_5 .C_ON=1'b0;
    defparam \ALU.d_RNI9DPVU_6_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI9DPVU_6_LC_10_3_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNI9DPVU_6_LC_10_3_5  (
            .in0(_gnd_net_),
            .in1(N__38648),
            .in2(N__27818),
            .in3(N__27815),
            .lcout(\ALU.d_RNI9DPVUZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIT1MQ7_7_LC_10_3_6 .C_ON=1'b0;
    defparam \ALU.d_RNIT1MQ7_7_LC_10_3_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIT1MQ7_7_LC_10_3_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \ALU.d_RNIT1MQ7_7_LC_10_3_6  (
            .in0(N__43689),
            .in1(N__40119),
            .in2(N__39083),
            .in3(N__46975),
            .lcout(\ALU.rshift_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIA9V4L_15_LC_10_3_7 .C_ON=1'b0;
    defparam \ALU.c_RNIA9V4L_15_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIA9V4L_15_LC_10_3_7 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ALU.c_RNIA9V4L_15_LC_10_3_7  (
            .in0(N__39010),
            .in1(N__30470),
            .in2(N__38715),
            .in3(N__27802),
            .lcout(\ALU.c_RNIA9V4LZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6I9AJ2_5_LC_10_4_0 .C_ON=1'b0;
    defparam \ALU.d_RNI6I9AJ2_5_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6I9AJ2_5_LC_10_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNI6I9AJ2_5_LC_10_4_0  (
            .in0(N__46363),
            .in1(N__27947),
            .in2(_gnd_net_),
            .in3(N__29528),
            .lcout(),
            .ltout(\ALU.a_15_m5_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIH1NE6F_5_LC_10_4_1 .C_ON=1'b0;
    defparam \ALU.d_RNIH1NE6F_5_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIH1NE6F_5_LC_10_4_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIH1NE6F_5_LC_10_4_1  (
            .in0(_gnd_net_),
            .in1(N__45923),
            .in2(N__27794),
            .in3(N__27791),
            .lcout(\ALU.d_RNIH1NE6FZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIRCOSL2_9_LC_10_4_2 .C_ON=1'b0;
    defparam \ALU.d_RNIRCOSL2_9_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIRCOSL2_9_LC_10_4_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNIRCOSL2_9_LC_10_4_2  (
            .in0(N__46362),
            .in1(N__30428),
            .in2(_gnd_net_),
            .in3(N__27776),
            .lcout(\ALU.a_15_m5_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_5_LC_10_4_3 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_5_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_5_LC_10_4_3 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.a_15_m2_ns_1_5_LC_10_4_3  (
            .in0(N__47178),
            .in1(N__44151),
            .in2(N__43929),
            .in3(N__43726),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISQNAA_5_LC_10_4_4 .C_ON=1'b0;
    defparam \ALU.d_RNISQNAA_5_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISQNAA_5_LC_10_4_4 .LUT_INIT=16'b1000011001100111;
    LogicCell40 \ALU.d_RNISQNAA_5_LC_10_4_4  (
            .in0(N__47179),
            .in1(N__40401),
            .in2(N__28100),
            .in3(N__28097),
            .lcout(),
            .ltout(\ALU.a_15_m2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQO6O01_5_LC_10_4_5 .C_ON=1'b0;
    defparam \ALU.d_RNIQO6O01_5_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQO6O01_5_LC_10_4_5 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \ALU.d_RNIQO6O01_5_LC_10_4_5  (
            .in0(N__44500),
            .in1(N__44152),
            .in2(N__27968),
            .in3(N__27965),
            .lcout(\ALU.a_15_m4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXbuffer_0_LC_10_5_0.C_ON=1'b0;
    defparam TXbuffer_0_LC_10_5_0.SEQ_MODE=4'b1000;
    defparam TXbuffer_0_LC_10_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_0_LC_10_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28937),
            .lcout(TXbufferZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47613),
            .ce(N__44551),
            .sr(_gnd_net_));
    defparam TXbuffer_2_LC_10_5_2.C_ON=1'b0;
    defparam TXbuffer_2_LC_10_5_2.SEQ_MODE=4'b1000;
    defparam TXbuffer_2_LC_10_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_2_LC_10_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28769),
            .lcout(TXbufferZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47613),
            .ce(N__44551),
            .sr(_gnd_net_));
    defparam TXbuffer_3_LC_10_5_3.C_ON=1'b0;
    defparam TXbuffer_3_LC_10_5_3.SEQ_MODE=4'b1000;
    defparam TXbuffer_3_LC_10_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_3_LC_10_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44915),
            .lcout(TXbufferZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47613),
            .ce(N__44551),
            .sr(_gnd_net_));
    defparam TXbuffer_4_LC_10_5_4.C_ON=1'b0;
    defparam TXbuffer_4_LC_10_5_4.SEQ_MODE=4'b1000;
    defparam TXbuffer_4_LC_10_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_4_LC_10_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27940),
            .lcout(TXbufferZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47613),
            .ce(N__44551),
            .sr(_gnd_net_));
    defparam TXbuffer_6_LC_10_5_6.C_ON=1'b0;
    defparam TXbuffer_6_LC_10_5_6.SEQ_MODE=4'b1000;
    defparam TXbuffer_6_LC_10_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_6_LC_10_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27908),
            .lcout(TXbufferZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47613),
            .ce(N__44551),
            .sr(_gnd_net_));
    defparam TXbuffer_7_LC_10_5_7.C_ON=1'b0;
    defparam TXbuffer_7_LC_10_5_7.SEQ_MODE=4'b1000;
    defparam TXbuffer_7_LC_10_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_7_LC_10_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27874),
            .lcout(TXbufferZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47613),
            .ce(N__44551),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI1BC602_12_LC_10_6_0 .C_ON=1'b0;
    defparam \ALU.c_RNI1BC602_12_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI1BC602_12_LC_10_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNI1BC602_12_LC_10_6_0  (
            .in0(N__44228),
            .in1(N__27836),
            .in2(_gnd_net_),
            .in3(N__28166),
            .lcout(),
            .ltout(\ALU.a_15_m4_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIC8RDN2_12_LC_10_6_1 .C_ON=1'b0;
    defparam \ALU.c_RNIC8RDN2_12_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIC8RDN2_12_LC_10_6_1 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \ALU.c_RNIC8RDN2_12_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__46383),
            .in2(N__28238),
            .in3(N__28187),
            .lcout(c_RNIC8RDN2_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_11_c_RNIQ9LMU_LC_10_6_2 .C_ON=1'b0;
    defparam \ALU.un2_addsub_cry_11_c_RNIQ9LMU_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_11_c_RNIQ9LMU_LC_10_6_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ALU.un2_addsub_cry_11_c_RNIQ9LMU_LC_10_6_2  (
            .in0(N__42459),
            .in1(N__40787),
            .in2(_gnd_net_),
            .in3(N__28235),
            .lcout(),
            .ltout(un2_addsub_cry_11_c_RNIQ9LMU_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_RNIGPL5M3_0_LC_10_6_3 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_RNIGPL5M3_0_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_RNIGPL5M3_0_LC_10_6_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \CONTROL.aluOperation_RNIGPL5M3_0_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__48339),
            .in2(N__28223),
            .in3(N__28220),
            .lcout(aluOperation_RNIGPL5M3_0),
            .ltout(aluOperation_RNIGPL5M3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_12_LC_10_6_4 .C_ON=1'b0;
    defparam \ALU.a_12_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \ALU.a_12_LC_10_6_4 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.a_12_LC_10_6_4  (
            .in0(N__48340),
            .in1(N__45836),
            .in2(N__28214),
            .in3(N__34031),
            .lcout(\ALU.aZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47619),
            .ce(N__44849),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIC6T9M_12_LC_10_6_5 .C_ON=1'b0;
    defparam \ALU.c_RNIC6T9M_12_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIC6T9M_12_LC_10_6_5 .LUT_INIT=16'b0101001100000011;
    LogicCell40 \ALU.c_RNIC6T9M_12_LC_10_6_5  (
            .in0(N__44437),
            .in1(N__28196),
            .in2(N__43189),
            .in3(N__43231),
            .lcout(\ALU.a_15_m3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI6VHRI1_0_LC_10_6_6 .C_ON=1'b0;
    defparam \ALU.d_RNI6VHRI1_0_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI6VHRI1_0_LC_10_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNI6VHRI1_0_LC_10_6_6  (
            .in0(N__44520),
            .in1(N__44959),
            .in2(_gnd_net_),
            .in3(N__28181),
            .lcout(\ALU.lshift_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_m2_1_0_LC_10_7_0 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_m2_1_0_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_m2_1_0_LC_10_7_0 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.mult_g0_0_0_m2_1_0_LC_10_7_0  (
            .in0(N__45281),
            .in1(N__28126),
            .in2(N__28159),
            .in3(N__35033),
            .lcout(\ALU.g0_0_0_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_9_LC_10_7_1 .C_ON=1'b0;
    defparam \ALU.b_9_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \ALU.b_9_LC_10_7_1 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.b_9_LC_10_7_1  (
            .in0(N__48435),
            .in1(N__36257),
            .in2(N__46084),
            .in3(N__36204),
            .lcout(\ALU.bZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47626),
            .ce(N__47393),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIUUJ01_9_LC_10_7_2 .C_ON=1'b0;
    defparam \ALU.f_RNIUUJ01_9_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIUUJ01_9_LC_10_7_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.f_RNIUUJ01_9_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__45284),
            .in2(N__28158),
            .in3(N__28125),
            .lcout(\ALU.f_RNIUUJ01Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_11_LC_10_7_3 .C_ON=1'b0;
    defparam \ALU.b_11_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \ALU.b_11_LC_10_7_3 .LUT_INIT=16'b0111010101000101;
    LogicCell40 \ALU.b_11_LC_10_7_3  (
            .in0(N__34246),
            .in1(N__48411),
            .in2(N__46083),
            .in3(N__34175),
            .lcout(\ALU.bZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47626),
            .ce(N__47393),
            .sr(_gnd_net_));
    defparam \ALU.b_12_LC_10_7_4 .C_ON=1'b0;
    defparam \ALU.b_12_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \ALU.b_12_LC_10_7_4 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.b_12_LC_10_7_4  (
            .in0(N__48409),
            .in1(N__45993),
            .in2(N__34088),
            .in3(N__34026),
            .lcout(\ALU.bZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47626),
            .ce(N__47393),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIILSD1_12_LC_10_7_5 .C_ON=1'b0;
    defparam \ALU.b_RNIILSD1_12_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIILSD1_12_LC_10_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.b_RNIILSD1_12_LC_10_7_5  (
            .in0(N__45283),
            .in1(N__28363),
            .in2(_gnd_net_),
            .in3(N__28342),
            .lcout(\ALU.b_RNIILSD1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_14_LC_10_7_6 .C_ON=1'b0;
    defparam \ALU.b_14_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \ALU.b_14_LC_10_7_6 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.b_14_LC_10_7_6  (
            .in0(N__48410),
            .in1(N__33815),
            .in2(N__46118),
            .in3(N__33756),
            .lcout(\ALU.bZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47626),
            .ce(N__47393),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIMPSD1_14_LC_10_7_7 .C_ON=1'b0;
    defparam \ALU.b_RNIMPSD1_14_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIMPSD1_14_LC_10_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.b_RNIMPSD1_14_LC_10_7_7  (
            .in0(N__28309),
            .in1(N__28288),
            .in2(_gnd_net_),
            .in3(N__45282),
            .lcout(\ALU.b_RNIMPSD1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI8DRP4_13_LC_10_8_0 .C_ON=1'b0;
    defparam \ALU.d_RNI8DRP4_13_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI8DRP4_13_LC_10_8_0 .LUT_INIT=16'b0111011100001010;
    LogicCell40 \ALU.d_RNI8DRP4_13_LC_10_8_0  (
            .in0(N__32983),
            .in1(N__28256),
            .in2(N__28250),
            .in3(N__31096),
            .lcout(),
            .ltout(\ALU.g0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIA7959_13_LC_10_8_1 .C_ON=1'b0;
    defparam \ALU.d_RNIA7959_13_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIA7959_13_LC_10_8_1 .LUT_INIT=16'b1010101100000000;
    LogicCell40 \ALU.d_RNIA7959_13_LC_10_8_1  (
            .in0(N__29612),
            .in1(N__29966),
            .in2(N__28277),
            .in3(N__38041),
            .lcout(\ALU.N_703_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIKNSD1_0_13_LC_10_8_2 .C_ON=1'b0;
    defparam \ALU.b_RNIKNSD1_0_13_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIKNSD1_0_13_LC_10_8_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.b_RNIKNSD1_0_13_LC_10_8_2  (
            .in0(N__45279),
            .in1(_gnd_net_),
            .in2(N__35614),
            .in3(N__35783),
            .lcout(\ALU.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO7LU_0_13_LC_10_8_3 .C_ON=1'b0;
    defparam \ALU.d_RNIO7LU_0_13_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO7LU_0_13_LC_10_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.d_RNIO7LU_0_13_LC_10_8_3  (
            .in0(N__35424),
            .in1(N__35461),
            .in2(_gnd_net_),
            .in3(N__45278),
            .lcout(\ALU.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_2_LC_10_8_5 .C_ON=1'b0;
    defparam \CONTROL.operand2_2_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_2_LC_10_8_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \CONTROL.operand2_2_LC_10_8_5  (
            .in0(N__34799),
            .in1(N__32213),
            .in2(N__34721),
            .in3(N__45280),
            .lcout(aluOperand2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47633),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIGJSD1_11_LC_10_8_6 .C_ON=1'b0;
    defparam \ALU.b_RNIGJSD1_11_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIGJSD1_11_LC_10_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_RNIGJSD1_11_LC_10_8_6  (
            .in0(N__45276),
            .in1(N__28468),
            .in2(_gnd_net_),
            .in3(N__28450),
            .lcout(\ALU.b_RNIGJSD1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIKNSD1_13_LC_10_8_7 .C_ON=1'b0;
    defparam \ALU.b_RNIKNSD1_13_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIKNSD1_13_LC_10_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.b_RNIKNSD1_13_LC_10_8_7  (
            .in0(N__35782),
            .in1(N__35607),
            .in2(_gnd_net_),
            .in3(N__45277),
            .lcout(\ALU.b_RNIKNSD1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_10_LC_10_9_0 .C_ON=1'b0;
    defparam \ALU.d_10_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \ALU.d_10_LC_10_9_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.d_10_LC_10_9_0  (
            .in0(N__48344),
            .in1(N__34343),
            .in2(N__46189),
            .in3(N__34395),
            .lcout(\ALU.dZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(N__43345),
            .sr(_gnd_net_));
    defparam \ALU.d_11_LC_10_9_1 .C_ON=1'b0;
    defparam \ALU.d_11_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \ALU.d_11_LC_10_9_1 .LUT_INIT=16'b0101110101010001;
    LogicCell40 \ALU.d_11_LC_10_9_1  (
            .in0(N__34250),
            .in1(N__46163),
            .in2(N__48575),
            .in3(N__34160),
            .lcout(\ALU.dZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(N__43345),
            .sr(_gnd_net_));
    defparam \ALU.d_12_LC_10_9_2 .C_ON=1'b0;
    defparam \ALU.d_12_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \ALU.d_12_LC_10_9_2 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.d_12_LC_10_9_2  (
            .in0(N__48345),
            .in1(N__34087),
            .in2(N__46190),
            .in3(N__34010),
            .lcout(\ALU.dZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(N__43345),
            .sr(_gnd_net_));
    defparam \ALU.d_14_LC_10_9_3 .C_ON=1'b0;
    defparam \ALU.d_14_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \ALU.d_14_LC_10_9_3 .LUT_INIT=16'b0101110101010001;
    LogicCell40 \ALU.d_14_LC_10_9_3  (
            .in0(N__33812),
            .in1(N__46165),
            .in2(N__48576),
            .in3(N__33740),
            .lcout(\ALU.dZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(N__43345),
            .sr(_gnd_net_));
    defparam \ALU.d_15_LC_10_9_4 .C_ON=1'b0;
    defparam \ALU.d_15_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \ALU.d_15_LC_10_9_4 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \ALU.d_15_LC_10_9_4  (
            .in0(N__48346),
            .in1(N__33659),
            .in2(N__46191),
            .in3(N__33591),
            .lcout(\ALU.dZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(N__43345),
            .sr(_gnd_net_));
    defparam \ALU.d_13_LC_10_9_5 .C_ON=1'b0;
    defparam \ALU.d_13_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \ALU.d_13_LC_10_9_5 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.d_13_LC_10_9_5  (
            .in0(N__48412),
            .in1(N__46164),
            .in2(N__33941),
            .in3(N__33864),
            .lcout(\ALU.dZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(N__43345),
            .sr(_gnd_net_));
    defparam \ALU.d_9_LC_10_9_6 .C_ON=1'b0;
    defparam \ALU.d_9_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \ALU.d_9_LC_10_9_6 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.d_9_LC_10_9_6  (
            .in0(N__48347),
            .in1(N__36260),
            .in2(N__46192),
            .in3(N__36178),
            .lcout(\ALU.dZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(N__43345),
            .sr(_gnd_net_));
    defparam \ALU.e_10_LC_10_10_0 .C_ON=1'b0;
    defparam \ALU.e_10_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.e_10_LC_10_10_0 .LUT_INIT=16'b0101010111000101;
    LogicCell40 \ALU.e_10_LC_10_10_0  (
            .in0(N__34344),
            .in1(N__34384),
            .in2(N__46147),
            .in3(N__48560),
            .lcout(\ALU.eZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(N__32457),
            .sr(_gnd_net_));
    defparam \ALU.e_11_LC_10_10_1 .C_ON=1'b0;
    defparam \ALU.e_11_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \ALU.e_11_LC_10_10_1 .LUT_INIT=16'b0101110101010001;
    LogicCell40 \ALU.e_11_LC_10_10_1  (
            .in0(N__34247),
            .in1(N__46060),
            .in2(N__48634),
            .in3(N__34147),
            .lcout(\ALU.eZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(N__32457),
            .sr(_gnd_net_));
    defparam \ALU.e_12_LC_10_10_2 .C_ON=1'b0;
    defparam \ALU.e_12_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.e_12_LC_10_10_2 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.e_12_LC_10_10_2  (
            .in0(N__48572),
            .in1(N__34090),
            .in2(N__46148),
            .in3(N__34000),
            .lcout(\ALU.eZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(N__32457),
            .sr(_gnd_net_));
    defparam \ALU.e_13_LC_10_10_3 .C_ON=1'b0;
    defparam \ALU.e_13_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \ALU.e_13_LC_10_10_3 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.e_13_LC_10_10_3  (
            .in0(N__48555),
            .in1(N__33934),
            .in2(N__46150),
            .in3(N__33853),
            .lcout(\ALU.eZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(N__32457),
            .sr(_gnd_net_));
    defparam \ALU.e_14_LC_10_10_4 .C_ON=1'b0;
    defparam \ALU.e_14_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \ALU.e_14_LC_10_10_4 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.e_14_LC_10_10_4  (
            .in0(N__48573),
            .in1(N__33814),
            .in2(N__46149),
            .in3(N__33727),
            .lcout(\ALU.eZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(N__32457),
            .sr(_gnd_net_));
    defparam \ALU.e_15_LC_10_10_5 .C_ON=1'b0;
    defparam \ALU.e_15_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \ALU.e_15_LC_10_10_5 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \ALU.e_15_LC_10_10_5  (
            .in0(N__48556),
            .in1(N__33660),
            .in2(N__46151),
            .in3(N__33589),
            .lcout(\ALU.eZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(N__32457),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIPER7_5_LC_10_10_6 .C_ON=1'b0;
    defparam \ALU.d_RNIPER7_5_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIPER7_5_LC_10_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIPER7_5_LC_10_10_6  (
            .in0(N__45063),
            .in1(N__31396),
            .in2(_gnd_net_),
            .in3(N__43396),
            .lcout(\ALU.d_RNIPER7Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_10_LC_10_11_0 .C_ON=1'b0;
    defparam \ALU.b_10_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.b_10_LC_10_11_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.b_10_LC_10_11_0  (
            .in0(N__48076),
            .in1(N__34345),
            .in2(N__46193),
            .in3(N__34394),
            .lcout(\ALU.bZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47651),
            .ce(N__47402),
            .sr(_gnd_net_));
    defparam \ALU.b_15_LC_10_11_1 .C_ON=1'b0;
    defparam \ALU.b_15_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.b_15_LC_10_11_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \ALU.b_15_LC_10_11_1  (
            .in0(N__48092),
            .in1(N__33661),
            .in2(N__46122),
            .in3(N__33590),
            .lcout(\ALU.bZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47651),
            .ce(N__47402),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_12_c_RNIG3PMU_LC_10_11_2 .C_ON=1'b0;
    defparam \ALU.un2_addsub_cry_12_c_RNIG3PMU_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_12_c_RNIG3PMU_LC_10_11_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ALU.un2_addsub_cry_12_c_RNIG3PMU_LC_10_11_2  (
            .in0(N__42518),
            .in1(N__40649),
            .in2(_gnd_net_),
            .in3(N__28700),
            .lcout(),
            .ltout(un2_addsub_cry_12_c_RNIG3PMU_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_RNI2J9SL3_0_LC_10_11_3 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_RNI2J9SL3_0_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_RNI2J9SL3_0_LC_10_11_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \CONTROL.aluOperation_RNI2J9SL3_0_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__48075),
            .in2(N__28688),
            .in3(N__28685),
            .lcout(aluOperation_RNI2J9SL3_0),
            .ltout(aluOperation_RNI2J9SL3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_13_LC_10_11_4 .C_ON=1'b0;
    defparam \ALU.b_13_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \ALU.b_13_LC_10_11_4 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.b_13_LC_10_11_4  (
            .in0(N__48077),
            .in1(N__46046),
            .in2(N__28670),
            .in3(N__33863),
            .lcout(\ALU.bZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47651),
            .ce(N__47402),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIFMN04_2_LC_10_11_5 .C_ON=1'b0;
    defparam \ALU.d_RNIIFMN04_2_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIFMN04_2_LC_10_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIIFMN04_2_LC_10_11_5  (
            .in0(N__46045),
            .in1(N__28667),
            .in2(_gnd_net_),
            .in3(N__28655),
            .lcout(\ALU.d_RNIIFMN04Z0Z_2 ),
            .ltout(\ALU.d_RNIIFMN04Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_2_LC_10_11_6 .C_ON=1'b0;
    defparam \ALU.b_2_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \ALU.b_2_LC_10_11_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \ALU.b_2_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(N__42151),
            .in2(N__28640),
            .in3(N__48093),
            .lcout(\ALU.bZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47651),
            .ce(N__47402),
            .sr(_gnd_net_));
    defparam \ALU.e_0_LC_10_12_0 .C_ON=1'b0;
    defparam \ALU.e_0_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.e_0_LC_10_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_0_LC_10_12_0  (
            .in0(N__48430),
            .in1(N__42321),
            .in2(_gnd_net_),
            .in3(N__42252),
            .lcout(\ALU.eZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47657),
            .ce(N__32468),
            .sr(_gnd_net_));
    defparam \ALU.e_2_LC_10_12_1 .C_ON=1'b0;
    defparam \ALU.e_2_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.e_2_LC_10_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_2_LC_10_12_1  (
            .in0(N__48567),
            .in1(N__42162),
            .in2(_gnd_net_),
            .in3(N__42078),
            .lcout(\ALU.eZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47657),
            .ce(N__32468),
            .sr(_gnd_net_));
    defparam \ALU.e_3_LC_10_12_2 .C_ON=1'b0;
    defparam \ALU.e_3_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.e_3_LC_10_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_3_LC_10_12_2  (
            .in0(N__48431),
            .in1(N__49468),
            .in2(_gnd_net_),
            .in3(N__49387),
            .lcout(\ALU.eZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47657),
            .ce(N__32468),
            .sr(_gnd_net_));
    defparam \ALU.e_6_LC_10_12_3 .C_ON=1'b0;
    defparam \ALU.e_6_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.e_6_LC_10_12_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.e_6_LC_10_12_3  (
            .in0(N__48932),
            .in1(N__48432),
            .in2(_gnd_net_),
            .in3(N__48881),
            .lcout(\ALU.eZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47657),
            .ce(N__32468),
            .sr(_gnd_net_));
    defparam \ALU.e_7_LC_10_12_4 .C_ON=1'b0;
    defparam \ALU.e_7_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.e_7_LC_10_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.e_7_LC_10_12_4  (
            .in0(N__48713),
            .in1(N__48569),
            .in2(_gnd_net_),
            .in3(N__48777),
            .lcout(\ALU.eZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47657),
            .ce(N__32468),
            .sr(_gnd_net_));
    defparam \ALU.e_8_LC_10_12_5 .C_ON=1'b0;
    defparam \ALU.e_8_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.e_8_LC_10_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_8_LC_10_12_5  (
            .in0(N__48568),
            .in1(N__47886),
            .in2(_gnd_net_),
            .in3(N__47794),
            .lcout(\ALU.eZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47657),
            .ce(N__32468),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_fast_1_LC_10_13_0 .C_ON=1'b0;
    defparam \CONTROL.operand2_fast_1_LC_10_13_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_fast_1_LC_10_13_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \CONTROL.operand2_fast_1_LC_10_13_0  (
            .in0(N__34764),
            .in1(N__31014),
            .in2(N__34709),
            .in3(N__34566),
            .lcout(aluOperand2_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47665),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_1_rep1_LC_10_13_1 .C_ON=1'b0;
    defparam \CONTROL.operand2_1_rep1_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_1_rep1_LC_10_13_1 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \CONTROL.operand2_1_rep1_LC_10_13_1  (
            .in0(N__34567),
            .in1(N__34765),
            .in2(N__34708),
            .in3(N__34994),
            .lcout(aluOperand2_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47665),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_fast_2_LC_10_13_2 .C_ON=1'b0;
    defparam \CONTROL.operand2_fast_2_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_fast_2_LC_10_13_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \CONTROL.operand2_fast_2_LC_10_13_2  (
            .in0(N__34867),
            .in1(N__32224),
            .in2(N__34787),
            .in3(N__34685),
            .lcout(aluOperand2_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47665),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIRMVJ_2_LC_10_13_3 .C_ON=1'b0;
    defparam \ALU.e_RNIRMVJ_2_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIRMVJ_2_LC_10_13_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \ALU.e_RNIRMVJ_2_LC_10_13_3  (
            .in0(N__28780),
            .in1(N__28759),
            .in2(N__34868),
            .in3(_gnd_net_),
            .lcout(\ALU.e_RNIRMVJZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIV2CO_2_LC_10_13_4 .C_ON=1'b0;
    defparam \ALU.g_RNIV2CO_2_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIV2CO_2_LC_10_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.g_RNIV2CO_2_LC_10_13_4  (
            .in0(N__29089),
            .in1(N__34855),
            .in2(_gnd_net_),
            .in3(N__31894),
            .lcout(),
            .ltout(\ALU.g_RNIV2COZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIPKSL1_2_LC_10_13_5 .C_ON=1'b0;
    defparam \ALU.e_RNIPKSL1_2_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIPKSL1_2_LC_10_13_5 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \ALU.e_RNIPKSL1_2_LC_10_13_5  (
            .in0(N__31013),
            .in1(N__31577),
            .in2(N__28742),
            .in3(N__28739),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIAUJU2_2_LC_10_13_6 .C_ON=1'b0;
    defparam \ALU.d_RNIAUJU2_2_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIAUJU2_2_LC_10_13_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIAUJU2_2_LC_10_13_6  (
            .in0(N__33089),
            .in1(N__28811),
            .in2(N__28733),
            .in3(N__31949),
            .lcout(\ALU.operand2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNINIVJ_0_LC_10_13_7 .C_ON=1'b0;
    defparam \ALU.e_RNINIVJ_0_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNINIVJ_0_LC_10_13_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_RNINIVJ_0_LC_10_13_7  (
            .in0(N__34854),
            .in1(N__28948),
            .in2(_gnd_net_),
            .in3(N__28926),
            .lcout(\ALU.e_RNINIVJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIM8LL_5_LC_10_14_0 .C_ON=1'b0;
    defparam \ALU.g_RNIM8LL_5_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIM8LL_5_LC_10_14_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_RNIM8LL_5_LC_10_14_0  (
            .in0(N__32025),
            .in1(N__31825),
            .in2(_gnd_net_),
            .in3(N__29026),
            .lcout(\ALU.g_RNIM8LLZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNI1TVJ_5_LC_10_14_1 .C_ON=1'b0;
    defparam \ALU.e_RNI1TVJ_5_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNI1TVJ_5_LC_10_14_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.e_RNI1TVJ_5_LC_10_14_1  (
            .in0(N__34863),
            .in1(N__44628),
            .in2(_gnd_net_),
            .in3(N__28861),
            .lcout(),
            .ltout(\ALU.e_RNI1TVJZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIOJPU1_5_LC_10_14_2 .C_ON=1'b0;
    defparam \ALU.e_RNIOJPU1_5_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIOJPU1_5_LC_10_14_2 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \ALU.e_RNIOJPU1_5_LC_10_14_2  (
            .in0(N__28892),
            .in1(N__34993),
            .in2(N__28886),
            .in3(N__31263),
            .lcout(\ALU.operand2_7_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_5_LC_10_14_3 .C_ON=1'b0;
    defparam \ALU.e_5_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.e_5_LC_10_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.e_5_LC_10_14_3  (
            .in0(N__48426),
            .in1(N__49130),
            .in2(_gnd_net_),
            .in3(N__49045),
            .lcout(\ALU.eZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47672),
            .ce(N__32467),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIRUBO_0_LC_10_14_4 .C_ON=1'b0;
    defparam \ALU.g_RNIRUBO_0_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIRUBO_0_LC_10_14_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.g_RNIRUBO_0_LC_10_14_4  (
            .in0(N__29134),
            .in1(N__34862),
            .in2(_gnd_net_),
            .in3(N__31933),
            .lcout(\ALU.g_RNIRUBOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIG6R7_1_LC_10_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNIG6R7_1_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIG6R7_1_LC_10_14_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNIG6R7_1_LC_10_14_5  (
            .in0(N__31441),
            .in1(N__32027),
            .in2(_gnd_net_),
            .in3(N__36553),
            .lcout(\ALU.d_RNIG6R7Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI45J9_1_LC_10_14_6 .C_ON=1'b0;
    defparam \ALU.d_RNI45J9_1_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI45J9_1_LC_10_14_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ALU.d_RNI45J9_1_LC_10_14_6  (
            .in0(N__36554),
            .in1(_gnd_net_),
            .in2(N__35586),
            .in3(N__31442),
            .lcout(\ALU.d_RNI45J9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNII8R7_2_LC_10_14_7 .C_ON=1'b0;
    defparam \ALU.d_RNII8R7_2_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNII8R7_2_LC_10_14_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_RNII8R7_2_LC_10_14_7  (
            .in0(N__31423),
            .in1(N__32026),
            .in2(_gnd_net_),
            .in3(N__42034),
            .lcout(\ALU.d_RNII8R7Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_0_LC_10_15_0 .C_ON=1'b0;
    defparam \ALU.c_0_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \ALU.c_0_LC_10_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_0_LC_10_15_0  (
            .in0(N__48631),
            .in1(N__42322),
            .in2(_gnd_net_),
            .in3(N__42254),
            .lcout(\ALU.cZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.c_1_LC_10_15_1 .C_ON=1'b0;
    defparam \ALU.c_1_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \ALU.c_1_LC_10_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_1_LC_10_15_1  (
            .in0(N__48421),
            .in1(N__41000),
            .in2(_gnd_net_),
            .in3(N__36613),
            .lcout(\ALU.cZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.c_2_LC_10_15_2 .C_ON=1'b0;
    defparam \ALU.c_2_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \ALU.c_2_LC_10_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_2_LC_10_15_2  (
            .in0(N__48632),
            .in1(N__42164),
            .in2(_gnd_net_),
            .in3(N__42092),
            .lcout(\ALU.cZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.c_3_LC_10_15_3 .C_ON=1'b0;
    defparam \ALU.c_3_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \ALU.c_3_LC_10_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_3_LC_10_15_3  (
            .in0(N__48422),
            .in1(N__49467),
            .in2(_gnd_net_),
            .in3(N__49388),
            .lcout(\ALU.cZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.c_4_LC_10_15_4 .C_ON=1'b0;
    defparam \ALU.c_4_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \ALU.c_4_LC_10_15_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.c_4_LC_10_15_4  (
            .in0(N__49218),
            .in1(N__48424),
            .in2(_gnd_net_),
            .in3(N__49285),
            .lcout(\ALU.cZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.c_5_LC_10_15_5 .C_ON=1'b0;
    defparam \ALU.c_5_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \ALU.c_5_LC_10_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_5_LC_10_15_5  (
            .in0(N__48423),
            .in1(N__49112),
            .in2(_gnd_net_),
            .in3(N__49047),
            .lcout(\ALU.cZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.c_6_LC_10_15_6 .C_ON=1'b0;
    defparam \ALU.c_6_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \ALU.c_6_LC_10_15_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.c_6_LC_10_15_6  (
            .in0(N__48943),
            .in1(N__48425),
            .in2(_gnd_net_),
            .in3(N__48892),
            .lcout(\ALU.cZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.c_7_LC_10_15_7 .C_ON=1'b0;
    defparam \ALU.c_7_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \ALU.c_7_LC_10_15_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.c_7_LC_10_15_7  (
            .in0(N__48715),
            .in1(N__48633),
            .in2(_gnd_net_),
            .in3(N__48749),
            .lcout(\ALU.cZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(N__31502),
            .sr(_gnd_net_));
    defparam \ALU.d_4_LC_10_16_7 .C_ON=1'b0;
    defparam \ALU.d_4_LC_10_16_7 .SEQ_MODE=4'b1000;
    defparam \ALU.d_4_LC_10_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_4_LC_10_16_7  (
            .in0(N__48629),
            .in1(N__49287),
            .in2(_gnd_net_),
            .in3(N__49219),
            .lcout(\ALU.dZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47682),
            .ce(N__43346),
            .sr(_gnd_net_));
    defparam \ALU.g_6_LC_10_17_5 .C_ON=1'b0;
    defparam \ALU.g_6_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \ALU.g_6_LC_10_17_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_6_LC_10_17_5  (
            .in0(N__48630),
            .in1(N__48893),
            .in2(_gnd_net_),
            .in3(N__48947),
            .lcout(\ALU.gZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47685),
            .ce(N__36104),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_21_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_21_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_21_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.gap_2_LC_11_1_2 .C_ON=1'b0;
    defparam \FTDI.gap_2_LC_11_1_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.gap_2_LC_11_1_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \FTDI.gap_2_LC_11_1_2  (
            .in0(N__29194),
            .in1(_gnd_net_),
            .in2(N__29219),
            .in3(N__29168),
            .lcout(\FTDI.gapZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.gap_1_LC_11_1_5 .C_ON=1'b0;
    defparam \FTDI.gap_1_LC_11_1_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.gap_1_LC_11_1_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \FTDI.gap_1_LC_11_1_5  (
            .in0(N__29167),
            .in1(N__29215),
            .in2(_gnd_net_),
            .in3(N__29193),
            .lcout(\FTDI.gapZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.gap_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNICVLM_0_LC_11_2_0 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNICVLM_0_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNICVLM_0_LC_11_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FTDI.TXstate_RNICVLM_0_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__30377),
            .in2(_gnd_net_),
            .in3(N__29518),
            .lcout(\FTDI.N_169_0 ),
            .ltout(\FTDI.N_169_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_0_LC_11_2_1 .C_ON=1'b0;
    defparam \FTDI.TXstate_0_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_0_LC_11_2_1 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \FTDI.TXstate_0_LC_11_2_1  (
            .in0(N__32322),
            .in1(N__29159),
            .in2(N__29153),
            .in3(N__29494),
            .lcout(\FTDI.TXstateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_1_LC_11_2_2 .C_ON=1'b0;
    defparam \FTDI.TXstate_1_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_1_LC_11_2_2 .LUT_INIT=16'b1010101001001000;
    LogicCell40 \FTDI.TXstate_1_LC_11_2_2  (
            .in0(N__29495),
            .in1(N__44744),
            .in2(N__29150),
            .in3(N__29597),
            .lcout(\FTDI.TXstateZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_2_LC_11_2_4 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_2_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_2_LC_11_2_4 .LUT_INIT=16'b1101011100000111;
    LogicCell40 \FTDI.TXstate_RNO_0_2_LC_11_2_4  (
            .in0(N__44719),
            .in1(N__29467),
            .in2(N__32327),
            .in3(N__30379),
            .lcout(),
            .ltout(\FTDI.TXstate_cnst_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_2_LC_11_2_5 .C_ON=1'b0;
    defparam \FTDI.TXstate_2_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_2_LC_11_2_5 .LUT_INIT=16'b1100111100001111;
    LogicCell40 \FTDI.TXstate_2_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(N__30410),
            .in2(N__29141),
            .in3(N__30341),
            .lcout(\FTDI.un3_TX_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXstate_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_1_1_LC_11_2_6 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_1_1_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_1_1_LC_11_2_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \FTDI.TXstate_RNO_1_1_LC_11_2_6  (
            .in0(_gnd_net_),
            .in1(N__32321),
            .in2(_gnd_net_),
            .in3(N__29517),
            .lcout(),
            .ltout(\FTDI.N_217_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_1_LC_11_2_7 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_1_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_1_LC_11_2_7 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \FTDI.TXstate_RNO_0_1_LC_11_2_7  (
            .in0(N__30378),
            .in1(N__44718),
            .in2(N__29600),
            .in3(N__29493),
            .lcout(\FTDI.N_216_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNINQ101_0_LC_11_3_0 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNINQ101_0_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNINQ101_0_LC_11_3_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \FTDI.TXstate_RNINQ101_0_LC_11_3_0  (
            .in0(N__30384),
            .in1(N__29519),
            .in2(_gnd_net_),
            .in3(N__29490),
            .lcout(\FTDI.N_170_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNIEFF51_0_LC_11_3_1 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNIEFF51_0_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNIEFF51_0_LC_11_3_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \FTDI.TXstate_RNIEFF51_0_LC_11_3_1  (
            .in0(N__29520),
            .in1(N__29492),
            .in2(N__44748),
            .in3(N__32319),
            .lcout(\FTDI.TXready ),
            .ltout(\FTDI.TXready_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_1_LC_11_3_2 .C_ON=1'b0;
    defparam \FTDI.baudAcc_1_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \FTDI.baudAcc_1_LC_11_3_2 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \FTDI.baudAcc_1_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__29563),
            .in2(N__29591),
            .in3(N__29588),
            .lcout(\FTDI.baudAccZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNID2HKH1_5_LC_11_3_3 .C_ON=1'b0;
    defparam \ALU.d_RNID2HKH1_5_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNID2HKH1_5_LC_11_3_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNID2HKH1_5_LC_11_3_3  (
            .in0(N__43179),
            .in1(N__29552),
            .in2(_gnd_net_),
            .in3(N__29534),
            .lcout(\ALU.a_15_m3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_RNO_0_3_LC_11_3_6 .C_ON=1'b0;
    defparam \FTDI.TXstate_RNO_0_3_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \FTDI.TXstate_RNO_0_3_LC_11_3_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \FTDI.TXstate_RNO_0_3_LC_11_3_6  (
            .in0(N__30385),
            .in1(N__29521),
            .in2(_gnd_net_),
            .in3(N__29491),
            .lcout(),
            .ltout(\FTDI.TXstate_e_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.TXstate_3_LC_11_3_7 .C_ON=1'b0;
    defparam \FTDI.TXstate_3_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXstate_3_LC_11_3_7 .LUT_INIT=16'b1111001010101010;
    LogicCell40 \FTDI.TXstate_3_LC_11_3_7  (
            .in0(N__44717),
            .in1(N__29468),
            .in2(N__29456),
            .in3(N__32320),
            .lcout(\FTDI.TXstateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.baudAcc_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI1OCN4_15_LC_11_4_0 .C_ON=1'b0;
    defparam \ALU.c_RNI1OCN4_15_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI1OCN4_15_LC_11_4_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \ALU.c_RNI1OCN4_15_LC_11_4_0  (
            .in0(N__29453),
            .in1(N__32666),
            .in2(_gnd_net_),
            .in3(N__29437),
            .lcout(),
            .ltout(\ALU.c_RNI1OCN4Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI68L5A_15_LC_11_4_1 .C_ON=1'b0;
    defparam \ALU.c_RNI68L5A_15_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI68L5A_15_LC_11_4_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.c_RNI68L5A_15_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__43172),
            .in2(N__30560),
            .in3(N__30443),
            .lcout(\ALU.a_15_m3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIKUKV3_15_LC_11_4_2 .C_ON=1'b0;
    defparam \ALU.c_RNIKUKV3_15_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIKUKV3_15_LC_11_4_2 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \ALU.c_RNIKUKV3_15_LC_11_4_2  (
            .in0(N__30557),
            .in1(N__30535),
            .in2(N__43747),
            .in3(N__35223),
            .lcout(\ALU.N_621_1 ),
            .ltout(\ALU.N_621_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI8597C_15_LC_11_4_3 .C_ON=1'b0;
    defparam \ALU.c_RNI8597C_15_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI8597C_15_LC_11_4_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNI8597C_15_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__39151),
            .in2(N__30506),
            .in3(N__30502),
            .lcout(\ALU.N_578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI4JFV4_0_15_LC_11_4_5 .C_ON=1'b0;
    defparam \ALU.c_RNI4JFV4_0_15_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI4JFV4_0_15_LC_11_4_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ALU.c_RNI4JFV4_0_15_LC_11_4_5  (
            .in0(N__38713),
            .in1(N__39152),
            .in2(N__44525),
            .in3(N__30471),
            .lcout(\ALU.c_RNI4JFV4_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI36KJ21_9_LC_11_4_6 .C_ON=1'b0;
    defparam \ALU.d_RNI36KJ21_9_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI36KJ21_9_LC_11_4_6 .LUT_INIT=16'b0101001100000011;
    LogicCell40 \ALU.d_RNI36KJ21_9_LC_11_4_6  (
            .in0(N__44499),
            .in1(N__30437),
            .in2(N__43184),
            .in3(N__31751),
            .lcout(\ALU.d_RNI36KJ21Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.baudAcc_RNINKH42_2_LC_11_5_0 .C_ON=1'b0;
    defparam \FTDI.baudAcc_RNINKH42_2_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.baudAcc_RNINKH42_2_LC_11_5_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \FTDI.baudAcc_RNINKH42_2_LC_11_5_0  (
            .in0(N__30417),
            .in1(N__30336),
            .in2(N__44768),
            .in3(N__30386),
            .lcout(\FTDI.un1_TXstate_0_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TXstart_LC_11_5_1.C_ON=1'b0;
    defparam TXstart_LC_11_5_1.SEQ_MODE=4'b1000;
    defparam TXstart_LC_11_5_1.LUT_INIT=16'b0010111010101000;
    LogicCell40 TXstart_LC_11_5_1 (
            .in0(N__30337),
            .in1(N__30808),
            .in2(N__30322),
            .in3(N__41413),
            .lcout(TXstartZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47610),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m326dup_LC_11_5_2 .C_ON=1'b0;
    defparam \ALU.m326dup_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \ALU.m326dup_LC_11_5_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ALU.m326dup_LC_11_5_2  (
            .in0(N__30807),
            .in1(N__41409),
            .in2(_gnd_net_),
            .in3(N__30315),
            .lcout(m326dup),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g0_7_LC_11_5_4 .C_ON=1'b0;
    defparam \ALU.g0_7_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \ALU.g0_7_LC_11_5_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ALU.g0_7_LC_11_5_4  (
            .in0(N__30239),
            .in1(N__30218),
            .in2(N__30025),
            .in3(N__29754),
            .lcout(\ALU.N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testState_RNIB7C_2_LC_11_5_6.C_ON=1'b0;
    defparam testState_RNIB7C_2_LC_11_5_6.SEQ_MODE=4'b0000;
    defparam testState_RNIB7C_2_LC_11_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 testState_RNIB7C_2_LC_11_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30806),
            .lcout(testState_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIJTBO_14_LC_11_5_7 .C_ON=1'b0;
    defparam \ALU.a_RNIJTBO_14_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIJTBO_14_LC_11_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.a_RNIJTBO_14_LC_11_5_7  (
            .in0(N__30721),
            .in1(N__31378),
            .in2(_gnd_net_),
            .in3(N__45128),
            .lcout(\ALU.a_RNIJTBOZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_13_c_RNI2LH1U_LC_11_6_0 .C_ON=1'b0;
    defparam \ALU.un2_addsub_cry_13_c_RNI2LH1U_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_13_c_RNI2LH1U_LC_11_6_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ALU.un2_addsub_cry_13_c_RNI2LH1U_LC_11_6_0  (
            .in0(N__42458),
            .in1(N__40538),
            .in2(_gnd_net_),
            .in3(N__30704),
            .lcout(),
            .ltout(un2_addsub_cry_13_c_RNI2LH1U_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_RNIR872K3_0_LC_11_6_1 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_RNIR872K3_0_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_RNIR872K3_0_LC_11_6_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \CONTROL.aluOperation_RNIR872K3_0_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__48271),
            .in2(N__30686),
            .in3(N__30683),
            .lcout(aluOperation_RNIR872K3_0),
            .ltout(aluOperation_RNIR872K3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_14_LC_11_6_2 .C_ON=1'b0;
    defparam \ALU.h_14_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \ALU.h_14_LC_11_6_2 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.h_14_LC_11_6_2  (
            .in0(N__48272),
            .in1(N__45930),
            .in2(N__30668),
            .in3(N__33757),
            .lcout(\ALU.hZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47614),
            .ce(N__45567),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIEH3U1_14_LC_11_6_3 .C_ON=1'b0;
    defparam \ALU.c_RNIEH3U1_14_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIEH3U1_14_LC_11_6_3 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \ALU.c_RNIEH3U1_14_LC_11_6_3  (
            .in0(N__34495),
            .in1(N__31532),
            .in2(N__30665),
            .in3(N__33065),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIGLRP4_14_LC_11_6_4 .C_ON=1'b0;
    defparam \ALU.d_RNIGLRP4_14_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIGLRP4_14_LC_11_6_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIGLRP4_14_LC_11_6_4  (
            .in0(N__32971),
            .in1(N__30566),
            .in2(N__30656),
            .in3(N__30653),
            .lcout(\ALU.operand2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIQ9LU_14_LC_11_6_5 .C_ON=1'b0;
    defparam \ALU.d_RNIQ9LU_14_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIQ9LU_14_LC_11_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIQ9LU_14_LC_11_6_5  (
            .in0(N__30610),
            .in1(N__30589),
            .in2(_gnd_net_),
            .in3(N__45322),
            .lcout(\ALU.d_RNIQ9LUZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_8_LC_11_7_0 .C_ON=1'b0;
    defparam \ALU.a_8_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \ALU.a_8_LC_11_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_8_LC_11_7_0  (
            .in0(N__48267),
            .in1(N__47827),
            .in2(_gnd_net_),
            .in3(N__47777),
            .lcout(\ALU.aZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47620),
            .ce(N__44871),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_7_c_RNIQIKVO_LC_11_7_1 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_7_c_RNIQIKVO_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_7_c_RNIQIKVO_LC_11_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.un9_addsub_cry_7_c_RNIQIKVO_LC_11_7_1  (
            .in0(N__42463),
            .in1(N__39875),
            .in2(_gnd_net_),
            .in3(N__31082),
            .lcout(\ALU.un9_addsub_cry_7_c_RNIQIKVOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIOG1M_8_LC_11_7_2 .C_ON=1'b0;
    defparam \ALU.e_RNIOG1M_8_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIOG1M_8_LC_11_7_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.e_RNIOG1M_8_LC_11_7_2  (
            .in0(N__31060),
            .in1(N__31042),
            .in2(N__30973),
            .in3(N__32073),
            .lcout(),
            .ltout(\ALU.operand2_3_ns_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIJQCH1_8_LC_11_7_3 .C_ON=1'b0;
    defparam \ALU.g_RNIJQCH1_8_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIJQCH1_8_LC_11_7_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.g_RNIJQCH1_8_LC_11_7_3  (
            .in0(N__30937),
            .in1(N__30901),
            .in2(N__30878),
            .in3(N__35030),
            .lcout(\ALU.N_819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m715_LC_11_7_4 .C_ON=1'b0;
    defparam \ALU.m715_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.m715_LC_11_7_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ALU.m715_LC_11_7_4  (
            .in0(N__48265),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43728),
            .lcout(\ALU.addsub_0_sqmuxa ),
            .ltout(\ALU.addsub_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_8_c_RNIKTS9S_LC_11_7_5 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_8_c_RNIKTS9S_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_8_c_RNIKTS9S_LC_11_7_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ALU.un9_addsub_cry_8_c_RNIKTS9S_LC_11_7_5  (
            .in0(N__39623),
            .in1(_gnd_net_),
            .in2(N__30860),
            .in3(N__30857),
            .lcout(),
            .ltout(\ALU.un9_addsub_cry_8_c_RNIKTS9SZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_8_c_RNIPHQ7I3_LC_11_7_6 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_8_c_RNIPHQ7I3_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_8_c_RNIPHQ7I3_LC_11_7_6 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \ALU.un9_addsub_cry_8_c_RNIPHQ7I3_LC_11_7_6  (
            .in0(N__48266),
            .in1(_gnd_net_),
            .in2(N__30845),
            .in3(N__30842),
            .lcout(\ALU.a_15_ns_1_9 ),
            .ltout(\ALU.a_15_ns_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_9_LC_11_7_7 .C_ON=1'b0;
    defparam \ALU.a_9_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \ALU.a_9_LC_11_7_7 .LUT_INIT=16'b0010111100001101;
    LogicCell40 \ALU.a_9_LC_11_7_7  (
            .in0(N__45990),
            .in1(N__48268),
            .in2(N__30833),
            .in3(N__36203),
            .lcout(\ALU.aZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47620),
            .ce(N__44871),
            .sr(_gnd_net_));
    defparam \ALU.a_RNICNBO_11_LC_11_8_0 .C_ON=1'b0;
    defparam \ALU.a_RNICNBO_11_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNICNBO_11_LC_11_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.a_RNICNBO_11_LC_11_8_0  (
            .in0(N__32067),
            .in1(N__32482),
            .in2(_gnd_net_),
            .in3(N__30826),
            .lcout(),
            .ltout(\ALU.a_RNICNBOZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNITCKM1_11_LC_11_8_1 .C_ON=1'b0;
    defparam \ALU.c_RNITCKM1_11_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNITCKM1_11_LC_11_8_1 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \ALU.c_RNITCKM1_11_LC_11_8_1  (
            .in0(N__35031),
            .in1(N__31249),
            .in2(N__31193),
            .in3(N__31118),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJ4CI4_11_LC_11_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNIJ4CI4_11_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJ4CI4_11_LC_11_8_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIJ4CI4_11_LC_11_8_2  (
            .in0(N__32902),
            .in1(N__31142),
            .in2(N__31190),
            .in3(N__31187),
            .lcout(\ALU.operand2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIK3LU_11_LC_11_8_3 .C_ON=1'b0;
    defparam \ALU.d_RNIK3LU_11_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIK3LU_11_LC_11_8_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIK3LU_11_LC_11_8_3  (
            .in0(N__45275),
            .in1(N__31129),
            .in2(_gnd_net_),
            .in3(N__31153),
            .lcout(\ALU.d_RNIK3LUZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_11_LC_11_8_4 .C_ON=1'b0;
    defparam \ALU.h_11_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \ALU.h_11_LC_11_8_4 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.h_11_LC_11_8_4  (
            .in0(N__48348),
            .in1(N__34248),
            .in2(N__46117),
            .in3(N__34180),
            .lcout(\ALU.hZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47627),
            .ce(N__45538),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIG749_11_LC_11_8_5 .C_ON=1'b0;
    defparam \ALU.c_RNIG749_11_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIG749_11_LC_11_8_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.c_RNIG749_11_LC_11_8_5  (
            .in0(N__34105),
            .in1(N__32066),
            .in2(_gnd_net_),
            .in3(N__31300),
            .lcout(\ALU.c_RNIG749Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNILB49_13_LC_11_9_0 .C_ON=1'b0;
    defparam \ALU.c_RNILB49_13_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNILB49_13_LC_11_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ALU.c_RNILB49_13_LC_11_9_0  (
            .in0(N__35809),
            .in1(N__35794),
            .in2(_gnd_net_),
            .in3(N__45076),
            .lcout(\ALU.c_RNILB49Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNIHRBO_13_LC_11_9_1 .C_ON=1'b0;
    defparam \ALU.a_RNIHRBO_13_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNIHRBO_13_LC_11_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_RNIHRBO_13_LC_11_9_1  (
            .in0(N__45077),
            .in1(N__36031),
            .in2(_gnd_net_),
            .in3(N__36020),
            .lcout(),
            .ltout(\ALU.a_RNIHRBOZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIAD3U1_13_LC_11_9_2 .C_ON=1'b0;
    defparam \ALU.c_RNIAD3U1_13_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIAD3U1_13_LC_11_9_2 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.c_RNIAD3U1_13_LC_11_9_2  (
            .in0(N__33063),
            .in1(N__34468),
            .in2(N__31112),
            .in3(N__31109),
            .lcout(\ALU.operand2_7_ns_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_2_rep2_LC_11_9_3 .C_ON=1'b0;
    defparam \CONTROL.operand2_2_rep2_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_2_rep2_LC_11_9_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \CONTROL.operand2_2_rep2_LC_11_9_3  (
            .in0(N__45080),
            .in1(N__32214),
            .in2(N__34720),
            .in3(N__34797),
            .lcout(aluOperand2_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47634),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIPF49_15_LC_11_9_4 .C_ON=1'b0;
    defparam \ALU.c_RNIPF49_15_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIPF49_15_LC_11_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.c_RNIPF49_15_LC_11_9_4  (
            .in0(N__31522),
            .in1(N__45078),
            .in2(_gnd_net_),
            .in3(N__33535),
            .lcout(\ALU.c_RNIPF49Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_RNILVBO_15_LC_11_9_5 .C_ON=1'b0;
    defparam \ALU.a_RNILVBO_15_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNILVBO_15_LC_11_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_RNILVBO_15_LC_11_9_5  (
            .in0(N__45079),
            .in1(N__31360),
            .in2(_gnd_net_),
            .in3(N__31741),
            .lcout(),
            .ltout(\ALU.a_RNILVBOZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIIL3U1_15_LC_11_9_6 .C_ON=1'b0;
    defparam \ALU.c_RNIIL3U1_15_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIIL3U1_15_LC_11_9_6 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \ALU.c_RNIIL3U1_15_LC_11_9_6  (
            .in0(N__33064),
            .in1(N__34469),
            .in2(N__31349),
            .in3(N__31346),
            .lcout(),
            .ltout(\ALU.operand2_7_ns_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIOTRP4_15_LC_11_9_7 .C_ON=1'b0;
    defparam \ALU.d_RNIOTRP4_15_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIOTRP4_15_LC_11_9_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \ALU.d_RNIOTRP4_15_LC_11_9_7  (
            .in0(N__32946),
            .in1(N__33449),
            .in2(N__31340),
            .in3(N__31337),
            .lcout(\ALU.operand2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_10_LC_11_10_0 .C_ON=1'b0;
    defparam \ALU.c_10_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.c_10_LC_11_10_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.c_10_LC_11_10_0  (
            .in0(N__48561),
            .in1(N__34346),
            .in2(N__46152),
            .in3(N__34402),
            .lcout(\ALU.cZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(N__31497),
            .sr(_gnd_net_));
    defparam \ALU.c_11_LC_11_10_1 .C_ON=1'b0;
    defparam \ALU.c_11_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \ALU.c_11_LC_11_10_1 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.c_11_LC_11_10_1  (
            .in0(N__48483),
            .in1(N__34249),
            .in2(N__46156),
            .in3(N__34167),
            .lcout(\ALU.cZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(N__31497),
            .sr(_gnd_net_));
    defparam \ALU.c_12_LC_11_10_2 .C_ON=1'b0;
    defparam \ALU.c_12_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.c_12_LC_11_10_2 .LUT_INIT=16'b0111010101000101;
    LogicCell40 \ALU.c_12_LC_11_10_2  (
            .in0(N__34089),
            .in1(N__48485),
            .in2(N__46153),
            .in3(N__34020),
            .lcout(\ALU.cZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(N__31497),
            .sr(_gnd_net_));
    defparam \ALU.c_13_LC_11_10_3 .C_ON=1'b0;
    defparam \ALU.c_13_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \ALU.c_13_LC_11_10_3 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.c_13_LC_11_10_3  (
            .in0(N__48484),
            .in1(N__33921),
            .in2(N__46157),
            .in3(N__33871),
            .lcout(\ALU.cZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(N__31497),
            .sr(_gnd_net_));
    defparam \ALU.c_14_LC_11_10_4 .C_ON=1'b0;
    defparam \ALU.c_14_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \ALU.c_14_LC_11_10_4 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.c_14_LC_11_10_4  (
            .in0(N__48562),
            .in1(N__33813),
            .in2(N__46154),
            .in3(N__33747),
            .lcout(\ALU.cZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(N__31497),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIND49_14_LC_11_10_5 .C_ON=1'b0;
    defparam \ALU.c_RNIND49_14_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIND49_14_LC_11_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.c_RNIND49_14_LC_11_10_5  (
            .in0(N__33685),
            .in1(N__31543),
            .in2(_gnd_net_),
            .in3(N__45081),
            .lcout(\ALU.c_RNIND49Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_15_LC_11_10_6 .C_ON=1'b0;
    defparam \ALU.c_15_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \ALU.c_15_LC_11_10_6 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \ALU.c_15_LC_11_10_6  (
            .in0(N__48563),
            .in1(N__33654),
            .in2(N__46155),
            .in3(N__33601),
            .lcout(\ALU.cZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(N__31497),
            .sr(_gnd_net_));
    defparam \ALU.c_9_LC_11_10_7 .C_ON=1'b0;
    defparam \ALU.c_9_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \ALU.c_9_LC_11_10_7 .LUT_INIT=16'b0010000011111101;
    LogicCell40 \ALU.c_9_LC_11_10_7  (
            .in0(N__46098),
            .in1(N__48564),
            .in2(N__36202),
            .in3(N__36259),
            .lcout(\ALU.cZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(N__31497),
            .sr(_gnd_net_));
    defparam \ALU.h_1_LC_11_11_0 .C_ON=1'b0;
    defparam \ALU.h_1_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \ALU.h_1_LC_11_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.h_1_LC_11_11_0  (
            .in0(N__36606),
            .in1(N__48095),
            .in2(_gnd_net_),
            .in3(N__40981),
            .lcout(\ALU.hZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47646),
            .ce(N__45568),
            .sr(_gnd_net_));
    defparam \ALU.h_2_LC_11_11_1 .C_ON=1'b0;
    defparam \ALU.h_2_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \ALU.h_2_LC_11_11_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.h_2_LC_11_11_1  (
            .in0(N__48094),
            .in1(N__42150),
            .in2(_gnd_net_),
            .in3(N__42072),
            .lcout(\ALU.hZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47646),
            .ce(N__45568),
            .sr(_gnd_net_));
    defparam \ALU.h_3_LC_11_11_2 .C_ON=1'b0;
    defparam \ALU.h_3_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \ALU.h_3_LC_11_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.h_3_LC_11_11_2  (
            .in0(N__49460),
            .in1(N__48096),
            .in2(_gnd_net_),
            .in3(N__49382),
            .lcout(\ALU.hZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47646),
            .ce(N__45568),
            .sr(_gnd_net_));
    defparam \ALU.h_7_LC_11_11_3 .C_ON=1'b0;
    defparam \ALU.h_7_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \ALU.h_7_LC_11_11_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.h_7_LC_11_11_3  (
            .in0(N__48788),
            .in1(N__48700),
            .in2(_gnd_net_),
            .in3(N__48571),
            .lcout(\ALU.hZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47646),
            .ce(N__45568),
            .sr(_gnd_net_));
    defparam \ALU.h_5_LC_11_11_4 .C_ON=1'b0;
    defparam \ALU.h_5_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \ALU.h_5_LC_11_11_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.h_5_LC_11_11_4  (
            .in0(N__48570),
            .in1(N__49122),
            .in2(_gnd_net_),
            .in3(N__49027),
            .lcout(\ALU.hZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47646),
            .ce(N__45568),
            .sr(_gnd_net_));
    defparam \ALU.a_13_LC_11_12_0 .C_ON=1'b0;
    defparam \ALU.a_13_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.a_13_LC_11_12_0 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.a_13_LC_11_12_0  (
            .in0(N__48565),
            .in1(N__33920),
            .in2(N__46201),
            .in3(N__33880),
            .lcout(\ALU.aZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47652),
            .ce(N__44884),
            .sr(_gnd_net_));
    defparam \ALU.a_14_LC_11_12_1 .C_ON=1'b0;
    defparam \ALU.a_14_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.a_14_LC_11_12_1 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.a_14_LC_11_12_1  (
            .in0(N__48574),
            .in1(N__33817),
            .in2(N__46200),
            .in3(N__33758),
            .lcout(\ALU.aZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47652),
            .ce(N__44884),
            .sr(_gnd_net_));
    defparam \ALU.a_15_LC_11_12_2 .C_ON=1'b0;
    defparam \ALU.a_15_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.a_15_LC_11_12_2 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \ALU.a_15_LC_11_12_2  (
            .in0(N__48566),
            .in1(N__33662),
            .in2(N__46202),
            .in3(N__33603),
            .lcout(\ALU.aZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47652),
            .ce(N__44884),
            .sr(_gnd_net_));
    defparam \ALU.f_RNI0P6L_1_LC_11_12_3 .C_ON=1'b0;
    defparam \ALU.f_RNI0P6L_1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNI0P6L_1_LC_11_12_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ALU.f_RNI0P6L_1_LC_11_12_3  (
            .in0(N__36623),
            .in1(_gnd_net_),
            .in2(N__35581),
            .in3(N__36467),
            .lcout(\ALU.f_RNI0P6LZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNICQEJ_1_LC_11_12_4 .C_ON=1'b0;
    defparam \ALU.f_RNICQEJ_1_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNICQEJ_1_LC_11_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.f_RNICQEJ_1_LC_11_12_4  (
            .in0(N__36466),
            .in1(N__36622),
            .in2(_gnd_net_),
            .in3(N__32015),
            .lcout(\ALU.f_RNICQEJZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIQCLL_7_LC_11_12_5 .C_ON=1'b0;
    defparam \ALU.g_RNIQCLL_7_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIQCLL_7_LC_11_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_RNIQCLL_7_LC_11_12_5  (
            .in0(N__32014),
            .in1(N__31807),
            .in2(_gnd_net_),
            .in3(N__31690),
            .lcout(\ALU.g_RNIQCLLZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIL2FJ_5_LC_11_12_6 .C_ON=1'b0;
    defparam \ALU.f_RNIL2FJ_5_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIL2FJ_5_LC_11_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.f_RNIL2FJ_5_LC_11_12_6  (
            .in0(N__36433),
            .in1(N__48964),
            .in2(_gnd_net_),
            .in3(N__45103),
            .lcout(\ALU.f_RNIL2FJZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.m286_ns_LC_11_12_7 .C_ON=1'b0;
    defparam \ALU.m286_ns_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU.m286_ns_LC_11_12_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.m286_ns_LC_11_12_7  (
            .in0(N__31646),
            .in1(N__33359),
            .in2(_gnd_net_),
            .in3(N__31628),
            .lcout(N_287_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_2_rep1_LC_11_13_0 .C_ON=1'b0;
    defparam \CONTROL.operand2_2_rep1_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_2_rep1_LC_11_13_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \CONTROL.operand2_2_rep1_LC_11_13_0  (
            .in0(N__34686),
            .in1(N__34769),
            .in2(N__32065),
            .in3(N__32228),
            .lcout(aluOperand2_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47658),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIAOEJ_0_LC_11_13_4 .C_ON=1'b0;
    defparam \ALU.f_RNIAOEJ_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIAOEJ_0_LC_11_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.f_RNIAOEJ_0_LC_11_13_4  (
            .in0(N__35044),
            .in1(N__36286),
            .in2(_gnd_net_),
            .in3(N__32040),
            .lcout(\ALU.f_RNIAOEJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_fast_0_LC_11_13_6 .C_ON=1'b0;
    defparam \CONTROL.operand2_fast_0_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_fast_0_LC_11_13_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \CONTROL.operand2_fast_0_LC_11_13_6  (
            .in0(N__34687),
            .in1(N__34770),
            .in2(N__31593),
            .in3(N__41114),
            .lcout(aluOperand2_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47658),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIESEJ_2_LC_11_13_7 .C_ON=1'b0;
    defparam \ALU.f_RNIESEJ_2_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIESEJ_2_LC_11_13_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_RNIESEJ_2_LC_11_13_7  (
            .in0(N__32039),
            .in1(N__36451),
            .in2(_gnd_net_),
            .in3(N__31964),
            .lcout(\ALU.f_RNIESEJZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_0_LC_11_14_0 .C_ON=1'b0;
    defparam \ALU.g_0_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \ALU.g_0_LC_11_14_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_0_LC_11_14_0  (
            .in0(N__48622),
            .in1(N__42298),
            .in2(_gnd_net_),
            .in3(N__42265),
            .lcout(\ALU.gZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__36100),
            .sr(_gnd_net_));
    defparam \ALU.g_1_LC_11_14_1 .C_ON=1'b0;
    defparam \ALU.g_1_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \ALU.g_1_LC_11_14_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.g_1_LC_11_14_1  (
            .in0(N__40999),
            .in1(N__48624),
            .in2(_gnd_net_),
            .in3(N__36592),
            .lcout(\ALU.gZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__36100),
            .sr(_gnd_net_));
    defparam \ALU.g_2_LC_11_14_2 .C_ON=1'b0;
    defparam \ALU.g_2_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \ALU.g_2_LC_11_14_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.g_2_LC_11_14_2  (
            .in0(N__42161),
            .in1(N__48628),
            .in2(_gnd_net_),
            .in3(N__42097),
            .lcout(\ALU.gZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__36100),
            .sr(_gnd_net_));
    defparam \ALU.g_3_LC_11_14_3 .C_ON=1'b0;
    defparam \ALU.g_3_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \ALU.g_3_LC_11_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_3_LC_11_14_3  (
            .in0(N__48626),
            .in1(N__49469),
            .in2(_gnd_net_),
            .in3(N__49383),
            .lcout(\ALU.gZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__36100),
            .sr(_gnd_net_));
    defparam \ALU.g_4_LC_11_14_4 .C_ON=1'b0;
    defparam \ALU.g_4_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \ALU.g_4_LC_11_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_4_LC_11_14_4  (
            .in0(N__48623),
            .in1(N__49288),
            .in2(_gnd_net_),
            .in3(N__49204),
            .lcout(\ALU.gZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__36100),
            .sr(_gnd_net_));
    defparam \ALU.g_5_LC_11_14_5 .C_ON=1'b0;
    defparam \ALU.g_5_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \ALU.g_5_LC_11_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.g_5_LC_11_14_5  (
            .in0(N__48627),
            .in1(N__49123),
            .in2(_gnd_net_),
            .in3(N__49048),
            .lcout(\ALU.gZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__36100),
            .sr(_gnd_net_));
    defparam \ALU.g_7_LC_11_14_7 .C_ON=1'b0;
    defparam \ALU.g_7_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \ALU.g_7_LC_11_14_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.g_7_LC_11_14_7  (
            .in0(N__48787),
            .in1(N__48625),
            .in2(_gnd_net_),
            .in3(N__48714),
            .lcout(\ALU.gZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__36100),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJ17GT_15_LC_12_3_2 .C_ON=1'b0;
    defparam \ALU.c_RNIJ17GT_15_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJ17GT_15_LC_12_3_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIJ17GT_15_LC_12_3_2  (
            .in0(N__38735),
            .in1(N__31783),
            .in2(_gnd_net_),
            .in3(N__31772),
            .lcout(\ALU.N_634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_12_3_4 .C_ON=1'b0;
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_2_c_inv_LC_12_3_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \FTDI.un3_TX_cry_2_c_inv_LC_12_3_4  (
            .in0(N__32363),
            .in1(N__36517),
            .in2(_gnd_net_),
            .in3(N__32326),
            .lcout(\FTDI.un3_TX_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_12_LC_12_4_4.C_ON=1'b0;
    defparam testWord_12_LC_12_4_4.SEQ_MODE=4'b1000;
    defparam testWord_12_LC_12_4_4.LUT_INIT=16'b1110001011110000;
    LogicCell40 testWord_12_LC_12_4_4 (
            .in0(N__32294),
            .in1(N__41467),
            .in2(N__32184),
            .in3(N__41220),
            .lcout(testWordZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47605),
            .ce(N__41063),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_0_LC_12_5_0 .C_ON=1'b0;
    defparam \FTDI.TXshift_0_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_0_LC_12_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_0_LC_12_5_0  (
            .in0(N__44754),
            .in1(N__44675),
            .in2(_gnd_net_),
            .in3(N__32153),
            .lcout(\FTDI.TXshiftZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__44659),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_5_LC_12_5_1 .C_ON=1'b0;
    defparam \FTDI.TXshift_5_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_5_LC_12_5_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_5_LC_12_5_1  (
            .in0(N__32087),
            .in1(N__44612),
            .in2(_gnd_net_),
            .in3(N__44758),
            .lcout(\FTDI.TXshiftZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__44659),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_3_LC_12_5_3 .C_ON=1'b0;
    defparam \FTDI.TXshift_3_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_3_LC_12_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_3_LC_12_5_3  (
            .in0(N__32120),
            .in1(N__32144),
            .in2(_gnd_net_),
            .in3(N__44756),
            .lcout(\FTDI.TXshiftZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__44659),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_4_LC_12_5_4 .C_ON=1'b0;
    defparam \FTDI.TXshift_4_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_4_LC_12_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_4_LC_12_5_4  (
            .in0(N__44757),
            .in1(N__32135),
            .in2(_gnd_net_),
            .in3(N__32129),
            .lcout(\FTDI.TXshiftZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__44659),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_2_LC_12_5_5 .C_ON=1'b0;
    defparam \FTDI.TXshift_2_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_2_LC_12_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_2_LC_12_5_5  (
            .in0(N__32111),
            .in1(N__32105),
            .in2(_gnd_net_),
            .in3(N__44755),
            .lcout(\FTDI.TXshiftZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__44659),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_6_LC_12_5_6 .C_ON=1'b0;
    defparam \FTDI.TXshift_6_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_6_LC_12_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \FTDI.TXshift_6_LC_12_5_6  (
            .in0(N__44759),
            .in1(N__32558),
            .in2(_gnd_net_),
            .in3(N__32096),
            .lcout(\FTDI.TXshiftZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__44659),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_7_LC_12_5_7 .C_ON=1'b0;
    defparam \FTDI.TXshift_7_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_7_LC_12_5_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \FTDI.TXshift_7_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__32567),
            .in2(_gnd_net_),
            .in3(N__44753),
            .lcout(\FTDI.TXshiftZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_0C_net ),
            .ce(N__44659),
            .sr(_gnd_net_));
    defparam \ALU.un2_addsub_cry_10_c_RNIEBKOT_LC_12_6_0 .C_ON=1'b0;
    defparam \ALU.un2_addsub_cry_10_c_RNIEBKOT_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un2_addsub_cry_10_c_RNIEBKOT_LC_12_6_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \ALU.un2_addsub_cry_10_c_RNIEBKOT_LC_12_6_0  (
            .in0(N__42517),
            .in1(N__39212),
            .in2(_gnd_net_),
            .in3(N__32552),
            .lcout(un2_addsub_cry_10_c_RNIEBKOT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_11_LC_12_6_1 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_11_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_11_LC_12_6_1 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \ALU.a_15_m2_ns_1_11_LC_12_6_1  (
            .in0(N__43754),
            .in1(N__47259),
            .in2(N__43939),
            .in3(N__44203),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI55HKC_11_LC_12_6_2 .C_ON=1'b0;
    defparam \ALU.c_RNI55HKC_11_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI55HKC_11_LC_12_6_2 .LUT_INIT=16'b0110011110000110;
    LogicCell40 \ALU.c_RNI55HKC_11_LC_12_6_2  (
            .in0(N__47260),
            .in1(N__39368),
            .in2(N__32537),
            .in3(N__39476),
            .lcout(),
            .ltout(\ALU.a_15_m2_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIPTRDR1_11_LC_12_6_3 .C_ON=1'b0;
    defparam \ALU.c_RNIPTRDR1_11_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIPTRDR1_11_LC_12_6_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNIPTRDR1_11_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__44204),
            .in2(N__32534),
            .in3(N__32531),
            .lcout(),
            .ltout(\ALU.a_15_m4_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNID7K8N2_11_LC_12_6_4 .C_ON=1'b0;
    defparam \ALU.c_RNID7K8N2_11_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNID7K8N2_11_LC_12_6_4 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \ALU.c_RNID7K8N2_11_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__46353),
            .in2(N__32516),
            .in3(N__32513),
            .lcout(),
            .ltout(c_RNID7K8N2_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperation_RNI5QD2L3_0_LC_12_6_5 .C_ON=1'b0;
    defparam \CONTROL.aluOperation_RNI5QD2L3_0_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \CONTROL.aluOperation_RNI5QD2L3_0_LC_12_6_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \CONTROL.aluOperation_RNI5QD2L3_0_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__48269),
            .in2(N__32501),
            .in3(N__32498),
            .lcout(aluOperation_RNI5QD2L3_0),
            .ltout(aluOperation_RNI5QD2L3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_11_LC_12_6_6 .C_ON=1'b0;
    defparam \ALU.a_11_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \ALU.a_11_LC_12_6_6 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \ALU.a_11_LC_12_6_6  (
            .in0(N__48270),
            .in1(N__46040),
            .in2(N__32492),
            .in3(N__34181),
            .lcout(\ALU.aZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47611),
            .ce(N__44872),
            .sr(_gnd_net_));
    defparam \ALU.e_9_LC_12_7_0 .C_ON=1'b0;
    defparam \ALU.e_9_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \ALU.e_9_LC_12_7_0 .LUT_INIT=16'b0010000011111101;
    LogicCell40 \ALU.e_9_LC_12_7_0  (
            .in0(N__45992),
            .in1(N__48328),
            .in2(N__36209),
            .in3(N__36258),
            .lcout(\ALU.eZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47615),
            .ce(N__32435),
            .sr(_gnd_net_));
    defparam \ALU.g_RNIVGLL_9_LC_12_7_2 .C_ON=1'b0;
    defparam \ALU.g_RNIVGLL_9_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.g_RNIVGLL_9_LC_12_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.g_RNIVGLL_9_LC_12_7_2  (
            .in0(N__36123),
            .in1(N__32715),
            .in2(_gnd_net_),
            .in3(N__45112),
            .lcout(),
            .ltout(\ALU.g_RNIVGLLZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIURH32_9_LC_12_7_3 .C_ON=1'b0;
    defparam \ALU.e_RNIURH32_9_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIURH32_9_LC_12_7_3 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \ALU.e_RNIURH32_9_LC_12_7_3  (
            .in0(N__33062),
            .in1(N__34475),
            .in2(N__32852),
            .in3(N__38345),
            .lcout(\ALU.operand2_7_ns_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_m2_0_1_LC_12_7_4 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_m2_0_1_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_m2_0_1_LC_12_7_4 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \ALU.mult_g0_0_0_m2_0_1_LC_12_7_4  (
            .in0(N__45321),
            .in1(N__38364),
            .in2(N__38401),
            .in3(N__35032),
            .lcout(\ALU.g0_0_0_m2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_m2_LC_12_7_5 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_m2_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_m2_LC_12_7_5 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.mult_g0_0_0_m2_LC_12_7_5  (
            .in0(N__32840),
            .in1(N__32796),
            .in2(N__32759),
            .in3(N__34474),
            .lcout(),
            .ltout(\ALU.N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_m4_LC_12_7_6 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_m4_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_m4_LC_12_7_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \ALU.mult_g0_0_0_m4_LC_12_7_6  (
            .in0(N__32684),
            .in1(_gnd_net_),
            .in2(N__32741),
            .in3(N__32970),
            .lcout(\ALU.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_g0_0_0_m2_0_LC_12_7_7 .C_ON=1'b0;
    defparam \ALU.mult_g0_0_0_m2_0_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_g0_0_0_m2_0_LC_12_7_7 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.mult_g0_0_0_m2_0_LC_12_7_7  (
            .in0(N__32716),
            .in1(N__34473),
            .in2(N__32693),
            .in3(N__36124),
            .lcout(\ALU.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_15_LC_12_8_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_15_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_15_LC_12_8_0 .LUT_INIT=16'b0011010100111111;
    LogicCell40 \ALU.a_15_m2_ns_1_15_LC_12_8_0  (
            .in0(N__44205),
            .in1(N__43937),
            .in2(N__47321),
            .in3(N__43675),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIMPCHC_15_LC_12_8_1 .C_ON=1'b0;
    defparam \ALU.c_RNIMPCHC_15_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIMPCHC_15_LC_12_8_1 .LUT_INIT=16'b0110011110000110;
    LogicCell40 \ALU.c_RNIMPCHC_15_LC_12_8_1  (
            .in0(N__47314),
            .in1(N__32674),
            .in2(N__32618),
            .in3(N__32615),
            .lcout(),
            .ltout(\ALU.a_15_m2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIM5JEB2_15_LC_12_8_2 .C_ON=1'b0;
    defparam \ALU.c_RNIM5JEB2_15_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIM5JEB2_15_LC_12_8_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.c_RNIM5JEB2_15_LC_12_8_2  (
            .in0(N__44206),
            .in1(_gnd_net_),
            .in2(N__32585),
            .in3(N__32582),
            .lcout(),
            .ltout(\ALU.a_15_m4_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIR4QHM2_15_LC_12_8_3 .C_ON=1'b0;
    defparam \ALU.c_RNIR4QHM2_15_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIR4QHM2_15_LC_12_8_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.c_RNIR4QHM2_15_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__46352),
            .in2(N__33521),
            .in3(N__33518),
            .lcout(),
            .ltout(\ALU.c_RNIR4QHM2Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_14_c_RNI1G6N93_LC_12_8_4 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_14_c_RNI1G6N93_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_14_c_RNI1G6N93_LC_12_8_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.un9_addsub_cry_14_c_RNI1G6N93_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__48273),
            .in2(N__33506),
            .in3(N__40487),
            .lcout(\ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93 ),
            .ltout(\ALU.un9_addsub_cry_14_c_RNI1G6NZ0Z93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_15_LC_12_8_5 .C_ON=1'b0;
    defparam \ALU.h_15_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \ALU.h_15_LC_12_8_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \ALU.h_15_LC_12_8_5  (
            .in0(N__48274),
            .in1(N__45903),
            .in2(N__33503),
            .in3(N__33604),
            .lcout(\ALU.hZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47621),
            .ce(N__45572),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISBLU_15_LC_12_8_6 .C_ON=1'b0;
    defparam \ALU.d_RNISBLU_15_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISBLU_15_LC_12_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNISBLU_15_LC_12_8_6  (
            .in0(N__33487),
            .in1(N__33472),
            .in2(_gnd_net_),
            .in3(N__45299),
            .lcout(\ALU.d_RNISBLUZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.aluOperationZ0Z_5_LC_12_9_1 .C_ON=1'b0;
    defparam \CONTROL.aluOperationZ0Z_5_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \CONTROL.aluOperationZ0Z_5_LC_12_9_1 .LUT_INIT=16'b1110111001001110;
    LogicCell40 \CONTROL.aluOperationZ0Z_5_LC_12_9_1  (
            .in0(N__33443),
            .in1(N__33163),
            .in2(N__33395),
            .in3(N__33354),
            .lcout(aluOperation_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47628),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_1_l_ofx_LC_12_9_2 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_1_l_ofx_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_1_l_ofx_LC_12_9_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \ALU.mult_madd_axb_1_l_ofx_LC_12_9_2  (
            .in0(N__37796),
            .in1(N__33149),
            .in2(N__37786),
            .in3(N__37479),
            .lcout(\ALU.madd_axb_1_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_0_rep2_LC_12_9_4 .C_ON=1'b0;
    defparam \CONTROL.operand2_0_rep2_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_0_rep2_LC_12_9_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \CONTROL.operand2_0_rep2_LC_12_9_4  (
            .in0(N__34714),
            .in1(N__34796),
            .in2(N__41113),
            .in3(N__33048),
            .lcout(aluOperand2_0_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47628),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_0_LC_12_9_5 .C_ON=1'b0;
    defparam \CONTROL.operand2_0_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_0_LC_12_9_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \CONTROL.operand2_0_LC_12_9_5  (
            .in0(N__34794),
            .in1(N__34715),
            .in2(N__32959),
            .in3(N__41107),
            .lcout(aluOperand2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47628),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIEFIJ_10_LC_12_9_6 .C_ON=1'b0;
    defparam \ALU.c_RNIEFIJ_10_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIEFIJ_10_LC_12_9_6 .LUT_INIT=16'b0000101001110111;
    LogicCell40 \ALU.c_RNIEFIJ_10_LC_12_9_6  (
            .in0(N__35029),
            .in1(N__34917),
            .in2(N__34269),
            .in3(N__34882),
            .lcout(\ALU.g0_7_m4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CONTROL.operand2_1_LC_12_9_7 .C_ON=1'b0;
    defparam \CONTROL.operand2_1_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \CONTROL.operand2_1_LC_12_9_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \CONTROL.operand2_1_LC_12_9_7  (
            .in0(N__34795),
            .in1(N__34716),
            .in2(N__34568),
            .in3(N__34488),
            .lcout(aluOperand2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47628),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.g_10_LC_12_10_0 .C_ON=1'b0;
    defparam \ALU.g_10_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \ALU.g_10_LC_12_10_0 .LUT_INIT=16'b0100000011101111;
    LogicCell40 \ALU.g_10_LC_12_10_0  (
            .in0(N__48486),
            .in1(N__34403),
            .in2(N__46158),
            .in3(N__34342),
            .lcout(\ALU.gZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47635),
            .ce(N__36093),
            .sr(_gnd_net_));
    defparam \ALU.g_11_LC_12_10_1 .C_ON=1'b0;
    defparam \ALU.g_11_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \ALU.g_11_LC_12_10_1 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.g_11_LC_12_10_1  (
            .in0(N__48490),
            .in1(N__34214),
            .in2(N__46000),
            .in3(N__34179),
            .lcout(\ALU.gZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47635),
            .ce(N__36093),
            .sr(_gnd_net_));
    defparam \ALU.g_12_LC_12_10_2 .C_ON=1'b0;
    defparam \ALU.g_12_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \ALU.g_12_LC_12_10_2 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.g_12_LC_12_10_2  (
            .in0(N__48487),
            .in1(N__34091),
            .in2(N__46159),
            .in3(N__34025),
            .lcout(\ALU.gZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47635),
            .ce(N__36093),
            .sr(_gnd_net_));
    defparam \ALU.g_13_LC_12_10_3 .C_ON=1'b0;
    defparam \ALU.g_13_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \ALU.g_13_LC_12_10_3 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.g_13_LC_12_10_3  (
            .in0(N__48491),
            .in1(N__33939),
            .in2(N__46001),
            .in3(N__33872),
            .lcout(\ALU.gZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47635),
            .ce(N__36093),
            .sr(_gnd_net_));
    defparam \ALU.g_14_LC_12_10_4 .C_ON=1'b0;
    defparam \ALU.g_14_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \ALU.g_14_LC_12_10_4 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.g_14_LC_12_10_4  (
            .in0(N__48488),
            .in1(N__33818),
            .in2(N__46160),
            .in3(N__33748),
            .lcout(\ALU.gZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47635),
            .ce(N__36093),
            .sr(_gnd_net_));
    defparam \ALU.g_15_LC_12_10_5 .C_ON=1'b0;
    defparam \ALU.g_15_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \ALU.g_15_LC_12_10_5 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \ALU.g_15_LC_12_10_5  (
            .in0(N__48492),
            .in1(N__33653),
            .in2(N__46002),
            .in3(N__33605),
            .lcout(\ALU.gZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47635),
            .ce(N__36093),
            .sr(_gnd_net_));
    defparam \ALU.g_9_LC_12_10_6 .C_ON=1'b0;
    defparam \ALU.g_9_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \ALU.g_9_LC_12_10_6 .LUT_INIT=16'b0111001100100011;
    LogicCell40 \ALU.g_9_LC_12_10_6  (
            .in0(N__48489),
            .in1(N__36264),
            .in2(N__46161),
            .in3(N__36195),
            .lcout(\ALU.gZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47635),
            .ce(N__36093),
            .sr(_gnd_net_));
    defparam \ALU.a_RNI85LF1_13_LC_12_11_0 .C_ON=1'b0;
    defparam \ALU.a_RNI85LF1_13_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_RNI85LF1_13_LC_12_11_0 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \ALU.a_RNI85LF1_13_LC_12_11_0  (
            .in0(N__36038),
            .in1(N__36019),
            .in2(N__36003),
            .in3(N__35898),
            .lcout(),
            .ltout(\ALU.dout_3_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIFEHQ1_13_LC_12_11_1 .C_ON=1'b0;
    defparam \ALU.c_RNIFEHQ1_13_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIFEHQ1_13_LC_12_11_1 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \ALU.c_RNIFEHQ1_13_LC_12_11_1  (
            .in0(N__35810),
            .in1(N__35377),
            .in2(N__35798),
            .in3(N__35795),
            .lcout(\ALU.N_712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_RNIRBBD1_13_LC_12_11_2 .C_ON=1'b0;
    defparam \ALU.b_RNIRBBD1_13_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.b_RNIRBBD1_13_LC_12_11_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \ALU.b_RNIRBBD1_13_LC_12_11_2  (
            .in0(N__35781),
            .in1(N__35752),
            .in2(N__35615),
            .in3(N__35532),
            .lcout(),
            .ltout(\ALU.dout_6_ns_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI4TJ02_13_LC_12_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNI4TJ02_13_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI4TJ02_13_LC_12_11_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \ALU.d_RNI4TJ02_13_LC_12_11_3  (
            .in0(N__35462),
            .in1(N__35434),
            .in2(N__35405),
            .in3(N__35378),
            .lcout(),
            .ltout(\ALU.N_760_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNINMUU3_13_LC_12_11_4 .C_ON=1'b0;
    defparam \ALU.c_RNINMUU3_13_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNINMUU3_13_LC_12_11_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \ALU.c_RNINMUU3_13_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__35252),
            .in2(N__35246),
            .in3(N__35229),
            .lcout(\ALU.aluOut_13 ),
            .ltout(\ALU.aluOut_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNI7KNC7_13_LC_12_11_5 .C_ON=1'b0;
    defparam \ALU.c_RNI7KNC7_13_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNI7KNC7_13_LC_12_11_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.c_RNI7KNC7_13_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35072),
            .in3(N__38325),
            .lcout(\ALU.a13_b_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.f_0_LC_12_12_0 .C_ON=1'b0;
    defparam \ALU.f_0_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.f_0_LC_12_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_0_LC_12_12_0  (
            .in0(N__48493),
            .in1(N__42296),
            .in2(_gnd_net_),
            .in3(N__42266),
            .lcout(\ALU.fZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.f_1_LC_12_12_1 .C_ON=1'b0;
    defparam \ALU.f_1_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.f_1_LC_12_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_1_LC_12_12_1  (
            .in0(N__48582),
            .in1(N__40959),
            .in2(_gnd_net_),
            .in3(N__36591),
            .lcout(\ALU.fZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.f_2_LC_12_12_2 .C_ON=1'b0;
    defparam \ALU.f_2_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.f_2_LC_12_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_2_LC_12_12_2  (
            .in0(N__48494),
            .in1(N__42146),
            .in2(_gnd_net_),
            .in3(N__42096),
            .lcout(\ALU.fZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.f_3_LC_12_12_3 .C_ON=1'b0;
    defparam \ALU.f_3_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.f_3_LC_12_12_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.f_3_LC_12_12_3  (
            .in0(N__49361),
            .in1(N__48496),
            .in2(_gnd_net_),
            .in3(N__49442),
            .lcout(\ALU.fZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.f_4_LC_12_12_4 .C_ON=1'b0;
    defparam \ALU.f_4_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.f_4_LC_12_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.f_4_LC_12_12_4  (
            .in0(N__49212),
            .in1(N__48584),
            .in2(_gnd_net_),
            .in3(N__49262),
            .lcout(\ALU.fZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.f_5_LC_12_12_5 .C_ON=1'b0;
    defparam \ALU.f_5_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.f_5_LC_12_12_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.f_5_LC_12_12_5  (
            .in0(N__49090),
            .in1(N__48497),
            .in2(_gnd_net_),
            .in3(N__49043),
            .lcout(\ALU.fZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.f_6_LC_12_12_6 .C_ON=1'b0;
    defparam \ALU.f_6_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \ALU.f_6_LC_12_12_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_6_LC_12_12_6  (
            .in0(N__48495),
            .in1(N__48867),
            .in2(_gnd_net_),
            .in3(N__48931),
            .lcout(\ALU.fZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.f_7_LC_12_12_7 .C_ON=1'b0;
    defparam \ALU.f_7_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \ALU.f_7_LC_12_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_7_LC_12_12_7  (
            .in0(N__48583),
            .in1(N__48789),
            .in2(_gnd_net_),
            .in3(N__48696),
            .lcout(\ALU.fZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(N__36380),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIO75MA_0_LC_12_13_1 .C_ON=1'b0;
    defparam \ALU.d_RNIO75MA_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIO75MA_0_LC_12_13_1 .LUT_INIT=16'b0101100110101001;
    LogicCell40 \ALU.d_RNIO75MA_0_LC_12_13_1  (
            .in0(N__38037),
            .in1(N__36329),
            .in2(N__42526),
            .in3(N__38248),
            .lcout(\ALU.d_RNIO75MAZ0Z_0 ),
            .ltout(\ALU.d_RNIO75MAZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_0_LC_12_13_2 .C_ON=1'b0;
    defparam \ALU.b_0_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \ALU.b_0_LC_12_13_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.b_0_LC_12_13_2  (
            .in0(N__48590),
            .in1(_gnd_net_),
            .in2(N__36302),
            .in3(N__42253),
            .lcout(\ALU.bZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47653),
            .ce(N__47397),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_0_l_ofx_LC_12_13_4 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_0_l_ofx_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_0_l_ofx_LC_12_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALU.mult_madd_axb_0_l_ofx_LC_12_13_4  (
            .in0(N__38249),
            .in1(N__38036),
            .in2(N__37502),
            .in3(N__37762),
            .lcout(\ALU.madd_axb_0_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.mult_madd_axb_0_LC_12_13_5 .C_ON=1'b0;
    defparam \ALU.mult_madd_axb_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU.mult_madd_axb_0_LC_12_13_5 .LUT_INIT=16'b0110110010100000;
    LogicCell40 \ALU.mult_madd_axb_0_LC_12_13_5  (
            .in0(N__37763),
            .in1(N__37480),
            .in2(N__38047),
            .in3(N__38247),
            .lcout(),
            .ltout(\ALU.mult_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIEICQ63_1_LC_12_13_6 .C_ON=1'b0;
    defparam \ALU.d_RNIEICQ63_1_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIEICQ63_1_LC_12_13_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIEICQ63_1_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__46004),
            .in2(N__36647),
            .in3(N__36644),
            .lcout(\ALU.d_RNIEICQ63Z0Z_1 ),
            .ltout(\ALU.d_RNIEICQ63Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_1_LC_12_13_7 .C_ON=1'b0;
    defparam \ALU.b_1_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \ALU.b_1_LC_12_13_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.b_1_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__48589),
            .in2(N__36626),
            .in3(N__40979),
            .lcout(\ALU.bZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47653),
            .ce(N__47397),
            .sr(_gnd_net_));
    defparam \ALU.d_1_LC_12_14_7 .C_ON=1'b0;
    defparam \ALU.d_1_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \ALU.d_1_LC_12_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_1_LC_12_14_7  (
            .in0(N__48591),
            .in1(N__40980),
            .in2(_gnd_net_),
            .in3(N__36590),
            .lcout(\ALU.dZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47659),
            .ce(N__43344),
            .sr(_gnd_net_));
    defparam \ALU.h_4_LC_12_16_3 .C_ON=1'b0;
    defparam \ALU.h_4_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \ALU.h_4_LC_12_16_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.h_4_LC_12_16_3  (
            .in0(N__49213),
            .in1(N__48588),
            .in2(_gnd_net_),
            .in3(N__49289),
            .lcout(\ALU.hZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47673),
            .ce(N__45573),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_2_c_LC_13_2_0 .C_ON=1'b1;
    defparam \FTDI.un3_TX_cry_2_c_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_2_c_LC_13_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \FTDI.un3_TX_cry_2_c_LC_13_2_0  (
            .in0(_gnd_net_),
            .in1(N__36518),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_2_0_),
            .carryout(\FTDI.un3_TX_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_13_2_1 .C_ON=1'b1;
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_13_2_1 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_3_c_inv_LC_13_2_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \FTDI.un3_TX_cry_3_c_inv_LC_13_2_1  (
            .in0(_gnd_net_),
            .in1(N__36506),
            .in2(_gnd_net_),
            .in3(N__44771),
            .lcout(\FTDI.un3_TX_axb_3 ),
            .ltout(),
            .carryin(\FTDI.un3_TX_cry_2 ),
            .carryout(\FTDI.un3_TX_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_13_2_2 .C_ON=1'b0;
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_13_2_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \FTDI.un3_TX_cry_3_c_RNIBAJU_LC_13_2_2  (
            .in0(N__44770),
            .in1(N__36500),
            .in2(_gnd_net_),
            .in3(N__36488),
            .lcout(FTDI_TX_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIU2HCP_0_LC_13_5_1 .C_ON=1'b0;
    defparam \ALU.d_RNIU2HCP_0_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIU2HCP_0_LC_13_5_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNIU2HCP_0_LC_13_5_1  (
            .in0(N__38744),
            .in1(N__39199),
            .in2(_gnd_net_),
            .in3(N__39181),
            .lcout(\ALU.N_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIMGKHG_13_LC_13_6_4 .C_ON=1'b0;
    defparam \ALU.c_RNIMGKHG_13_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIMGKHG_13_LC_13_6_4 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ALU.c_RNIMGKHG_13_LC_13_6_4  (
            .in0(N__39070),
            .in1(N__38765),
            .in2(N__38739),
            .in3(N__38444),
            .lcout(\ALU.rshift_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.e_RNIR49H_9_LC_13_6_7 .C_ON=1'b0;
    defparam \ALU.e_RNIR49H_9_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \ALU.e_RNIR49H_9_LC_13_6_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \ALU.e_RNIR49H_9_LC_13_6_7  (
            .in0(N__38391),
            .in1(N__38371),
            .in2(N__45135),
            .in3(_gnd_net_),
            .lcout(\ALU.e_RNIR49HZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIKQQR6_0_LC_13_7_0 .C_ON=1'b1;
    defparam \ALU.d_RNIKQQR6_0_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIKQQR6_0_LC_13_7_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALU.d_RNIKQQR6_0_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__38338),
            .in2(N__38051),
            .in3(N__37254),
            .lcout(\ALU.a0_b_2 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\ALU.un9_addsub_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_0_c_RNI2U096_LC_13_7_1 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_0_c_RNI2U096_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_0_c_RNI2U096_LC_13_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_0_c_RNI2U096_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__37787),
            .in2(N__37501),
            .in3(N__37259),
            .lcout(\ALU.un9_addsub_cry_0_c_RNI2UZ0Z096 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_0 ),
            .carryout(\ALU.un9_addsub_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_1_c_RNI6TD17_LC_13_7_2 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_1_c_RNI6TD17_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_1_c_RNI6TD17_LC_13_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_1_c_RNI6TD17_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__37255),
            .in2(N__37001),
            .in3(N__36698),
            .lcout(\ALU.un9_addsub_cry_1_c_RNI6TDZ0Z17 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_1 ),
            .carryout(\ALU.un9_addsub_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_2_c_RNIA3LG7_LC_13_7_3 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_2_c_RNIA3LG7_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_2_c_RNIA3LG7_LC_13_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_2_c_RNIA3LG7_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__41974),
            .in2(N__36695),
            .in3(N__36680),
            .lcout(\ALU.un9_addsub_cry_2_c_RNIA3LGZ0Z7 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_2 ),
            .carryout(\ALU.un9_addsub_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_3_c_RNI525R7_LC_13_7_4 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_3_c_RNI525R7_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_3_c_RNI525R7_LC_13_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_3_c_RNI525R7_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__42992),
            .in2(N__36677),
            .in3(N__36665),
            .lcout(\ALU.un9_addsub_cry_3_c_RNI525RZ0Z7 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_3 ),
            .carryout(\ALU.un9_addsub_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_4_c_RNIL4N97_LC_13_7_5 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_4_c_RNIL4N97_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_4_c_RNIL4N97_LC_13_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_4_c_RNIL4N97_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__40391),
            .in2(N__40223),
            .in3(N__40196),
            .lcout(\ALU.un9_addsub_cry_4_c_RNIL4NZ0Z97 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_4 ),
            .carryout(\ALU.un9_addsub_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_5_c_RNI6SCF7_LC_13_7_6 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_5_c_RNI6SCF7_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_5_c_RNI6SCF7_LC_13_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_5_c_RNI6SCF7_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__46733),
            .in2(N__40193),
            .in3(N__40175),
            .lcout(\ALU.un9_addsub_cry_5_c_RNI6SCFZ0Z7 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_5 ),
            .carryout(\ALU.un9_addsub_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_6_c_RNI2EFH8_LC_13_7_7 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_6_c_RNI2EFH8_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_6_c_RNI2EFH8_LC_13_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_6_c_RNI2EFH8_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__46976),
            .in2(N__40172),
            .in3(N__40124),
            .lcout(\ALU.un9_addsub_cry_6_c_RNI2EFHZ0Z8 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_6 ),
            .carryout(\ALU.un9_addsub_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_7_c_RNIU7F18_LC_13_8_0 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_7_c_RNIU7F18_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_7_c_RNIU7F18_LC_13_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_7_c_RNIU7F18_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__40121),
            .in2(N__39890),
            .in3(N__39863),
            .lcout(\ALU.un9_addsub_cry_7_c_RNIU7FZ0Z18 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\ALU.un9_addsub_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_8_c_RNIPV1S8_LC_13_8_1 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_8_c_RNIPV1S8_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_8_c_RNIPV1S8_LC_13_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_8_c_RNIPV1S8_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__39859),
            .in2(N__39641),
            .in3(N__39611),
            .lcout(\ALU.un9_addsub_cry_8_c_RNIPV1SZ0Z8 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_8 ),
            .carryout(\ALU.un9_addsub_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_9_c_RNI22U6K_LC_13_8_2 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_9_c_RNI22U6K_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_9_c_RNI22U6K_LC_13_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_9_c_RNI22U6K_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__39605),
            .in2(N__39506),
            .in3(N__39479),
            .lcout(\ALU.un9_addsub_cry_9_c_RNI22U6KZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_9 ),
            .carryout(\ALU.un9_addsub_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_10_c_RNI9C0K9_LC_13_8_3 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_10_c_RNI9C0K9_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_10_c_RNI9C0K9_LC_13_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_10_c_RNI9C0K9_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__39467),
            .in2(N__39398),
            .in3(N__39203),
            .lcout(\ALU.un9_addsub_cry_10_c_RNI9C0KZ0Z9 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_10 ),
            .carryout(\ALU.un9_addsub_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_11_c_RNI10BQK_LC_13_8_4 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_11_c_RNI10BQK_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_11_c_RNI10BQK_LC_13_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_11_c_RNI10BQK_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__40853),
            .in2(N__40805),
            .in3(N__40775),
            .lcout(\ALU.un9_addsub_cry_11_c_RNI10BQKZ0 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_11 ),
            .carryout(\ALU.un9_addsub_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_12_c_RNIBB5Q9_LC_13_8_5 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_12_c_RNIBB5Q9_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_12_c_RNIBB5Q9_LC_13_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_12_c_RNIBB5Q9_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__40711),
            .in2(N__40664),
            .in3(N__40637),
            .lcout(\ALU.un9_addsub_cry_12_c_RNIBB5QZ0Z9 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_12 ),
            .carryout(\ALU.un9_addsub_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_13_c_RNI4JGF9_LC_13_8_6 .C_ON=1'b1;
    defparam \ALU.un9_addsub_cry_13_c_RNI4JGF9_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_13_c_RNI4JGF9_LC_13_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU.un9_addsub_cry_13_c_RNI4JGF9_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__40634),
            .in2(N__40559),
            .in3(N__40526),
            .lcout(\ALU.un9_addsub_cry_13_c_RNI4JGFZ0Z9 ),
            .ltout(),
            .carryin(\ALU.un9_addsub_cry_13 ),
            .carryout(\ALU.un9_addsub_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_14_c_RNIS374J_LC_13_8_7 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_14_c_RNIS374J_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_14_c_RNIS374J_LC_13_8_7 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ALU.un9_addsub_cry_14_c_RNIS374J_LC_13_8_7  (
            .in0(N__42495),
            .in1(N__40523),
            .in2(N__40508),
            .in3(N__40490),
            .lcout(\ALU.un9_addsub_cry_14_c_RNIS374JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_3_LC_13_9_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_3_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_3_LC_13_9_0 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.a_15_m2_ns_1_3_LC_13_9_0  (
            .in0(N__47303),
            .in1(N__44198),
            .in2(N__43952),
            .in3(N__43761),
            .lcout(\ALU.a_15_m2_ns_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.c_RNIJK5GK1_15_LC_13_9_1 .C_ON=1'b0;
    defparam \ALU.c_RNIJK5GK1_15_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.c_RNIJK5GK1_15_LC_13_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.c_RNIJK5GK1_15_LC_13_9_1  (
            .in0(N__44527),
            .in1(N__40481),
            .in2(_gnd_net_),
            .in3(N__40466),
            .lcout(),
            .ltout(\ALU.rshift_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI3V2CP1_3_LC_13_9_2 .C_ON=1'b0;
    defparam \ALU.d_RNI3V2CP1_3_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI3V2CP1_3_LC_13_9_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \ALU.d_RNI3V2CP1_3_LC_13_9_2  (
            .in0(N__43185),
            .in1(_gnd_net_),
            .in2(N__40454),
            .in3(N__40451),
            .lcout(),
            .ltout(\ALU.d_RNI3V2CP1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBRAVJ2_3_LC_13_9_3 .C_ON=1'b0;
    defparam \ALU.d_RNIBRAVJ2_3_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBRAVJ2_3_LC_13_9_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNIBRAVJ2_3_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__46391),
            .in2(N__40436),
            .in3(N__41588),
            .lcout(\ALU.a_15_m5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJTNHA_3_LC_13_9_4 .C_ON=1'b0;
    defparam \ALU.d_RNIJTNHA_3_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJTNHA_3_LC_13_9_4 .LUT_INIT=16'b1000011001100111;
    LogicCell40 \ALU.d_RNIJTNHA_3_LC_13_9_4  (
            .in0(N__47304),
            .in1(N__42005),
            .in2(N__41747),
            .in3(N__41735),
            .lcout(),
            .ltout(\ALU.a_15_m2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI95MLP_3_LC_13_9_5 .C_ON=1'b0;
    defparam \ALU.d_RNI95MLP_3_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI95MLP_3_LC_13_9_5 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \ALU.d_RNI95MLP_3_LC_13_9_5  (
            .in0(N__44526),
            .in1(N__44202),
            .in2(N__41609),
            .in3(N__41606),
            .lcout(\ALU.d_RNI95MLPZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIE8SJN5_3_LC_13_9_6 .C_ON=1'b0;
    defparam \ALU.d_RNIE8SJN5_3_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIE8SJN5_3_LC_13_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIE8SJN5_3_LC_13_9_6  (
            .in0(N__45893),
            .in1(N__41582),
            .in2(_gnd_net_),
            .in3(N__41573),
            .lcout(\ALU.d_RNIE8SJN5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam testWord_10_LC_13_10_0.C_ON=1'b0;
    defparam testWord_10_LC_13_10_0.SEQ_MODE=4'b1000;
    defparam testWord_10_LC_13_10_0.LUT_INIT=16'b1110001011110000;
    LogicCell40 testWord_10_LC_13_10_0 (
            .in0(N__41567),
            .in1(N__41500),
            .in2(N__41108),
            .in3(N__41231),
            .lcout(testWordZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47629),
            .ce(N__41061),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_0_c_RNIEMTLK_LC_13_10_1 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_0_c_RNIEMTLK_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_0_c_RNIEMTLK_LC_13_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.un9_addsub_cry_0_c_RNIEMTLK_LC_13_10_1  (
            .in0(N__42502),
            .in1(N__41021),
            .in2(_gnd_net_),
            .in3(N__41012),
            .lcout(\ALU.un9_addsub_cry_0_c_RNIEMTLKZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_1_c_RNIM56UL_LC_13_10_2 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_1_c_RNIM56UL_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_1_c_RNIM56UL_LC_13_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.un9_addsub_cry_1_c_RNIM56UL_LC_13_10_2  (
            .in0(N__42506),
            .in1(N__40925),
            .in2(_gnd_net_),
            .in3(N__40916),
            .lcout(\ALU.un9_addsub_cry_1_c_RNIM56ULZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_2_c_RNIMN63N_LC_13_10_3 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_2_c_RNIMN63N_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_2_c_RNIMN63N_LC_13_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.un9_addsub_cry_2_c_RNIMN63N_LC_13_10_3  (
            .in0(N__40901),
            .in1(N__42507),
            .in2(_gnd_net_),
            .in3(N__40892),
            .lcout(\ALU.un9_addsub_cry_2_c_RNIMN63NZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_3_c_RNI4L7RO_LC_13_10_4 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_3_c_RNI4L7RO_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_3_c_RNI4L7RO_LC_13_10_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.un9_addsub_cry_3_c_RNI4L7RO_LC_13_10_4  (
            .in0(N__40877),
            .in1(N__42503),
            .in2(_gnd_net_),
            .in3(N__40862),
            .lcout(\ALU.un9_addsub_cry_3_c_RNI4L7ROZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_4_c_RNIUEDLM_LC_13_10_5 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_4_c_RNIUEDLM_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_4_c_RNIUEDLM_LC_13_10_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.un9_addsub_cry_4_c_RNIUEDLM_LC_13_10_5  (
            .in0(N__42504),
            .in1(N__42563),
            .in2(_gnd_net_),
            .in3(N__42554),
            .lcout(\ALU.un9_addsub_cry_4_c_RNIUEDLMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.un9_addsub_cry_5_c_RNI26HCN_LC_13_10_6 .C_ON=1'b0;
    defparam \ALU.un9_addsub_cry_5_c_RNI26HCN_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \ALU.un9_addsub_cry_5_c_RNI26HCN_LC_13_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.un9_addsub_cry_5_c_RNI26HCN_LC_13_10_6  (
            .in0(N__42539),
            .in1(N__42505),
            .in2(_gnd_net_),
            .in3(N__42419),
            .lcout(\ALU.un9_addsub_cry_5_c_RNI26HCNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_7_LC_13_11_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_7_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_7_LC_13_11_0 .LUT_INIT=16'b0001110100111111;
    LogicCell40 \ALU.a_15_m2_ns_1_7_LC_13_11_0  (
            .in0(N__44226),
            .in1(N__47320),
            .in2(N__43963),
            .in3(N__43767),
            .lcout(\ALU.a_15_m2_ns_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIP43E91_7_LC_13_11_2 .C_ON=1'b0;
    defparam \ALU.d_RNIP43E91_7_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIP43E91_7_LC_13_11_2 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \ALU.d_RNIP43E91_7_LC_13_11_2  (
            .in0(N__42404),
            .in1(N__44537),
            .in2(N__46748),
            .in3(N__44227),
            .lcout(),
            .ltout(\ALU.d_RNIP43E91Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIL4SQK2_7_LC_13_11_3 .C_ON=1'b0;
    defparam \ALU.d_RNIL4SQK2_7_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIL4SQK2_7_LC_13_11_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ALU.d_RNIL4SQK2_7_LC_13_11_3  (
            .in0(N__46393),
            .in1(_gnd_net_),
            .in2(N__42389),
            .in3(N__42386),
            .lcout(),
            .ltout(\ALU.a_15_m5_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIIIPM081_7_LC_13_11_4 .C_ON=1'b0;
    defparam \ALU.d_RNIIIPM081_7_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIIIPM081_7_LC_13_11_4 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ALU.d_RNIIIPM081_7_LC_13_11_4  (
            .in0(N__46003),
            .in1(N__42371),
            .in2(N__42356),
            .in3(N__42353),
            .lcout(\ALU.d_RNIIIPM081Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_0_LC_13_12_0 .C_ON=1'b0;
    defparam \ALU.d_0_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.d_0_LC_13_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_0_LC_13_12_0  (
            .in0(N__48578),
            .in1(N__42297),
            .in2(_gnd_net_),
            .in3(N__42264),
            .lcout(\ALU.dZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47641),
            .ce(N__43340),
            .sr(_gnd_net_));
    defparam \ALU.d_2_LC_13_12_2 .C_ON=1'b0;
    defparam \ALU.d_2_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.d_2_LC_13_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_2_LC_13_12_2  (
            .in0(N__48579),
            .in1(N__42126),
            .in2(_gnd_net_),
            .in3(N__42098),
            .lcout(\ALU.dZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47641),
            .ce(N__43340),
            .sr(_gnd_net_));
    defparam \ALU.d_3_LC_13_12_3 .C_ON=1'b0;
    defparam \ALU.d_3_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.d_3_LC_13_12_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.d_3_LC_13_12_3  (
            .in0(N__49441),
            .in1(N__48580),
            .in2(_gnd_net_),
            .in3(N__49360),
            .lcout(\ALU.dZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47641),
            .ce(N__43340),
            .sr(_gnd_net_));
    defparam \ALU.d_5_LC_13_12_5 .C_ON=1'b0;
    defparam \ALU.d_5_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.d_5_LC_13_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_5_LC_13_12_5  (
            .in0(N__48585),
            .in1(N__49044),
            .in2(_gnd_net_),
            .in3(N__49089),
            .lcout(\ALU.dZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47641),
            .ce(N__43340),
            .sr(_gnd_net_));
    defparam \ALU.d_6_LC_13_12_6 .C_ON=1'b0;
    defparam \ALU.d_6_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \ALU.d_6_LC_13_12_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.d_6_LC_13_12_6  (
            .in0(N__48917),
            .in1(N__48587),
            .in2(_gnd_net_),
            .in3(N__48863),
            .lcout(\ALU.dZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47641),
            .ce(N__43340),
            .sr(_gnd_net_));
    defparam \ALU.d_7_LC_13_12_7 .C_ON=1'b0;
    defparam \ALU.d_7_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \ALU.d_7_LC_13_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_7_LC_13_12_7  (
            .in0(N__48586),
            .in1(N__48790),
            .in2(_gnd_net_),
            .in3(N__48684),
            .lcout(\ALU.dZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47641),
            .ce(N__43340),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIHUEJ_3_LC_13_13_6 .C_ON=1'b0;
    defparam \ALU.f_RNIHUEJ_3_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIHUEJ_3_LC_13_13_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.f_RNIHUEJ_3_LC_13_13_6  (
            .in0(N__43261),
            .in1(N__49303),
            .in2(_gnd_net_),
            .in3(N__45119),
            .lcout(\ALU.f_RNIHUEJZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_4_LC_13_14_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_4_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_4_LC_13_14_0 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.a_15_m2_ns_1_4_LC_13_14_0  (
            .in0(N__47323),
            .in1(N__44224),
            .in2(N__43967),
            .in3(N__43768),
            .lcout(\ALU.a_15_m2_ns_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNISSLDG1_6_LC_13_14_1 .C_ON=1'b0;
    defparam \ALU.d_RNISSLDG1_6_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNISSLDG1_6_LC_13_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNISSLDG1_6_LC_13_14_1  (
            .in0(N__44540),
            .in1(N__43232),
            .in2(_gnd_net_),
            .in3(N__43211),
            .lcout(),
            .ltout(\ALU.rshift_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIC1CRK1_4_LC_13_14_2 .C_ON=1'b0;
    defparam \ALU.d_RNIC1CRK1_4_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIC1CRK1_4_LC_13_14_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ALU.d_RNIC1CRK1_4_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__43193),
            .in2(N__43025),
            .in3(N__43022),
            .lcout(),
            .ltout(\ALU.a_15_m3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIBK80K2_4_LC_13_14_3 .C_ON=1'b0;
    defparam \ALU.d_RNIBK80K2_4_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIBK80K2_4_LC_13_14_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ALU.d_RNIBK80K2_4_LC_13_14_3  (
            .in0(N__46384),
            .in1(_gnd_net_),
            .in2(N__43001),
            .in3(N__44942),
            .lcout(\ALU.a_15_m5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNINL83B_4_LC_13_14_4 .C_ON=1'b0;
    defparam \ALU.d_RNINL83B_4_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNINL83B_4_LC_13_14_4 .LUT_INIT=16'b1000011001100111;
    LogicCell40 \ALU.d_RNINL83B_4_LC_13_14_4  (
            .in0(N__47324),
            .in1(N__42993),
            .in2(N__42707),
            .in3(N__42697),
            .lcout(),
            .ltout(\ALU.a_15_m2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI0SA7U_4_LC_13_14_5 .C_ON=1'b0;
    defparam \ALU.d_RNI0SA7U_4_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI0SA7U_4_LC_13_14_5 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \ALU.d_RNI0SA7U_4_LC_13_14_5  (
            .in0(N__44225),
            .in1(N__44539),
            .in2(N__44972),
            .in3(N__44969),
            .lcout(\ALU.a_15_m4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMA3938_4_LC_13_14_6 .C_ON=1'b0;
    defparam \ALU.d_RNIMA3938_4_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMA3938_4_LC_13_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.d_RNIMA3938_4_LC_13_14_6  (
            .in0(N__46085),
            .in1(N__44936),
            .in2(_gnd_net_),
            .in3(N__44921),
            .lcout(\ALU.d_RNIMA3938Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_3_LC_13_15_3 .C_ON=1'b0;
    defparam \ALU.a_3_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \ALU.a_3_LC_13_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.a_3_LC_13_15_3  (
            .in0(N__48577),
            .in1(N__49450),
            .in2(_gnd_net_),
            .in3(N__49378),
            .lcout(a_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47660),
            .ce(N__44888),
            .sr(_gnd_net_));
    defparam \FTDI.TXshift_1_LC_14_5_5 .C_ON=1'b0;
    defparam \FTDI.TXshift_1_LC_14_5_5 .SEQ_MODE=4'b1000;
    defparam \FTDI.TXshift_1_LC_14_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \FTDI.TXshift_1_LC_14_5_5  (
            .in0(N__44780),
            .in1(N__44567),
            .in2(_gnd_net_),
            .in3(N__44769),
            .lcout(\FTDI.TXshiftZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVFTDI.TXshift_1C_net ),
            .ce(N__44666),
            .sr(_gnd_net_));
    defparam TXbuffer_5_LC_14_7_5.C_ON=1'b0;
    defparam TXbuffer_5_LC_14_7_5.SEQ_MODE=4'b1000;
    defparam TXbuffer_5_LC_14_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_5_LC_14_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44645),
            .lcout(TXbufferZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47608),
            .ce(N__44558),
            .sr(_gnd_net_));
    defparam TXbuffer_1_LC_14_7_7.C_ON=1'b0;
    defparam TXbuffer_1_LC_14_7_7.SEQ_MODE=4'b1000;
    defparam TXbuffer_1_LC_14_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 TXbuffer_1_LC_14_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44600),
            .lcout(TXbufferZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47608),
            .ce(N__44558),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIJ75U41_6_LC_14_8_2 .C_ON=1'b0;
    defparam \ALU.d_RNIJ75U41_6_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIJ75U41_6_LC_14_8_2 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \ALU.d_RNIJ75U41_6_LC_14_8_2  (
            .in0(N__44219),
            .in1(N__46400),
            .in2(N__44538),
            .in3(N__44240),
            .lcout(\ALU.d_RNIJ75U41Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.a_15_m2_ns_1_6_LC_14_9_0 .C_ON=1'b0;
    defparam \ALU.a_15_m2_ns_1_6_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \ALU.a_15_m2_ns_1_6_LC_14_9_0 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \ALU.a_15_m2_ns_1_6_LC_14_9_0  (
            .in0(N__47309),
            .in1(N__44223),
            .in2(N__43962),
            .in3(N__43763),
            .lcout(),
            .ltout(\ALU.a_15_m2_ns_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIMBENA_6_LC_14_9_1 .C_ON=1'b0;
    defparam \ALU.d_RNIMBENA_6_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIMBENA_6_LC_14_9_1 .LUT_INIT=16'b1000011001100111;
    LogicCell40 \ALU.d_RNIMBENA_6_LC_14_9_1  (
            .in0(N__47310),
            .in1(N__46727),
            .in2(N__46484),
            .in3(N__46481),
            .lcout(\ALU.a_15_m2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNI7VNOJ2_6_LC_14_9_3 .C_ON=1'b0;
    defparam \ALU.d_RNI7VNOJ2_6_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNI7VNOJ2_6_LC_14_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ALU.d_RNI7VNOJ2_6_LC_14_9_3  (
            .in0(N__46392),
            .in1(N__46229),
            .in2(_gnd_net_),
            .in3(N__46208),
            .lcout(),
            .ltout(\ALU.a_15_m5_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILPR7TQ_6_LC_14_9_4 .C_ON=1'b0;
    defparam \ALU.d_RNILPR7TQ_6_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILPR7TQ_6_LC_14_9_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.d_RNILPR7TQ_6_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__46033),
            .in2(N__45638),
            .in3(N__45635),
            .lcout(\ALU.d_RNILPR7TQZ0Z_6 ),
            .ltout(\ALU.d_RNILPR7TQZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.h_6_LC_14_9_5 .C_ON=1'b0;
    defparam \ALU.h_6_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \ALU.h_6_LC_14_9_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \ALU.h_6_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__48509),
            .in2(N__45626),
            .in3(N__48856),
            .lcout(\ALU.hZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47616),
            .ce(N__45557),
            .sr(_gnd_net_));
    defparam \ALU.f_RNIJ0FJ_4_LC_14_10_3 .C_ON=1'b0;
    defparam \ALU.f_RNIJ0FJ_4_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \ALU.f_RNIJ0FJ_4_LC_14_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.f_RNIJ0FJ_4_LC_14_10_3  (
            .in0(N__45121),
            .in1(N__45409),
            .in2(_gnd_net_),
            .in3(N__49144),
            .lcout(\ALU.f_RNIJ0FJZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIU60L_7_LC_14_11_6 .C_ON=1'b0;
    defparam \ALU.d_RNIU60L_7_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIU60L_7_LC_14_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNIU60L_7_LC_14_11_6  (
            .in0(N__45373),
            .in1(N__45349),
            .in2(_gnd_net_),
            .in3(N__45312),
            .lcout(\ALU.d_RNIU60LZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.d_RNILAR7_3_LC_14_11_7 .C_ON=1'b0;
    defparam \ALU.d_RNILAR7_3_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNILAR7_3_LC_14_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ALU.d_RNILAR7_3_LC_14_11_7  (
            .in0(N__45175),
            .in1(N__45148),
            .in2(_gnd_net_),
            .in3(N__45120),
            .lcout(\ALU.d_RNILAR7Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU.b_3_LC_14_12_0 .C_ON=1'b0;
    defparam \ALU.b_3_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \ALU.b_3_LC_14_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_3_LC_14_12_0  (
            .in0(N__48592),
            .in1(N__49443),
            .in2(_gnd_net_),
            .in3(N__49368),
            .lcout(\ALU.bZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47636),
            .ce(N__47401),
            .sr(_gnd_net_));
    defparam \ALU.b_4_LC_14_12_1 .C_ON=1'b0;
    defparam \ALU.b_4_LC_14_12_1 .SEQ_MODE=4'b1000;
    defparam \ALU.b_4_LC_14_12_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ALU.b_4_LC_14_12_1  (
            .in0(N__49244),
            .in1(N__48595),
            .in2(_gnd_net_),
            .in3(N__49211),
            .lcout(\ALU.bZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47636),
            .ce(N__47401),
            .sr(_gnd_net_));
    defparam \ALU.b_5_LC_14_12_2 .C_ON=1'b0;
    defparam \ALU.b_5_LC_14_12_2 .SEQ_MODE=4'b1000;
    defparam \ALU.b_5_LC_14_12_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_5_LC_14_12_2  (
            .in0(N__48593),
            .in1(N__49094),
            .in2(_gnd_net_),
            .in3(N__49049),
            .lcout(\ALU.bZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47636),
            .ce(N__47401),
            .sr(_gnd_net_));
    defparam \ALU.b_6_LC_14_12_3 .C_ON=1'b0;
    defparam \ALU.b_6_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \ALU.b_6_LC_14_12_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ALU.b_6_LC_14_12_3  (
            .in0(N__48916),
            .in1(N__48596),
            .in2(_gnd_net_),
            .in3(N__48880),
            .lcout(\ALU.bZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47636),
            .ce(N__47401),
            .sr(_gnd_net_));
    defparam \ALU.b_7_LC_14_12_4 .C_ON=1'b0;
    defparam \ALU.b_7_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \ALU.b_7_LC_14_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_7_LC_14_12_4  (
            .in0(N__48594),
            .in1(N__48791),
            .in2(_gnd_net_),
            .in3(N__48695),
            .lcout(\ALU.bZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47636),
            .ce(N__47401),
            .sr(_gnd_net_));
    defparam \ALU.b_8_LC_14_12_5 .C_ON=1'b0;
    defparam \ALU.b_8_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \ALU.b_8_LC_14_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ALU.b_8_LC_14_12_5  (
            .in0(N__48581),
            .in1(N__47892),
            .in2(_gnd_net_),
            .in3(N__47810),
            .lcout(\ALU.bZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47636),
            .ce(N__47401),
            .sr(_gnd_net_));
    defparam \ALU.d_RNIHRFPB_7_LC_14_13_6 .C_ON=1'b0;
    defparam \ALU.d_RNIHRFPB_7_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \ALU.d_RNIHRFPB_7_LC_14_13_6 .LUT_INIT=16'b1001010100101011;
    LogicCell40 \ALU.d_RNIHRFPB_7_LC_14_13_6  (
            .in0(N__47322),
            .in1(N__47105),
            .in2(N__46991),
            .in3(N__46964),
            .lcout(\ALU.a_15_m2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
