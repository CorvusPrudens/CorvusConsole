module dromdata(
    input wire CLK,
    input wire [15:0] address,
    output wire [15:0] data
    );

    (* rom_style = "block" *) reg [15:0] dintern = 16'b0;

    always @( * ) begin
        case (address)
        16'h0000: dintern = 16'h001F;
        16'h0001: dintern = 16'h0011;
        16'h0002: dintern = 16'h001F;
        16'h0003: dintern = 16'h001F;
        16'h0004: dintern = 16'h0011;
        16'h0005: dintern = 16'h001F;
        16'h0006: dintern = 16'h001F;
        16'h0007: dintern = 16'h0011;
        16'h0008: dintern = 16'h001F;
        16'h0009: dintern = 16'h001F;
        16'h000A: dintern = 16'h0011;
        16'h000B: dintern = 16'h001F;
        16'h000C: dintern = 16'h001F;
        16'h000D: dintern = 16'h0011;
        16'h000E: dintern = 16'h001F;
        16'h000F: dintern = 16'h001F;
        16'h0010: dintern = 16'h0011;
        16'h0011: dintern = 16'h001F;
        16'h0012: dintern = 16'h001F;
        16'h0013: dintern = 16'h0011;
        16'h0014: dintern = 16'h001F;
        16'h0015: dintern = 16'h001F;
        16'h0016: dintern = 16'h0011;
        16'h0017: dintern = 16'h001F;
        16'h0018: dintern = 16'h001F;
        16'h0019: dintern = 16'h0011;
        16'h001A: dintern = 16'h001F;
        16'h001B: dintern = 16'h001F;
        16'h001C: dintern = 16'h0011;
        16'h001D: dintern = 16'h001F;
        16'h001E: dintern = 16'h001F;
        16'h001F: dintern = 16'h0011;
        16'h0020: dintern = 16'h001F;
        16'h0021: dintern = 16'h001F;
        16'h0022: dintern = 16'h0011;
        16'h0023: dintern = 16'h001F;
        16'h0024: dintern = 16'h001F;
        16'h0025: dintern = 16'h0011;
        16'h0026: dintern = 16'h001F;
        16'h0027: dintern = 16'h001F;
        16'h0028: dintern = 16'h0011;
        16'h0029: dintern = 16'h001F;
        16'h002A: dintern = 16'h001F;
        16'h002B: dintern = 16'h0011;
        16'h002C: dintern = 16'h001F;
        16'h002D: dintern = 16'h001F;
        16'h002E: dintern = 16'h0011;
        16'h002F: dintern = 16'h001F;
        16'h0030: dintern = 16'h001F;
        16'h0031: dintern = 16'h0011;
        16'h0032: dintern = 16'h001F;
        16'h0033: dintern = 16'h001F;
        16'h0034: dintern = 16'h0011;
        16'h0035: dintern = 16'h001F;
        16'h0036: dintern = 16'h001F;
        16'h0037: dintern = 16'h0011;
        16'h0038: dintern = 16'h001F;
        16'h0039: dintern = 16'h001F;
        16'h003A: dintern = 16'h0011;
        16'h003B: dintern = 16'h001F;
        16'h003C: dintern = 16'h001F;
        16'h003D: dintern = 16'h0011;
        16'h003E: dintern = 16'h001F;
        16'h003F: dintern = 16'h001F;
        16'h0040: dintern = 16'h0011;
        16'h0041: dintern = 16'h001F;
        16'h0042: dintern = 16'h001F;
        16'h0043: dintern = 16'h0011;
        16'h0044: dintern = 16'h001F;
        16'h0045: dintern = 16'h001F;
        16'h0046: dintern = 16'h0011;
        16'h0047: dintern = 16'h001F;
        16'h0048: dintern = 16'h001F;
        16'h0049: dintern = 16'h0011;
        16'h004A: dintern = 16'h001F;
        16'h004B: dintern = 16'h001F;
        16'h004C: dintern = 16'h0011;
        16'h004D: dintern = 16'h001F;
        16'h004E: dintern = 16'h001F;
        16'h004F: dintern = 16'h0011;
        16'h0050: dintern = 16'h001F;
        16'h0051: dintern = 16'h001F;
        16'h0052: dintern = 16'h0011;
        16'h0053: dintern = 16'h001F;
        16'h0054: dintern = 16'h001F;
        16'h0055: dintern = 16'h0011;
        16'h0056: dintern = 16'h001F;
        16'h0057: dintern = 16'h001F;
        16'h0058: dintern = 16'h0011;
        16'h0059: dintern = 16'h001F;
        16'h005A: dintern = 16'h001F;
        16'h005B: dintern = 16'h0011;
        16'h005C: dintern = 16'h001F;
        16'h005D: dintern = 16'h001F;
        16'h005E: dintern = 16'h001F;
        16'h005F: dintern = 16'h001F;
        16'h0060: dintern = 16'h0000;
        16'h0061: dintern = 16'h0000;
        16'h0062: dintern = 16'h0000;
        16'h0063: dintern = 16'h0000;
        16'h0064: dintern = 16'h0017;
        16'h0065: dintern = 16'h0000;
        16'h0066: dintern = 16'h0003;
        16'h0067: dintern = 16'h0000;
        16'h0068: dintern = 16'h0003;
        16'h0069: dintern = 16'h001F;
        16'h006A: dintern = 16'h000A;
        16'h006B: dintern = 16'h001F;
        16'h006C: dintern = 16'h000A;
        16'h006D: dintern = 16'h001F;
        16'h006E: dintern = 16'h0005;
        16'h006F: dintern = 16'h0009;
        16'h0070: dintern = 16'h0004;
        16'h0071: dintern = 16'h0012;
        16'h0072: dintern = 16'h000F;
        16'h0073: dintern = 16'h0017;
        16'h0074: dintern = 16'h001C;
        16'h0075: dintern = 16'h0000;
        16'h0076: dintern = 16'h0003;
        16'h0077: dintern = 16'h0000;
        16'h0078: dintern = 16'h0000;
        16'h0079: dintern = 16'h000E;
        16'h007A: dintern = 16'h0011;
        16'h007B: dintern = 16'h0011;
        16'h007C: dintern = 16'h000E;
        16'h007D: dintern = 16'h0000;
        16'h007E: dintern = 16'h0005;
        16'h007F: dintern = 16'h0002;
        16'h0080: dintern = 16'h0005;
        16'h0081: dintern = 16'h0004;
        16'h0082: dintern = 16'h000E;
        16'h0083: dintern = 16'h0004;
        16'h0084: dintern = 16'h0010;
        16'h0085: dintern = 16'h0008;
        16'h0086: dintern = 16'h0000;
        16'h0087: dintern = 16'h0004;
        16'h0088: dintern = 16'h0004;
        16'h0089: dintern = 16'h0004;
        16'h008A: dintern = 16'h0000;
        16'h008B: dintern = 16'h0010;
        16'h008C: dintern = 16'h0000;
        16'h008D: dintern = 16'h0018;
        16'h008E: dintern = 16'h0004;
        16'h008F: dintern = 16'h0003;
        16'h0090: dintern = 16'h001E;
        16'h0091: dintern = 16'h0011;
        16'h0092: dintern = 16'h000F;
        16'h0093: dintern = 16'h0002;
        16'h0094: dintern = 16'h001F;
        16'h0095: dintern = 16'h0000;
        16'h0096: dintern = 16'h0019;
        16'h0097: dintern = 16'h0015;
        16'h0098: dintern = 16'h0012;
        16'h0099: dintern = 16'h0011;
        16'h009A: dintern = 16'h0015;
        16'h009B: dintern = 16'h000A;
        16'h009C: dintern = 16'h0007;
        16'h009D: dintern = 16'h0004;
        16'h009E: dintern = 16'h001F;
        16'h009F: dintern = 16'h0017;
        16'h00A0: dintern = 16'h0015;
        16'h00A1: dintern = 16'h0009;
        16'h00A2: dintern = 16'h001E;
        16'h00A3: dintern = 16'h0015;
        16'h00A4: dintern = 16'h001D;
        16'h00A5: dintern = 16'h0019;
        16'h00A6: dintern = 16'h0005;
        16'h00A7: dintern = 16'h0003;
        16'h00A8: dintern = 16'h001F;
        16'h00A9: dintern = 16'h0015;
        16'h00AA: dintern = 16'h001F;
        16'h00AB: dintern = 16'h0017;
        16'h00AC: dintern = 16'h0015;
        16'h00AD: dintern = 16'h000F;
        16'h00AE: dintern = 16'h0000;
        16'h00AF: dintern = 16'h000A;
        16'h00B0: dintern = 16'h0000;
        16'h00B1: dintern = 16'h0010;
        16'h00B2: dintern = 16'h000A;
        16'h00B3: dintern = 16'h0000;
        16'h00B4: dintern = 16'h0004;
        16'h00B5: dintern = 16'h000A;
        16'h00B6: dintern = 16'h0011;
        16'h00B7: dintern = 16'h000A;
        16'h00B8: dintern = 16'h000A;
        16'h00B9: dintern = 16'h000A;
        16'h00BA: dintern = 16'h0011;
        16'h00BB: dintern = 16'h000A;
        16'h00BC: dintern = 16'h0004;
        16'h00BD: dintern = 16'h0001;
        16'h00BE: dintern = 16'h0015;
        16'h00BF: dintern = 16'h0003;
        16'h00C0: dintern = 16'h000E;
        16'h00C1: dintern = 16'h0015;
        16'h00C2: dintern = 16'h0016;
        16'h00C3: dintern = 16'h001E;
        16'h00C4: dintern = 16'h0005;
        16'h00C5: dintern = 16'h001E;
        16'h00C6: dintern = 16'h001F;
        16'h00C7: dintern = 16'h0015;
        16'h00C8: dintern = 16'h000A;
        16'h00C9: dintern = 16'h000E;
        16'h00CA: dintern = 16'h0011;
        16'h00CB: dintern = 16'h0011;
        16'h00CC: dintern = 16'h001F;
        16'h00CD: dintern = 16'h0011;
        16'h00CE: dintern = 16'h000E;
        16'h00CF: dintern = 16'h001F;
        16'h00D0: dintern = 16'h0015;
        16'h00D1: dintern = 16'h0015;
        16'h00D2: dintern = 16'h001F;
        16'h00D3: dintern = 16'h0005;
        16'h00D4: dintern = 16'h0005;
        16'h00D5: dintern = 16'h000E;
        16'h00D6: dintern = 16'h0015;
        16'h00D7: dintern = 16'h001D;
        16'h00D8: dintern = 16'h001F;
        16'h00D9: dintern = 16'h0004;
        16'h00DA: dintern = 16'h001F;
        16'h00DB: dintern = 16'h0011;
        16'h00DC: dintern = 16'h001F;
        16'h00DD: dintern = 16'h0011;
        16'h00DE: dintern = 16'h0008;
        16'h00DF: dintern = 16'h0010;
        16'h00E0: dintern = 16'h000F;
        16'h00E1: dintern = 16'h001F;
        16'h00E2: dintern = 16'h0004;
        16'h00E3: dintern = 16'h001B;
        16'h00E4: dintern = 16'h001F;
        16'h00E5: dintern = 16'h0010;
        16'h00E6: dintern = 16'h0010;
        16'h00E7: dintern = 16'h001F;
        16'h00E8: dintern = 16'h0006;
        16'h00E9: dintern = 16'h001F;
        16'h00EA: dintern = 16'h001F;
        16'h00EB: dintern = 16'h000E;
        16'h00EC: dintern = 16'h001F;
        16'h00ED: dintern = 16'h000E;
        16'h00EE: dintern = 16'h0011;
        16'h00EF: dintern = 16'h000E;
        16'h00F0: dintern = 16'h001F;
        16'h00F1: dintern = 16'h0005;
        16'h00F2: dintern = 16'h0002;
        16'h00F3: dintern = 16'h000E;
        16'h00F4: dintern = 16'h0019;
        16'h00F5: dintern = 16'h001E;
        16'h00F6: dintern = 16'h001F;
        16'h00F7: dintern = 16'h000D;
        16'h00F8: dintern = 16'h0016;
        16'h00F9: dintern = 16'h0012;
        16'h00FA: dintern = 16'h0015;
        16'h00FB: dintern = 16'h0009;
        16'h00FC: dintern = 16'h0001;
        16'h00FD: dintern = 16'h001F;
        16'h00FE: dintern = 16'h0001;
        16'h00FF: dintern = 16'h000F;
        16'h0100: dintern = 16'h0010;
        16'h0101: dintern = 16'h001F;
        16'h0102: dintern = 16'h0007;
        16'h0103: dintern = 16'h0018;
        16'h0104: dintern = 16'h0007;
        16'h0105: dintern = 16'h001F;
        16'h0106: dintern = 16'h000C;
        16'h0107: dintern = 16'h001F;
        16'h0108: dintern = 16'h001B;
        16'h0109: dintern = 16'h0004;
        16'h010A: dintern = 16'h001B;
        16'h010B: dintern = 16'h0003;
        16'h010C: dintern = 16'h001C;
        16'h010D: dintern = 16'h0003;
        16'h010E: dintern = 16'h0019;
        16'h010F: dintern = 16'h0015;
        16'h0110: dintern = 16'h0013;
        16'h0111: dintern = 16'h001F;
        16'h0112: dintern = 16'h0011;
        16'h0113: dintern = 16'h0011;
        16'h0114: dintern = 16'h0002;
        16'h0115: dintern = 16'h0004;
        16'h0116: dintern = 16'h0008;
        16'h0117: dintern = 16'h0011;
        16'h0118: dintern = 16'h0011;
        16'h0119: dintern = 16'h001F;
        16'h011A: dintern = 16'h0002;
        16'h011B: dintern = 16'h0001;
        16'h011C: dintern = 16'h0002;
        16'h011D: dintern = 16'h0010;
        16'h011E: dintern = 16'h0010;
        16'h011F: dintern = 16'h0010;
        16'h0120: dintern = 16'h0001;
        16'h0121: dintern = 16'h0002;
        16'h0122: dintern = 16'h0000;
        16'h0123: dintern = 16'h001A;
        16'h0124: dintern = 16'h0016;
        16'h0125: dintern = 16'h001C;
        16'h0126: dintern = 16'h001F;
        16'h0127: dintern = 16'h0012;
        16'h0128: dintern = 16'h000C;
        16'h0129: dintern = 16'h000C;
        16'h012A: dintern = 16'h0012;
        16'h012B: dintern = 16'h0012;
        16'h012C: dintern = 16'h000C;
        16'h012D: dintern = 16'h0012;
        16'h012E: dintern = 16'h001F;
        16'h012F: dintern = 16'h000C;
        16'h0130: dintern = 16'h001A;
        16'h0131: dintern = 16'h0016;
        16'h0132: dintern = 16'h0004;
        16'h0133: dintern = 16'h001E;
        16'h0134: dintern = 16'h0005;
        16'h0135: dintern = 16'h000C;
        16'h0136: dintern = 16'h002A;
        16'h0137: dintern = 16'h001E;
        16'h0138: dintern = 16'h001F;
        16'h0139: dintern = 16'h0002;
        16'h013A: dintern = 16'h001C;
        16'h013B: dintern = 16'h0000;
        16'h013C: dintern = 16'h001D;
        16'h013D: dintern = 16'h0000;
        16'h013E: dintern = 16'h0010;
        16'h013F: dintern = 16'h0020;
        16'h0140: dintern = 16'h001D;
        16'h0141: dintern = 16'h001F;
        16'h0142: dintern = 16'h000C;
        16'h0143: dintern = 16'h0012;
        16'h0144: dintern = 16'h0011;
        16'h0145: dintern = 16'h001F;
        16'h0146: dintern = 16'h0010;
        16'h0147: dintern = 16'h001E;
        16'h0148: dintern = 16'h000E;
        16'h0149: dintern = 16'h001E;
        16'h014A: dintern = 16'h001E;
        16'h014B: dintern = 16'h0002;
        16'h014C: dintern = 16'h001C;
        16'h014D: dintern = 16'h000C;
        16'h014E: dintern = 16'h0012;
        16'h014F: dintern = 16'h000C;
        16'h0150: dintern = 16'h003E;
        16'h0151: dintern = 16'h0012;
        16'h0152: dintern = 16'h000C;
        16'h0153: dintern = 16'h000C;
        16'h0154: dintern = 16'h0012;
        16'h0155: dintern = 16'h003E;
        16'h0156: dintern = 16'h001C;
        16'h0157: dintern = 16'h0002;
        16'h0158: dintern = 16'h0002;
        16'h0159: dintern = 16'h0014;
        16'h015A: dintern = 16'h001E;
        16'h015B: dintern = 16'h000A;
        16'h015C: dintern = 16'h0002;
        16'h015D: dintern = 16'h001F;
        16'h015E: dintern = 16'h0012;
        16'h015F: dintern = 16'h000E;
        16'h0160: dintern = 16'h0010;
        16'h0161: dintern = 16'h001E;
        16'h0162: dintern = 16'h000E;
        16'h0163: dintern = 16'h0018;
        16'h0164: dintern = 16'h000E;
        16'h0165: dintern = 16'h001E;
        16'h0166: dintern = 16'h001C;
        16'h0167: dintern = 16'h001E;
        16'h0168: dintern = 16'h0012;
        16'h0169: dintern = 16'h000C;
        16'h016A: dintern = 16'h0012;
        16'h016B: dintern = 16'h0006;
        16'h016C: dintern = 16'h0028;
        16'h016D: dintern = 16'h001E;
        16'h016E: dintern = 16'h001A;
        16'h016F: dintern = 16'h001E;
        16'h0170: dintern = 16'h0016;
        16'h0171: dintern = 16'h0004;
        16'h0172: dintern = 16'h001B;
        16'h0173: dintern = 16'h0011;
        16'h0174: dintern = 16'h0000;
        16'h0175: dintern = 16'h001B;
        16'h0176: dintern = 16'h0000;
        16'h0177: dintern = 16'h0011;
        16'h0178: dintern = 16'h001B;
        16'h0179: dintern = 16'h0004;
        16'h017A: dintern = 16'h0002;
        16'h017B: dintern = 16'h0003;
        16'h017C: dintern = 16'h0001;
        16'h017D: dintern = 16'h001F;
        16'h017E: dintern = 16'h001F;
        16'h017F: dintern = 16'h001F;
        16'h0180: dintern = 16'h0000;
        16'h0181: dintern = 16'h0000;
        16'h0182: dintern = 16'h0000;
        16'h0183: dintern = 16'h4600;
        16'h0184: dintern = 16'hE700;
        16'h0185: dintern = 16'h7700;
        16'h0186: dintern = 16'h3BC0;
        16'h0187: dintern = 16'h0FE0;
        16'h0188: dintern = 16'h17E0;
        16'h0189: dintern = 16'h1F20;
        16'h018A: dintern = 16'h0FE0;
        16'h018B: dintern = 16'h0400;
        16'h018C: dintern = 16'h0000;
        16'h018D: dintern = 16'h0000;
        16'h018E: dintern = 16'h0000;
        16'h018F: dintern = 16'h0000;
        16'h0190: dintern = 16'h0000;
        16'h0191: dintern = 16'h0000;
        16'h0192: dintern = 16'h0000;
        16'h0193: dintern = 16'h6000;
        16'h0194: dintern = 16'h3000;
        16'h0195: dintern = 16'h3700;
        16'h0196: dintern = 16'h17C0;
        16'h0197: dintern = 16'h09E0;
        16'h0198: dintern = 16'h0FE0;
        16'h0199: dintern = 16'h1F20;
        16'h019A: dintern = 16'h1FE0;
        16'h019B: dintern = 16'h1800;
        16'h019C: dintern = 16'h0000;
        16'h019D: dintern = 16'h0000;
        16'h019E: dintern = 16'h0000;
        16'h019F: dintern = 16'h0000;
        16'h01A0: dintern = 16'h0000;
        16'h01A1: dintern = 16'h0000;
        16'h01A2: dintern = 16'h0000;
        16'h01A3: dintern = 16'h3000;
        16'h01A4: dintern = 16'h3800;
        16'h01A5: dintern = 16'h1BC0;
        16'h01A6: dintern = 16'h1BE0;
        16'h01A7: dintern = 16'h0A70;
        16'h01A8: dintern = 16'h05F0;
        16'h01A9: dintern = 16'h0790;
        16'h01AA: dintern = 16'h0FF0;
        16'h01AB: dintern = 16'h0C00;
        16'h01AC: dintern = 16'h0800;
        16'h01AD: dintern = 16'h0000;
        16'h01AE: dintern = 16'h0000;
        16'h01AF: dintern = 16'h0000;
        16'h01B0: dintern = 16'h0000;
        16'h01B1: dintern = 16'h0000;
        16'h01B2: dintern = 16'h0000;
        16'h01B3: dintern = 16'h0800;
        16'h01B4: dintern = 16'h1800;
        16'h01B5: dintern = 16'h1DE0;
        16'h01B6: dintern = 16'h0DF0;
        16'h01B7: dintern = 16'h07B8;
        16'h01B8: dintern = 16'h0678;
        16'h01B9: dintern = 16'h07C8;
        16'h01BA: dintern = 16'h0F78;
        16'h01BB: dintern = 16'h0E00;
        16'h01BC: dintern = 16'h0C00;
        16'h01BD: dintern = 16'h0000;
        16'h01BE: dintern = 16'h0000;
        16'h01BF: dintern = 16'h0000;
        16'h01C0: dintern = 16'h0000;
        16'h01C1: dintern = 16'h0000;
        16'h01C2: dintern = 16'h0000;
        16'h01C3: dintern = 16'h0000;
        16'h01C4: dintern = 16'h1800;
        16'h01C5: dintern = 16'h1BC0;
        16'h01C6: dintern = 16'h1BE0;
        16'h01C7: dintern = 16'h0F70;
        16'h01C8: dintern = 16'h0CF0;
        16'h01C9: dintern = 16'h1F90;
        16'h01CA: dintern = 16'h3EF0;
        16'h01CB: dintern = 16'h7C00;
        16'h01CC: dintern = 16'h7800;
        16'h01CD: dintern = 16'h0000;
        16'h01CE: dintern = 16'h0000;
        16'h01CF: dintern = 16'h0000;
        16'h01D0: dintern = 16'h0000;
        16'h01D1: dintern = 16'h0000;
        16'h01D2: dintern = 16'h0000;
        16'h01D3: dintern = 16'h0000;
        16'h01D4: dintern = 16'h1300;
        16'h01D5: dintern = 16'h1BC0;
        16'h01D6: dintern = 16'h1FE0;
        16'h01D7: dintern = 16'h0CF0;
        16'h01D8: dintern = 16'h37F0;
        16'h01D9: dintern = 16'hFF90;
        16'h01DA: dintern = 16'hFCF0;
        16'h01DB: dintern = 16'hC000;
        16'h01DC: dintern = 16'h0000;
        16'h01DD: dintern = 16'h0000;
        16'h01DE: dintern = 16'h0000;
        16'h01DF: dintern = 16'h0000;
        16'h01E0: dintern = 16'h0000;
        16'h01E1: dintern = 16'h0000;
        16'h01E2: dintern = 16'h0000;
        16'h01E3: dintern = 16'h0000;
        16'h01E4: dintern = 16'h0600;
        16'h01E5: dintern = 16'h2780;
        16'h01E6: dintern = 16'h33C0;
        16'h01E7: dintern = 16'h1FE0;
        16'h01E8: dintern = 16'hDFE0;
        16'h01E9: dintern = 16'hE720;
        16'h01EA: dintern = 16'h9FE0;
        16'h01EB: dintern = 16'h0000;
        16'h01EC: dintern = 16'h0000;
        16'h01ED: dintern = 16'h0000;
        16'h01EE: dintern = 16'h0000;
        16'h01EF: dintern = 16'h0000;
        16'h01F0: dintern = 16'h0000;
        16'h01F1: dintern = 16'h0000;
        16'h01F2: dintern = 16'h0000;
        16'h01F3: dintern = 16'h0C00;
        16'h01F4: dintern = 16'h0E00;
        16'h01F5: dintern = 16'h1700;
        16'h01F6: dintern = 16'h3F80;
        16'h01F7: dintern = 16'hBFC0;
        16'h01F8: dintern = 16'hDE40;
        16'h01F9: dintern = 16'h0FC0;
        16'h01FA: dintern = 16'h0640;
        16'h01FB: dintern = 16'h0000;
        16'h01FC: dintern = 16'h0000;
        16'h01FD: dintern = 16'h0000;
        16'h01FE: dintern = 16'h0000;
        16'h01FF: dintern = 16'h0000;
        16'h0200: dintern = 16'h0000;
        16'h0201: dintern = 16'h0000;
        16'h0202: dintern = 16'h0C00;
        16'h0203: dintern = 16'h0E00;
        16'h0204: dintern = 16'h0700;
        16'h0205: dintern = 16'h0380;
        16'h0206: dintern = 16'hAFC0;
        16'h0207: dintern = 16'hBFE0;
        16'h0208: dintern = 16'h7E60;
        16'h0209: dintern = 16'h37E0;
        16'h020A: dintern = 16'h0E60;
        16'h020B: dintern = 16'h0000;
        16'h020C: dintern = 16'h0000;
        16'h020D: dintern = 16'h0000;
        16'h020E: dintern = 16'h0000;
        16'h020F: dintern = 16'h0000;
        16'h0210: dintern = 16'h0000;
        16'h0211: dintern = 16'h0000;
        16'h0212: dintern = 16'h0600;
        16'h0213: dintern = 16'h0600;
        16'h0214: dintern = 16'h0300;
        16'h0215: dintern = 16'h6380;
        16'h0216: dintern = 16'h2FC0;
        16'h0217: dintern = 16'h1FE0;
        16'h0218: dintern = 16'h3F20;
        16'h0219: dintern = 16'h37E0;
        16'h021A: dintern = 16'h3720;
        16'h021B: dintern = 16'h0300;
        16'h021C: dintern = 16'h0000;
        16'h021D: dintern = 16'h0000;
        16'h021E: dintern = 16'h0000;
        16'h021F: dintern = 16'h0000;
        16'h0220: dintern = 16'h0000;
        16'h0221: dintern = 16'h0000;
        16'h0222: dintern = 16'h0180;
        16'h0223: dintern = 16'h01C0;
        16'h0224: dintern = 16'h31C0;
        16'h0225: dintern = 16'h38E0;
        16'h0226: dintern = 16'h0FE0;
        16'h0227: dintern = 16'h1FF0;
        16'h0228: dintern = 16'h1F90;
        16'h0229: dintern = 16'h3BF0;
        16'h022A: dintern = 16'h3B90;
        16'h022B: dintern = 16'h3180;
        16'h022C: dintern = 16'h0180;
        16'h022D: dintern = 16'h0000;
        16'h022E: dintern = 16'h0000;
        16'h022F: dintern = 16'h0000;
        16'h0230: dintern = 16'h0000;
        16'h0231: dintern = 16'h00C0;
        16'h0232: dintern = 16'h00C0;
        16'h0233: dintern = 16'h0060;
        16'h0234: dintern = 16'h1860;
        16'h0235: dintern = 16'h14F0;
        16'h0236: dintern = 16'h0FF0;
        16'h0237: dintern = 16'h0FF8;
        16'h0238: dintern = 16'h1FC8;
        16'h0239: dintern = 16'h1DF8;
        16'h023A: dintern = 16'h3CC8;
        16'h023B: dintern = 16'h38C0;
        16'h023C: dintern = 16'h30C0;
        16'h023D: dintern = 16'h00C0;
        16'h023E: dintern = 16'h0000;
        16'h023F: dintern = 16'h0000;
        16'h0240: dintern = 16'h0000;
        16'h0241: dintern = 16'h00C0;
        16'h0242: dintern = 16'h00C0;
        16'h0243: dintern = 16'h00C0;
        16'h0244: dintern = 16'h00E0;
        16'h0245: dintern = 16'h11E0;
        16'h0246: dintern = 16'h17E0;
        16'h0247: dintern = 16'h0FF0;
        16'h0248: dintern = 16'h1F90;
        16'h0249: dintern = 16'h1BF0;
        16'h024A: dintern = 16'h7990;
        16'h024B: dintern = 16'h61C0;
        16'h024C: dintern = 16'h00C0;
        16'h024D: dintern = 16'h00C0;
        16'h024E: dintern = 16'h0000;
        16'h024F: dintern = 16'h0000;
        16'h0250: dintern = 16'h0000;
        16'h0251: dintern = 16'h0000;
        16'h0252: dintern = 16'h0180;
        16'h0253: dintern = 16'h0180;
        16'h0254: dintern = 16'h0380;
        16'h0255: dintern = 16'hE7C0;
        16'h0256: dintern = 16'hFFC0;
        16'h0257: dintern = 16'hBFE0;
        16'h0258: dintern = 16'h0F20;
        16'h0259: dintern = 16'h1FE0;
        16'h025A: dintern = 16'h0F20;
        16'h025B: dintern = 16'h0600;
        16'h025C: dintern = 16'h0400;
        16'h025D: dintern = 16'h0000;
        16'h025E: dintern = 16'h0000;
        16'h025F: dintern = 16'h0000;
        16'h0260: dintern = 16'h0000;
        16'h0261: dintern = 16'h0000;
        16'h0262: dintern = 16'h0000;
        16'h0263: dintern = 16'h0000;
        16'h0264: dintern = 16'h0000;
        16'h0265: dintern = 16'h0000;
        16'h0266: dintern = 16'h0000;
        16'h0267: dintern = 16'h0000;
        16'h0268: dintern = 16'h0000;
        16'h0269: dintern = 16'h0000;
        16'h026A: dintern = 16'h0000;
        16'h026B: dintern = 16'h0000;
        16'h026C: dintern = 16'h0000;
        16'h026D: dintern = 16'h0000;
        16'h026E: dintern = 16'h0000;
        16'h026F: dintern = 16'h0000;
        16'h0270: dintern = 16'h0000;
        16'h0271: dintern = 16'h0000;
        16'h0272: dintern = 16'h0000;
        16'h0273: dintern = 16'h0000;
        16'h0274: dintern = 16'h0000;
        16'h0275: dintern = 16'h0000;
        16'h0276: dintern = 16'h0000;
        16'h0277: dintern = 16'h0000;
        16'h0278: dintern = 16'h0000;
        16'h0279: dintern = 16'h0000;
        16'h027A: dintern = 16'h0000;
        16'h027B: dintern = 16'h0000;
        16'h027C: dintern = 16'h0000;
        16'h027D: dintern = 16'h0000;
        16'h027E: dintern = 16'h0000;
        16'h027F: dintern = 16'h0000;
        16'h0280: dintern = 16'h0000;
        16'h0281: dintern = 16'h0000;
        16'h0282: dintern = 16'hFFFF;
        16'h0283: dintern = 16'h00FF;
        16'h0284: dintern = 16'h2020;
        16'h0285: dintern = 16'h0020;
        16'h0286: dintern = 16'h7D6E;
        16'h0287: dintern = 16'h00AB;
        16'h0288: dintern = 16'h22C5;
        16'h0289: dintern = 16'h0033;
        16'h028A: dintern = 16'h0049;
        16'h028B: dintern = 16'h0020;
        16'h028C: dintern = 16'h006E;
        16'h028D: dintern = 16'h006F;
        16'h028E: dintern = 16'h0077;
        16'h028F: dintern = 16'h0020;
        16'h0290: dintern = 16'h0068;
        16'h0291: dintern = 16'h0061;
        16'h0292: dintern = 16'h0076;
        16'h0293: dintern = 16'h0065;
        16'h0294: dintern = 16'h0020;
        16'h0295: dintern = 16'h002A;
        16'h0296: dintern = 16'h0073;
        16'h0297: dintern = 16'h0069;
        16'h0298: dintern = 16'h006D;
        16'h0299: dintern = 16'h0070;
        16'h029A: dintern = 16'h006C;
        16'h029B: dintern = 16'h0065;
        16'h029C: dintern = 16'h002A;
        16'h029D: dintern = 16'h0020;
        16'h029E: dintern = 16'h0077;
        16'h029F: dintern = 16'h006F;
        16'h02A0: dintern = 16'h0072;
        16'h02A1: dintern = 16'h006B;
        16'h02A2: dintern = 16'h0069;
        16'h02A3: dintern = 16'h006E;
        16'h02A4: dintern = 16'h0067;
        16'h02A5: dintern = 16'h0020;
        16'h02A6: dintern = 16'h0073;
        16'h02A7: dintern = 16'h0070;
        16'h02A8: dintern = 16'h0072;
        16'h02A9: dintern = 16'h0069;
        16'h02AA: dintern = 16'h0074;
        16'h02AB: dintern = 16'h0065;
        16'h02AC: dintern = 16'h0020;
        16'h02AD: dintern = 16'h0061;
        16'h02AE: dintern = 16'h006E;
        16'h02AF: dintern = 16'h0064;
        16'h02B0: dintern = 16'h0020;
        16'h02B1: dintern = 16'h0074;
        16'h02B2: dintern = 16'h0065;
        16'h02B3: dintern = 16'h0078;
        16'h02B4: dintern = 16'h0074;
        16'h02B5: dintern = 16'h0020;
        16'h02B6: dintern = 16'h0067;
        16'h02B7: dintern = 16'h0072;
        16'h02B8: dintern = 16'h0061;
        16'h02B9: dintern = 16'h0070;
        16'h02BA: dintern = 16'h0068;
        16'h02BB: dintern = 16'h0069;
        16'h02BC: dintern = 16'h0063;
        16'h02BD: dintern = 16'h0073;
        16'h02BE: dintern = 16'h0000;
        default: dintern = 16'h0;
    endcase
  end

  assign data = dintern;

endmodule
